module DSP (Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    Tile_X0Y0_E1BEG,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2BEG,
    Tile_X0Y0_E2BEGb,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6BEG,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4BEG,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_NN4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_SS4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W1END,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W2END,
    Tile_X0Y0_W2MID,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_W6END,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y0_WW4END,
    Tile_X0Y1_E1BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2BEG,
    Tile_X0Y1_E2BEGb,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6BEG,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4BEG,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_NN4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_SS4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W1END,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W2END,
    Tile_X0Y1_W2MID,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_W6END,
    Tile_X0Y1_WW4BEG,
    Tile_X0Y1_WW4END);
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 output [3:0] Tile_X0Y0_E1BEG;
 input [3:0] Tile_X0Y0_E1END;
 output [7:0] Tile_X0Y0_E2BEG;
 output [7:0] Tile_X0Y0_E2BEGb;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 output [11:0] Tile_X0Y0_E6BEG;
 input [11:0] Tile_X0Y0_E6END;
 output [15:0] Tile_X0Y0_EE4BEG;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 output [15:0] Tile_X0Y0_NN4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 input [15:0] Tile_X0Y0_SS4END;
 output [3:0] Tile_X0Y0_W1BEG;
 input [3:0] Tile_X0Y0_W1END;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 input [7:0] Tile_X0Y0_W2END;
 input [7:0] Tile_X0Y0_W2MID;
 output [11:0] Tile_X0Y0_W6BEG;
 input [11:0] Tile_X0Y0_W6END;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [15:0] Tile_X0Y0_WW4END;
 output [3:0] Tile_X0Y1_E1BEG;
 input [3:0] Tile_X0Y1_E1END;
 output [7:0] Tile_X0Y1_E2BEG;
 output [7:0] Tile_X0Y1_E2BEGb;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 output [11:0] Tile_X0Y1_E6BEG;
 input [11:0] Tile_X0Y1_E6END;
 output [15:0] Tile_X0Y1_EE4BEG;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 input [15:0] Tile_X0Y1_NN4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [15:0] Tile_X0Y1_SS4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 input [3:0] Tile_X0Y1_W1END;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 input [7:0] Tile_X0Y1_W2END;
 input [7:0] Tile_X0Y1_W2MID;
 output [11:0] Tile_X0Y1_W6BEG;
 input [11:0] Tile_X0Y1_W6END;
 output [15:0] Tile_X0Y1_WW4BEG;
 input [15:0] Tile_X0Y1_WW4END;

 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net750;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire \Tile_X0Y1_DSP_bot.A0 ;
 wire \Tile_X0Y1_DSP_bot.A1 ;
 wire \Tile_X0Y1_DSP_bot.A2 ;
 wire \Tile_X0Y1_DSP_bot.A3 ;
 wire \Tile_X0Y1_DSP_bot.B0 ;
 wire \Tile_X0Y1_DSP_bot.B1 ;
 wire \Tile_X0Y1_DSP_bot.B2 ;
 wire \Tile_X0Y1_DSP_bot.B3 ;
 wire \Tile_X0Y1_DSP_bot.C0 ;
 wire \Tile_X0Y1_DSP_bot.C1 ;
 wire \Tile_X0Y1_DSP_bot.C2 ;
 wire \Tile_X0Y1_DSP_bot.C3 ;
 wire \Tile_X0Y1_DSP_bot.C4 ;
 wire \Tile_X0Y1_DSP_bot.C5 ;
 wire \Tile_X0Y1_DSP_bot.C6 ;
 wire \Tile_X0Y1_DSP_bot.C7 ;
 wire \Tile_X0Y1_DSP_bot.C8 ;
 wire \Tile_X0Y1_DSP_bot.C9 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net707;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net723;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net691;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net665;
 wire net605;
 wire net713;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net616;
 wire net617;
 wire Tile_X0Y1_UserCLK_regs;
 wire clknet_0_Tile_X0Y1_UserCLK;
 wire clknet_1_0__leaf_Tile_X0Y1_UserCLK;
 wire clknet_0_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs;
 wire clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net657;
 wire net658;
 wire net662;
 wire net663;
 wire net664;
 wire net666;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net684;
 wire net688;
 wire net689;
 wire net690;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net714;
 wire net715;
 wire net716;
 wire net721;
 wire net722;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;

 sky130_fd_sc_hd__nor2_1 _1906_ (.A(_0740_),
    .B(_0829_),
    .Y(_0910_));
 sky130_fd_sc_hd__nor2_1 _1907_ (.A(_0450_),
    .B(_0601_),
    .Y(_0911_));
 sky130_fd_sc_hd__and3b_1 _1908_ (.A_N(_0601_),
    .B(_0575_),
    .C(_0574_),
    .X(_0912_));
 sky130_fd_sc_hd__xnor2_1 _1909_ (.A(_0889_),
    .B(_0911_),
    .Y(_0913_));
 sky130_fd_sc_hd__or3_1 _1910_ (.A(_0740_),
    .B(_0829_),
    .C(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__xnor2_1 _1911_ (.A(_0910_),
    .B(_0913_),
    .Y(_0915_));
 sky130_fd_sc_hd__a21o_1 _1912_ (.A1(_0909_),
    .A2(_0915_),
    .B1(_0908_),
    .X(_0916_));
 sky130_fd_sc_hd__xor2_1 _1913_ (.A(_0886_),
    .B(_0891_),
    .X(_0917_));
 sky130_fd_sc_hd__nand2_1 _1914_ (.A(_0916_),
    .B(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__xnor2_1 _1915_ (.A(_0916_),
    .B(_0917_),
    .Y(_0919_));
 sky130_fd_sc_hd__a21bo_1 _1916_ (.A1(_0889_),
    .A2(_0911_),
    .B1_N(_0914_),
    .X(_0920_));
 sky130_fd_sc_hd__mux4_2 _1917_ (.A0(net179),
    .A1(net125),
    .A2(net71),
    .A3(net233),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _1918_ (.A0(_0921_),
    .A1(_0173_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0922_));
 sky130_fd_sc_hd__mux4_2 _1919_ (.A0(net973),
    .A1(net968),
    .A2(net987),
    .A3(net992),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0923_));
 sky130_fd_sc_hd__or2_1 _1920_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .B(net983),
    .X(_0924_));
 sky130_fd_sc_hd__o211a_1 _1921_ (.A1(_0121_),
    .A2(net998),
    .B1(_0924_),
    .C1(_0122_),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _1922_ (.A0(net1019),
    .A1(net1015),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0926_));
 sky130_fd_sc_hd__a21o_1 _1923_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .A2(_0926_),
    .B1(_0123_),
    .X(_0927_));
 sky130_fd_sc_hd__o221a_1 _1924_ (.A1(_0923_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .B1(_0925_),
    .B2(_0927_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0928_));
 sky130_fd_sc_hd__a211o_1 _1925_ (.A1(_0323_),
    .A2(_0324_),
    .B1(_0121_),
    .C1(_0348_),
    .X(_0929_));
 sky130_fd_sc_hd__a211o_1 _1926_ (.A1(_0527_),
    .A2(_0528_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .C1(_0522_),
    .X(_0930_));
 sky130_fd_sc_hd__or2_1 _1927_ (.A(net74),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0931_));
 sky130_fd_sc_hd__o211a_1 _1928_ (.A1(net210),
    .A2(_0121_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .C1(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__a311o_1 _1929_ (.A1(_0929_),
    .A2(_0122_),
    .A3(_0930_),
    .B1(_0932_),
    .C1(_0123_),
    .X(_0933_));
 sky130_fd_sc_hd__mux4_1 _1930_ (.A0(net174),
    .A1(net182),
    .A2(net120),
    .A3(net128),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0934_));
 sky130_fd_sc_hd__o21ba_1 _1931_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0934_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0935_));
 sky130_fd_sc_hd__a21o_1 _1932_ (.A1(_0935_),
    .A2(_0933_),
    .B1(_0928_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__a211o_1 _1933_ (.A1(_0933_),
    .A2(_0935_),
    .B1(_0928_),
    .C1(_0120_),
    .X(_0936_));
 sky130_fd_sc_hd__o21a_1 _1934_ (.A1(net223),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .X(_0937_));
 sky130_fd_sc_hd__mux2_1 _1935_ (.A0(net187),
    .A1(net133),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0938_));
 sky130_fd_sc_hd__a221o_1 _1936_ (.A1(_0937_),
    .A2(_0936_),
    .B1(_0938_),
    .B2(_0124_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0939_));
 sky130_fd_sc_hd__mux4_2 _1937_ (.A0(net188),
    .A1(net134),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(net224),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0940_));
 sky130_fd_sc_hd__inv_2 _1938_ (.A(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__a21oi_2 _1939_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0941_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .Y(_0942_));
 sky130_fd_sc_hd__a22o_4 _1940_ (.A1(_0922_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .B1(_0939_),
    .B2(_0942_),
    .X(\Tile_X0Y1_DSP_bot.B1 ));
 sky130_fd_sc_hd__nand2b_1 _1941_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ),
    .B(net1061),
    .Y(_0943_));
 sky130_fd_sc_hd__o21ai_4 _1942_ (.A1(\Tile_X0Y1_DSP_bot.B1 ),
    .A2(net1061),
    .B1(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__nor2_4 _1943_ (.A(net626),
    .B(_0492_),
    .Y(_0945_));
 sky130_fd_sc_hd__nand2_2 _1944_ (.A(_0920_),
    .B(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__xnor2_1 _1945_ (.A(_0920_),
    .B(_0945_),
    .Y(_0947_));
 sky130_fd_sc_hd__o21ai_1 _1946_ (.A1(_0919_),
    .A2(_0947_),
    .B1(_0918_),
    .Y(_0948_));
 sky130_fd_sc_hd__xor2_1 _1947_ (.A(_0895_),
    .B(_0896_),
    .X(_0949_));
 sky130_fd_sc_hd__xor2_1 _1948_ (.A(_0948_),
    .B(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__a32oi_1 _1949_ (.A1(_0920_),
    .A2(_0945_),
    .A3(_0950_),
    .B1(_0949_),
    .B2(_0948_),
    .Y(_0951_));
 sky130_fd_sc_hd__and2b_1 _1950_ (.A_N(_0951_),
    .B(_0904_),
    .X(_0952_));
 sky130_fd_sc_hd__and2b_1 _1951_ (.A_N(_0904_),
    .B(_0951_),
    .X(_0953_));
 sky130_fd_sc_hd__nor2_1 _1952_ (.A(_0952_),
    .B(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__xnor2_2 _1953_ (.A(_0946_),
    .B(_0950_),
    .Y(_0955_));
 sky130_fd_sc_hd__o22ai_2 _1954_ (.A1(_0709_),
    .A2(_0785_),
    .B1(net624),
    .B2(_0661_),
    .Y(_0956_));
 sky130_fd_sc_hd__nand2_2 _1955_ (.A(_0906_),
    .B(_0956_),
    .Y(_0957_));
 sky130_fd_sc_hd__nor2_1 _1956_ (.A(net662),
    .B(_0829_),
    .Y(_0958_));
 sky130_fd_sc_hd__nor2_4 _1957_ (.A(_0676_),
    .B(_0450_),
    .Y(_0959_));
 sky130_fd_sc_hd__xor2_2 _1958_ (.A(_0912_),
    .B(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__xnor2_2 _1959_ (.A(_0960_),
    .B(_0958_),
    .Y(_0961_));
 sky130_fd_sc_hd__or2_1 _1960_ (.A(_0957_),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__xnor2_1 _1961_ (.A(_0909_),
    .B(_0915_),
    .Y(_0963_));
 sky130_fd_sc_hd__nor2_1 _1962_ (.A(_0962_),
    .B(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__xor2_1 _1963_ (.A(_0962_),
    .B(_0963_),
    .X(_0965_));
 sky130_fd_sc_hd__a22o_1 _1964_ (.A1(_0912_),
    .A2(_0959_),
    .B1(_0960_),
    .B2(_0958_),
    .X(_0966_));
 sky130_fd_sc_hd__mux4_2 _1965_ (.A0(net126),
    .A1(net233),
    .A2(net92),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_0967_));
 sky130_fd_sc_hd__mux4_1 _1966_ (.A0(net204),
    .A1(net129),
    .A2(net75),
    .A3(net219),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_4 _1967_ (.A0(_0968_),
    .A1(_0967_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .X(_0969_));
 sky130_fd_sc_hd__a211o_1 _1968_ (.A1(_0533_),
    .A2(_0535_),
    .B1(_0125_),
    .C1(_0507_),
    .X(_0970_));
 sky130_fd_sc_hd__o21a_1 _1969_ (.A1(net227),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_1 _1970_ (.A0(net137),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_0972_));
 sky130_fd_sc_hd__a221o_1 _1971_ (.A1(_0970_),
    .A2(_0971_),
    .B1(_0972_),
    .B2(_0126_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_4 _1972_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .A1(net228),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0974_));
 sky130_fd_sc_hd__nand2_1 _1973_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__mux2_1 _1974_ (.A0(net192),
    .A1(net138),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0976_));
 sky130_fd_sc_hd__inv_1 _1975_ (.A(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__o211a_1 _1976_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .A2(_0977_),
    .B1(_0975_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .X(_0978_));
 sky130_fd_sc_hd__nor2_1 _1977_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__a22o_4 _1978_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0969_),
    .B1(_0979_),
    .B2(_0973_),
    .X(\Tile_X0Y1_DSP_bot.B0 ));
 sky130_fd_sc_hd__nand2b_1 _1979_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ),
    .B(net1061),
    .Y(_0980_));
 sky130_fd_sc_hd__o21ai_4 _1980_ (.A1(\Tile_X0Y1_DSP_bot.B0 ),
    .A2(net1061),
    .B1(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__nor2_1 _1981_ (.A(_0492_),
    .B(net625),
    .Y(_0982_));
 sky130_fd_sc_hd__xnor2_1 _1982_ (.A(_0966_),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__o21ai_1 _1983_ (.A1(net722),
    .A2(_0944_),
    .B1(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__or3_1 _1984_ (.A(net722),
    .B(net626),
    .C(_0983_),
    .X(_0985_));
 sky130_fd_sc_hd__and2_1 _1985_ (.A(_0984_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__a21o_1 _1986_ (.A1(_0965_),
    .A2(_0986_),
    .B1(_0964_),
    .X(_0987_));
 sky130_fd_sc_hd__xor2_1 _1987_ (.A(_0919_),
    .B(_0947_),
    .X(_0988_));
 sky130_fd_sc_hd__and2_1 _1988_ (.A(_0987_),
    .B(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__a21bo_1 _1989_ (.A1(_0966_),
    .A2(_0982_),
    .B1_N(_0985_),
    .X(_0990_));
 sky130_fd_sc_hd__xor2_1 _1990_ (.A(_0987_),
    .B(_0988_),
    .X(_0991_));
 sky130_fd_sc_hd__a21oi_1 _1991_ (.A1(_0990_),
    .A2(_0991_),
    .B1(_0989_),
    .Y(_0992_));
 sky130_fd_sc_hd__and2b_1 _1992_ (.A_N(_0992_),
    .B(_0955_),
    .X(_0993_));
 sky130_fd_sc_hd__xnor2_2 _1993_ (.A(_0955_),
    .B(_0992_),
    .Y(_0994_));
 sky130_fd_sc_hd__xor2_1 _1994_ (.A(_0990_),
    .B(_0991_),
    .X(_0995_));
 sky130_fd_sc_hd__xor2_2 _1995_ (.A(_0957_),
    .B(_0961_),
    .X(_0996_));
 sky130_fd_sc_hd__nor2_1 _1996_ (.A(_0601_),
    .B(_0829_),
    .Y(_0997_));
 sky130_fd_sc_hd__nor2_1 _1997_ (.A(_0450_),
    .B(_0785_),
    .Y(_0998_));
 sky130_fd_sc_hd__a31oi_4 _1998_ (.A1(_0677_),
    .A2(_0575_),
    .A3(_0574_),
    .B1(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__and3_4 _1999_ (.A(_0784_),
    .B(_0575_),
    .C(_0574_),
    .X(_1000_));
 sky130_fd_sc_hd__nand2_4 _2000_ (.A(_0959_),
    .B(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__a21o_1 _2001_ (.A1(_0959_),
    .A2(_1000_),
    .B1(_0999_),
    .X(_1002_));
 sky130_fd_sc_hd__xor2_4 _2002_ (.A(_0997_),
    .B(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__or3_4 _2003_ (.A(_1003_),
    .B(net624),
    .C(net665),
    .X(_1004_));
 sky130_fd_sc_hd__inv_1 _2004_ (.A(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__xor2_4 _2005_ (.A(_0996_),
    .B(_1004_),
    .X(_1006_));
 sky130_fd_sc_hd__or2_1 _2006_ (.A(_0740_),
    .B(net626),
    .X(_1007_));
 sky130_fd_sc_hd__o31ai_4 _2007_ (.A1(_0601_),
    .A2(_0829_),
    .A3(_0999_),
    .B1(_1001_),
    .Y(_1008_));
 sky130_fd_sc_hd__nor2_8 _2008_ (.A(net625),
    .B(net722),
    .Y(_1009_));
 sky130_fd_sc_hd__xnor2_4 _2009_ (.A(_1009_),
    .B(_1008_),
    .Y(_1010_));
 sky130_fd_sc_hd__xnor2_4 _2010_ (.A(_1010_),
    .B(_1007_),
    .Y(_1011_));
 sky130_fd_sc_hd__nor2_1 _2011_ (.A(_1011_),
    .B(_1006_),
    .Y(_1012_));
 sky130_fd_sc_hd__a21o_1 _2012_ (.A1(_0996_),
    .A2(_1005_),
    .B1(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__xnor2_2 _2013_ (.A(_0965_),
    .B(_0986_),
    .Y(_1014_));
 sky130_fd_sc_hd__and2b_1 _2014_ (.A_N(_1014_),
    .B(_1013_),
    .X(_1015_));
 sky130_fd_sc_hd__a2bb2o_4 _2015_ (.A1_N(_1007_),
    .A2_N(_1010_),
    .B1(_1008_),
    .B2(_1009_),
    .X(_1016_));
 sky130_fd_sc_hd__xnor2_2 _2016_ (.A(_1013_),
    .B(_1014_),
    .Y(_1017_));
 sky130_fd_sc_hd__a21oi_2 _2017_ (.A1(_1016_),
    .A2(_1017_),
    .B1(_1015_),
    .Y(_1018_));
 sky130_fd_sc_hd__and2b_1 _2018_ (.A_N(_1018_),
    .B(_0995_),
    .X(_1019_));
 sky130_fd_sc_hd__xnor2_1 _2019_ (.A(_0995_),
    .B(_1018_),
    .Y(_1020_));
 sky130_fd_sc_hd__xor2_4 _2020_ (.A(_1016_),
    .B(_1017_),
    .X(_1021_));
 sky130_fd_sc_hd__xor2_4 _2021_ (.A(_1003_),
    .B(_0905_),
    .X(_1022_));
 sky130_fd_sc_hd__or2_4 _2022_ (.A(_0729_),
    .B(net626),
    .X(_1023_));
 sky130_fd_sc_hd__and3b_1 _2023_ (.A_N(net624),
    .B(_0575_),
    .C(_0574_),
    .X(_1024_));
 sky130_fd_sc_hd__nor2_1 _2024_ (.A(_0450_),
    .B(net624),
    .Y(_1025_));
 sky130_fd_sc_hd__and3_1 _2025_ (.A(_0827_),
    .B(_0677_),
    .C(_0828_),
    .X(_1026_));
 sky130_fd_sc_hd__a31o_1 _2026_ (.A1(_0574_),
    .A2(_0575_),
    .A3(_0784_),
    .B1(_1025_),
    .X(_1027_));
 sky130_fd_sc_hd__a21bo_1 _2027_ (.A1(_0998_),
    .A2(_1024_),
    .B1_N(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__a22o_4 _2028_ (.A1(_0998_),
    .A2(_1024_),
    .B1(_1027_),
    .B2(_1026_),
    .X(_1029_));
 sky130_fd_sc_hd__nor2_1 _2029_ (.A(_0740_),
    .B(net625),
    .Y(_1030_));
 sky130_fd_sc_hd__xnor2_4 _2030_ (.A(_1030_),
    .B(_1029_),
    .Y(_1031_));
 sky130_fd_sc_hd__xnor2_4 _2031_ (.A(_1023_),
    .B(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__nor2_8 _2032_ (.A(_1022_),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__xor2_4 _2033_ (.A(_1011_),
    .B(_1006_),
    .X(_1034_));
 sky130_fd_sc_hd__nand2_4 _2034_ (.A(_1033_),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__o2bb2a_4 _2035_ (.A1_N(_1029_),
    .A2_N(_1030_),
    .B1(_1031_),
    .B2(_1023_),
    .X(_1036_));
 sky130_fd_sc_hd__xnor2_4 _2036_ (.A(_1034_),
    .B(_1033_),
    .Y(_1037_));
 sky130_fd_sc_hd__o21ai_4 _2037_ (.A1(_1036_),
    .A2(_1037_),
    .B1(_1035_),
    .Y(_1038_));
 sky130_fd_sc_hd__or2_4 _2038_ (.A(_1038_),
    .B(_1021_),
    .X(_1039_));
 sky130_fd_sc_hd__xnor2_4 _2039_ (.A(_1037_),
    .B(_1036_),
    .Y(_1040_));
 sky130_fd_sc_hd__xor2_2 _2040_ (.A(_1022_),
    .B(_1032_),
    .X(_1041_));
 sky130_fd_sc_hd__xnor2_1 _2041_ (.A(_1026_),
    .B(_1028_),
    .Y(_1042_));
 sky130_fd_sc_hd__nor2_1 _2042_ (.A(_0601_),
    .B(_0944_),
    .Y(_1043_));
 sky130_fd_sc_hd__and3b_2 _2043_ (.A_N(_0878_),
    .B(_0828_),
    .C(_0827_),
    .X(_1044_));
 sky130_fd_sc_hd__a2bb2o_1 _2044_ (.A1_N(net662),
    .A2_N(_0981_),
    .B1(_1000_),
    .B2(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__or4bb_1 _2045_ (.A(net662),
    .B(net625),
    .C_N(_1000_),
    .D_N(_1044_),
    .X(_1046_));
 sky130_fd_sc_hd__a21o_1 _2046_ (.A1(_1045_),
    .A2(_1046_),
    .B1(_1043_),
    .X(_1047_));
 sky130_fd_sc_hd__nand3_1 _2047_ (.A(_1043_),
    .B(_1045_),
    .C(_1046_),
    .Y(_1048_));
 sky130_fd_sc_hd__and3_4 _2048_ (.A(_1042_),
    .B(_1047_),
    .C(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__nand2_1 _2049_ (.A(_1046_),
    .B(_1048_),
    .Y(_1050_));
 sky130_fd_sc_hd__xnor2_2 _2050_ (.A(_1049_),
    .B(_1041_),
    .Y(_1051_));
 sky130_fd_sc_hd__and2b_1 _2051_ (.A_N(_1051_),
    .B(_1050_),
    .X(_1052_));
 sky130_fd_sc_hd__a21o_1 _2052_ (.A1(_1041_),
    .A2(_1049_),
    .B1(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__and2b_1 _2053_ (.A_N(_1040_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__xnor2_4 _2054_ (.A(_1053_),
    .B(_1040_),
    .Y(_1055_));
 sky130_fd_sc_hd__xor2_1 _2055_ (.A(_1051_),
    .B(_1050_),
    .X(_1056_));
 sky130_fd_sc_hd__o21ba_1 _2056_ (.A1(_0785_),
    .A2(_0829_),
    .B1_N(_1024_),
    .X(_1057_));
 sky130_fd_sc_hd__a21o_1 _2057_ (.A1(_1000_),
    .A2(_1044_),
    .B1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__nor2_4 _2058_ (.A(_0981_),
    .B(_0676_),
    .Y(_1059_));
 sky130_fd_sc_hd__nand2_2 _2059_ (.A(_1043_),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__o22a_1 _2060_ (.A1(_0676_),
    .A2(_0944_),
    .B1(net625),
    .B2(_0601_),
    .X(_1061_));
 sky130_fd_sc_hd__a21o_1 _2061_ (.A1(_1043_),
    .A2(_1059_),
    .B1(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__nor2_1 _2062_ (.A(_1062_),
    .B(_1058_),
    .Y(_1063_));
 sky130_fd_sc_hd__a21oi_1 _2063_ (.A1(_1047_),
    .A2(_1048_),
    .B1(_1042_),
    .Y(_1064_));
 sky130_fd_sc_hd__or3b_4 _2064_ (.A(_1049_),
    .B(_1064_),
    .C_N(_1063_),
    .X(_1065_));
 sky130_fd_sc_hd__o21bai_1 _2065_ (.A1(_1049_),
    .A2(_1064_),
    .B1_N(_1063_),
    .Y(_1066_));
 sky130_fd_sc_hd__nand3b_4 _2066_ (.A_N(_1060_),
    .B(_1065_),
    .C(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__and2_4 _2067_ (.A(_1067_),
    .B(_1065_),
    .X(_1068_));
 sky130_fd_sc_hd__nor2_1 _2068_ (.A(_1056_),
    .B(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__xor2_4 _2069_ (.A(_1068_),
    .B(_1056_),
    .X(_1070_));
 sky130_fd_sc_hd__a21bo_1 _2070_ (.A1(_1065_),
    .A2(_1066_),
    .B1_N(_1060_),
    .X(_1071_));
 sky130_fd_sc_hd__xor2_1 _2071_ (.A(_1058_),
    .B(_1062_),
    .X(_1072_));
 sky130_fd_sc_hd__nor2_1 _2072_ (.A(_0785_),
    .B(_0944_),
    .Y(_1073_));
 sky130_fd_sc_hd__and2_1 _2073_ (.A(_1059_),
    .B(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__xor2_2 _2074_ (.A(_1059_),
    .B(_1073_),
    .X(_1075_));
 sky130_fd_sc_hd__and2_1 _2075_ (.A(_1044_),
    .B(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__xnor2_1 _2076_ (.A(_1072_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__o21a_1 _2077_ (.A1(_1074_),
    .A2(_1076_),
    .B1(_1072_),
    .X(_1078_));
 sky130_fd_sc_hd__nand3_4 _2078_ (.A(_1071_),
    .B(_1067_),
    .C(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__xnor2_1 _2079_ (.A(_1074_),
    .B(_1077_),
    .Y(_1080_));
 sky130_fd_sc_hd__nor2_4 _2080_ (.A(_0878_),
    .B(_0981_),
    .Y(_1081_));
 sky130_fd_sc_hd__nand2_4 _2081_ (.A(_1073_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__xnor2_4 _2082_ (.A(_1075_),
    .B(_1044_),
    .Y(_1083_));
 sky130_fd_sc_hd__nor2_1 _2083_ (.A(_1082_),
    .B(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__and2_1 _2084_ (.A(_1080_),
    .B(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__a21o_1 _2085_ (.A1(_1067_),
    .A2(_1071_),
    .B1(_1078_),
    .X(_1086_));
 sky130_fd_sc_hd__nand3_4 _2086_ (.A(_1079_),
    .B(_1085_),
    .C(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__a21bo_1 _2087_ (.A1(_1085_),
    .A2(_1086_),
    .B1_N(_1079_),
    .X(_1088_));
 sky130_fd_sc_hd__a21o_1 _2088_ (.A1(_1070_),
    .A2(_1088_),
    .B1(_1069_),
    .X(_1089_));
 sky130_fd_sc_hd__a21o_1 _2089_ (.A1(_1055_),
    .A2(_1089_),
    .B1(_1054_),
    .X(_1090_));
 sky130_fd_sc_hd__a221o_1 _2090_ (.A1(_1021_),
    .A2(_1038_),
    .B1(_1055_),
    .B2(_1089_),
    .C1(_1054_),
    .X(_1091_));
 sky130_fd_sc_hd__xor2_2 _2091_ (.A(_1021_),
    .B(_1038_),
    .X(_1092_));
 sky130_fd_sc_hd__and3_1 _2092_ (.A(_1020_),
    .B(_1091_),
    .C(_1039_),
    .X(_1093_));
 sky130_fd_sc_hd__a31o_1 _2093_ (.A1(_1020_),
    .A2(_1039_),
    .A3(_1091_),
    .B1(_1019_),
    .X(_1094_));
 sky130_fd_sc_hd__a21o_1 _2094_ (.A1(_0994_),
    .A2(_1094_),
    .B1(_0993_),
    .X(_1095_));
 sky130_fd_sc_hd__a21o_1 _2095_ (.A1(_1095_),
    .A2(_0954_),
    .B1(_0952_),
    .X(_1096_));
 sky130_fd_sc_hd__a21o_1 _2096_ (.A1(_0903_),
    .A2(_1096_),
    .B1(_0901_),
    .X(_1097_));
 sky130_fd_sc_hd__nand2_4 _2097_ (.A(_0841_),
    .B(_0858_),
    .Y(_1098_));
 sky130_fd_sc_hd__nand2b_1 _2098_ (.A_N(_0859_),
    .B(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__a21o_4 _2099_ (.A1(_1097_),
    .A2(_1098_),
    .B1(_0859_),
    .X(_1100_));
 sky130_fd_sc_hd__nor2_1 _2100_ (.A(_0854_),
    .B(_0857_),
    .Y(_1101_));
 sky130_fd_sc_hd__o22ai_2 _2101_ (.A1(net722),
    .A2(_0620_),
    .B1(_0661_),
    .B2(_0492_),
    .Y(_1102_));
 sky130_fd_sc_hd__or2_1 _2102_ (.A(_0492_),
    .B(_0620_),
    .X(_1103_));
 sky130_fd_sc_hd__o31ai_2 _2103_ (.A1(_1103_),
    .A2(_0661_),
    .A3(net722),
    .B1(_1102_),
    .Y(_1104_));
 sky130_fd_sc_hd__o21ba_4 _2104_ (.A1(_0845_),
    .A2(_0848_),
    .B1_N(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__nor3b_1 _2105_ (.A(_0845_),
    .B(_0848_),
    .C_N(_1104_),
    .Y(_1106_));
 sky130_fd_sc_hd__inv_1 _2106_ (.A(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__or2_1 _2107_ (.A(_1105_),
    .B(_1106_),
    .X(_1108_));
 sky130_fd_sc_hd__xnor2_4 _2108_ (.A(_1108_),
    .B(_0851_),
    .Y(_1109_));
 sky130_fd_sc_hd__xnor2_4 _2109_ (.A(_1109_),
    .B(_1101_),
    .Y(_1110_));
 sky130_fd_sc_hd__a22oi_4 _2110_ (.A1(_0857_),
    .A2(_1109_),
    .B1(_1110_),
    .B2(_1100_),
    .Y(_1111_));
 sky130_fd_sc_hd__nor2_1 _2111_ (.A(_0843_),
    .B(_1103_),
    .Y(_1112_));
 sky130_fd_sc_hd__o31a_1 _2112_ (.A1(_0851_),
    .A2(_1105_),
    .A3(_0854_),
    .B1(_1107_),
    .X(_1113_));
 sky130_fd_sc_hd__xnor2_2 _2113_ (.A(_1113_),
    .B(_1112_),
    .Y(_1114_));
 sky130_fd_sc_hd__or2_4 _2114_ (.A(_1111_),
    .B(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__xnor2_2 _2115_ (.A(_1111_),
    .B(_1114_),
    .Y(_1116_));
 sky130_fd_sc_hd__nand2b_4 _2116_ (.A_N(_1116_),
    .B(_0432_),
    .Y(_1117_));
 sky130_fd_sc_hd__xor2_1 _2117_ (.A(_0432_),
    .B(_1116_),
    .X(_1118_));
 sky130_fd_sc_hd__nand2_1 _2118_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ),
    .Y(_1119_));
 sky130_fd_sc_hd__mux4_1 _2119_ (.A0(net1011),
    .A1(net1046),
    .A2(net1028),
    .A3(net1052),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_1120_));
 sky130_fd_sc_hd__mux4_1 _2120_ (.A0(net1042),
    .A1(net1033),
    .A2(net1007),
    .A3(net1054),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_1121_));
 sky130_fd_sc_hd__mux2_1 _2121_ (.A0(_1120_),
    .A1(_1121_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_1122_));
 sky130_fd_sc_hd__or2_1 _2122_ (.A(_0089_),
    .B(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__mux4_2 _2123_ (.A0(net619),
    .A1(net1258),
    .A2(net191),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_1124_));
 sky130_fd_sc_hd__mux4_1 _2124_ (.A0(net57),
    .A1(net59),
    .A2(net67),
    .A3(net95),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_1125_));
 sky130_fd_sc_hd__mux2_4 _2125_ (.A0(_1124_),
    .A1(_1125_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_1126_));
 sky130_fd_sc_hd__o21ai_4 _2126_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ),
    .A2(_1126_),
    .B1(_1123_),
    .Y(_1127_));
 sky130_fd_sc_hd__inv_1 _2127_ (.A(_1127_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ));
 sky130_fd_sc_hd__nand2_2 _2128_ (.A(_1127_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ),
    .Y(_1128_));
 sky130_fd_sc_hd__o21a_1 _2129_ (.A1(net105),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ),
    .X(_1129_));
 sky130_fd_sc_hd__mux2_1 _2130_ (.A0(net13),
    .A1(net69),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_1130_));
 sky130_fd_sc_hd__a221o_1 _2131_ (.A1(_1129_),
    .A2(_1128_),
    .B1(_1130_),
    .B2(_0090_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_1131_));
 sky130_fd_sc_hd__mux2_2 _2132_ (.A0(net690),
    .A1(net14),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_1132_));
 sky130_fd_sc_hd__inv_1 _2133_ (.A(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__mux2_1 _2134_ (.A0(net70),
    .A1(net106),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_1134_));
 sky130_fd_sc_hd__nand2_1 _2135_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ),
    .B(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hd__o211a_1 _2136_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ),
    .A2(_1133_),
    .B1(_1135_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_1136_));
 sky130_fd_sc_hd__nor2_1 _2137_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__mux4_2 _2138_ (.A0(net26),
    .A1(net116),
    .A2(net77),
    .A3(_0468_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_1138_));
 sky130_fd_sc_hd__mux4_2 _2139_ (.A0(net207),
    .A1(net6),
    .A2(net62),
    .A3(net98),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_4 _2140_ (.A0(_1139_),
    .A1(_1138_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_1140_));
 sky130_fd_sc_hd__a22o_1 _2141_ (.A1(_1137_),
    .A2(_1131_),
    .B1(_1140_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ));
 sky130_fd_sc_hd__mux2_4 _2142_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .X(_1141_));
 sky130_fd_sc_hd__nand2_4 _2143_ (.A(net1058),
    .B(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__xnor2_4 _2144_ (.A(_1110_),
    .B(_1100_),
    .Y(_1143_));
 sky130_fd_sc_hd__nand3_4 _2145_ (.A(_1143_),
    .B(_1142_),
    .C(_1119_),
    .Y(_1144_));
 sky130_fd_sc_hd__inv_2 _2146_ (.A(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__a21oi_4 _2147_ (.A1(_1119_),
    .A2(_1142_),
    .B1(_1143_),
    .Y(_1146_));
 sky130_fd_sc_hd__mux4_2 _2148_ (.A0(net190),
    .A1(net86),
    .A2(net10),
    .A3(net102),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_1 _2149_ (.A0(_1147_),
    .A1(_0520_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_1148_));
 sky130_fd_sc_hd__mux4_2 _2150_ (.A0(_0536_),
    .A1(_0081_),
    .A2(_0030_),
    .A3(_0158_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1149_));
 sky130_fd_sc_hd__mux4_2 _2151_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .A1(net109),
    .A2(net73),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1150_));
 sky130_fd_sc_hd__mux4_2 _2152_ (.A0(net710),
    .A1(net74),
    .A2(net18),
    .A3(net110),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_4 _2153_ (.A0(_1150_),
    .A1(_1151_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_1152_));
 sky130_fd_sc_hd__mux2_4 _2154_ (.A0(_1152_),
    .A1(_1148_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ));
 sky130_fd_sc_hd__mux2_2 _2155_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_4 _2156_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ),
    .A1(_1153_),
    .S(net1058),
    .X(_1154_));
 sky130_fd_sc_hd__xnor2_2 _2157_ (.A(_1097_),
    .B(_1099_),
    .Y(_1155_));
 sky130_fd_sc_hd__and2_1 _2158_ (.A(_1154_),
    .B(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__xor2_2 _2159_ (.A(_1154_),
    .B(_1155_),
    .X(_1157_));
 sky130_fd_sc_hd__mux4_2 _2160_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net16),
    .A2(net72),
    .A3(net108),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_1158_));
 sky130_fd_sc_hd__mux4_1 _2161_ (.A0(net1012),
    .A1(net1047),
    .A2(net1027),
    .A3(net1051),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1159_));
 sky130_fd_sc_hd__and2b_1 _2162_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__mux4_1 _2163_ (.A0(net1043),
    .A1(net1032),
    .A2(net1008),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_1161_));
 sky130_fd_sc_hd__a21bo_1 _2164_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_1161_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_1162_));
 sky130_fd_sc_hd__mux4_1 _2165_ (.A0(net620),
    .A1(net1258),
    .A2(net191),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_1163_));
 sky130_fd_sc_hd__mux4_1 _2166_ (.A0(net57),
    .A1(net59),
    .A2(net67),
    .A3(net1220),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_2 _2167_ (.A0(_1163_),
    .A1(_1164_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_1165_));
 sky130_fd_sc_hd__o22a_4 _2168_ (.A1(_1160_),
    .A2(_1162_),
    .B1(_1165_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _2169_ (.A0(net188),
    .A1(net8),
    .A2(net64),
    .A3(net116),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_1166_));
 sky130_fd_sc_hd__mux4_1 _2170_ (.A0(net207),
    .A1(net79),
    .A2(net7),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1167_));
 sky130_fd_sc_hd__mux4_1 _2171_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A1(net15),
    .A2(net71),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_1168_));
 sky130_fd_sc_hd__mux4_2 _2172_ (.A0(_1168_),
    .A1(_1166_),
    .A2(_1158_),
    .A3(_1167_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ));
 sky130_fd_sc_hd__mux2_1 _2173_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ),
    .S(net1064),
    .X(_1169_));
 sky130_fd_sc_hd__mux2_1 _2174_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ),
    .A1(_1169_),
    .S(net1058),
    .X(_1170_));
 sky130_fd_sc_hd__xnor2_2 _2175_ (.A(_0903_),
    .B(_1096_),
    .Y(_1171_));
 sky130_fd_sc_hd__and2b_1 _2176_ (.A_N(_1171_),
    .B(_1170_),
    .X(_1172_));
 sky130_fd_sc_hd__nand2b_1 _2177_ (.A_N(_1170_),
    .B(_1171_),
    .Y(_1173_));
 sky130_fd_sc_hd__nand2b_4 _2178_ (.A_N(_1172_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__mux4_2 _2179_ (.A0(net200),
    .A1(net8),
    .A2(net100),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_1175_));
 sky130_fd_sc_hd__mux4_2 _2180_ (.A0(net192),
    .A1(net25),
    .A2(net68),
    .A3(net104),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_1176_));
 sky130_fd_sc_hd__mux2_4 _2181_ (.A0(_1176_),
    .A1(_1175_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_1177_));
 sky130_fd_sc_hd__mux4_1 _2182_ (.A0(net1012),
    .A1(net1048),
    .A2(net1027),
    .A3(net1052),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_1178_));
 sky130_fd_sc_hd__nand2b_1 _2183_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .B(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hd__mux4_1 _2184_ (.A0(net1043),
    .A1(net1032),
    .A2(net1008),
    .A3(net1022),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_1180_));
 sky130_fd_sc_hd__nand2_1 _2185_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .B(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__mux4_1 _2186_ (.A0(net619),
    .A1(net3),
    .A2(net191),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_1182_));
 sky130_fd_sc_hd__mux4_1 _2187_ (.A0(net59),
    .A1(net67),
    .A2(net93),
    .A3(net1220),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(_1182_),
    .A1(_1183_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_1184_));
 sky130_fd_sc_hd__nor2_1 _2189_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__a31o_1 _2190_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ),
    .A2(_1179_),
    .A3(_1181_),
    .B1(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__inv_2 _2191_ (.A(_1186_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _2192_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .A1(net19),
    .A2(net111),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ),
    .X(_1187_));
 sky130_fd_sc_hd__mux2_1 _2193_ (.A0(_1187_),
    .A1(_0526_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_1188_));
 sky130_fd_sc_hd__mux2_4 _2194_ (.A0(_1188_),
    .A1(_1177_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ));
 sky130_fd_sc_hd__mux2_4 _2195_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ),
    .S(net1064),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_4 _2196_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ),
    .A1(_1189_),
    .S(net1058),
    .X(_1190_));
 sky130_fd_sc_hd__xnor2_1 _2197_ (.A(_0954_),
    .B(_1095_),
    .Y(_1191_));
 sky130_fd_sc_hd__and2b_1 _2198_ (.A_N(_1191_),
    .B(_1190_),
    .X(_1192_));
 sky130_fd_sc_hd__xnor2_1 _2199_ (.A(_1190_),
    .B(_1191_),
    .Y(_1193_));
 sky130_fd_sc_hd__and2_1 _2200_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ),
    .X(_1194_));
 sky130_fd_sc_hd__mux4_1 _2201_ (.A0(net974),
    .A1(net970),
    .A2(net989),
    .A3(net994),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1195_));
 sky130_fd_sc_hd__inv_1 _2202_ (.A(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__mux2_1 _2203_ (.A0(net979),
    .A1(net998),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_1197_));
 sky130_fd_sc_hd__and2b_1 _2204_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .B(net734),
    .X(_1198_));
 sky130_fd_sc_hd__a21bo_1 _2205_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .A2(net693),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1199_));
 sky130_fd_sc_hd__o221a_1 _2206_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .A2(_1197_),
    .B1(_1198_),
    .B2(_1199_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_1200_));
 sky130_fd_sc_hd__o21ai_1 _2207_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_1196_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .Y(_1201_));
 sky130_fd_sc_hd__mux4_2 _2208_ (.A0(_0410_),
    .A1(_0302_),
    .A2(net75),
    .A3(net1068),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1202_));
 sky130_fd_sc_hd__mux4_1 _2209_ (.A0(net175),
    .A1(net121),
    .A2(net183),
    .A3(net129),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_1203_));
 sky130_fd_sc_hd__and2b_1 _2210_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .B(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__a211o_1 _2211_ (.A1(_1202_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .B1(_1204_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_1205_));
 sky130_fd_sc_hd__o21a_1 _2212_ (.A1(_1200_),
    .A2(_1201_),
    .B1(_1205_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__mux2_2 _2213_ (.A0(_0410_),
    .A1(_0302_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1206_));
 sky130_fd_sc_hd__nand2b_1 _2214_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__mux2_1 _2215_ (.A0(net89),
    .A1(net231),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1208_));
 sky130_fd_sc_hd__nand2_1 _2216_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__mux4_1 _2217_ (.A0(net173),
    .A1(net177),
    .A2(net119),
    .A3(net123),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1210_));
 sky130_fd_sc_hd__nor2_1 _2218_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .B(_1210_),
    .Y(_1211_));
 sky130_fd_sc_hd__a311oi_1 _2219_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_1207_),
    .A3(_1209_),
    .B1(_1211_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .Y(_1212_));
 sky130_fd_sc_hd__mux2_1 _2220_ (.A0(net979),
    .A1(net984),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1213_));
 sky130_fd_sc_hd__inv_1 _2221_ (.A(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__mux2_1 _2222_ (.A0(net997),
    .A1(net693),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1215_));
 sky130_fd_sc_hd__o21ai_1 _2223_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .A2(_1214_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .Y(_1216_));
 sky130_fd_sc_hd__a21o_1 _2224_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .A2(_1215_),
    .B1(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__nand2b_1 _2225_ (.A_N(net968),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .Y(_1218_));
 sky130_fd_sc_hd__o21ba_1 _2226_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(net973),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1219_));
 sky130_fd_sc_hd__mux2_1 _2227_ (.A0(net987),
    .A1(net992),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1220_));
 sky130_fd_sc_hd__a221o_1 _2228_ (.A1(_1218_),
    .A2(_1219_),
    .B1(_1220_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1221_));
 sky130_fd_sc_hd__a31o_1 _2229_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1217_),
    .A3(_1221_),
    .B1(_1212_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(_0410_),
    .A1(_0302_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_1222_));
 sky130_fd_sc_hd__and2b_1 _2231_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .B(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(net75),
    .A1(net1068),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_1224_));
 sky130_fd_sc_hd__a21o_1 _2233_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .A2(_1224_),
    .B1(_0131_),
    .X(_1225_));
 sky130_fd_sc_hd__mux4_1 _2234_ (.A0(net175),
    .A1(net1218),
    .A2(net183),
    .A3(net129),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_1226_));
 sky130_fd_sc_hd__o221a_1 _2235_ (.A1(_1223_),
    .A2(_1225_),
    .B1(_1226_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .C1(_0132_),
    .X(_1227_));
 sky130_fd_sc_hd__mux4_1 _2236_ (.A0(net978),
    .A1(net998),
    .A2(net1019),
    .A3(net1002),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_1228_));
 sky130_fd_sc_hd__or2_1 _2237_ (.A(_0131_),
    .B(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__mux4_1 _2238_ (.A0(net973),
    .A1(net968),
    .A2(net987),
    .A3(net992),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_1230_));
 sky130_fd_sc_hd__or2_1 _2239_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .B(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__a31o_4 _2240_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .A2(_1229_),
    .A3(_1231_),
    .B1(_1227_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ));
 sky130_fd_sc_hd__mux2_1 _2241_ (.A0(_0410_),
    .A1(_0302_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_1 _2242_ (.A0(net69),
    .A1(net209),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1233_));
 sky130_fd_sc_hd__a21bo_1 _2243_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .A2(_1233_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .X(_1234_));
 sky130_fd_sc_hd__a21o_1 _2244_ (.A1(_0133_),
    .A2(_1232_),
    .B1(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__mux4_1 _2245_ (.A0(net173),
    .A1(net177),
    .A2(net119),
    .A3(net123),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1236_));
 sky130_fd_sc_hd__o21ba_1 _2246_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(_1236_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_1237_));
 sky130_fd_sc_hd__mux4_1 _2247_ (.A0(net973),
    .A1(net968),
    .A2(net987),
    .A3(net992),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1238_));
 sky130_fd_sc_hd__mux4_1 _2248_ (.A0(net979),
    .A1(net998),
    .A2(net984),
    .A3(net1002),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _2249_ (.A0(_1238_),
    .A1(_1239_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .X(_1240_));
 sky130_fd_sc_hd__a22o_1 _2250_ (.A1(_1235_),
    .A2(_1237_),
    .B1(_1240_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_1241_));
 sky130_fd_sc_hd__mux4_2 _2251_ (.A0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .A3(_1241_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1242_));
 sky130_fd_sc_hd__nand2_1 _2252_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .B(_0425_),
    .Y(_1243_));
 sky130_fd_sc_hd__o21ai_1 _2253_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .B1(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__mux4_1 _2254_ (.A0(net974),
    .A1(net969),
    .A2(net988),
    .A3(net993),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_1245_));
 sky130_fd_sc_hd__mux4_1 _2255_ (.A0(net978),
    .A1(net997),
    .A2(net983),
    .A3(net1014),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_1246_));
 sky130_fd_sc_hd__o21a_1 _2256_ (.A1(_0130_),
    .A2(_1246_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_1247_));
 sky130_fd_sc_hd__o21ai_1 _2257_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(_1245_),
    .B1(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__mux2_2 _2258_ (.A0(_0410_),
    .A1(net69),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_1249_));
 sky130_fd_sc_hd__inv_1 _2259_ (.A(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__mux2_1 _2260_ (.A0(net209),
    .A1(net211),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_1251_));
 sky130_fd_sc_hd__nand2_1 _2261_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .B(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__o211a_1 _2262_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_1250_),
    .B1(_1252_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_1253_));
 sky130_fd_sc_hd__mux4_1 _2263_ (.A0(net173),
    .A1(net177),
    .A2(net119),
    .A3(net123),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_1254_));
 sky130_fd_sc_hd__nor2_1 _2264_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .B(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__o31ai_2 _2265_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_1253_),
    .A3(_1255_),
    .B1(_1248_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ));
 sky130_fd_sc_hd__nor2_1 _2266_ (.A(_0127_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ),
    .Y(_1256_));
 sky130_fd_sc_hd__mux4_1 _2267_ (.A0(net973),
    .A1(net968),
    .A2(net987),
    .A3(net992),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1257_));
 sky130_fd_sc_hd__mux4_1 _2268_ (.A0(net978),
    .A1(net997),
    .A2(net1019),
    .A3(net1014),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1258_));
 sky130_fd_sc_hd__o21a_1 _2269_ (.A1(_0129_),
    .A2(_1258_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_1259_));
 sky130_fd_sc_hd__o21ai_1 _2270_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_1257_),
    .B1(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__nor2_1 _2271_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .B(_0302_),
    .Y(_1261_));
 sky130_fd_sc_hd__a211o_1 _2272_ (.A1(_0059_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .C1(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__mux2_1 _2273_ (.A0(net209),
    .A1(net1068),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1263_));
 sky130_fd_sc_hd__nand2_1 _2274_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .B(_1263_),
    .Y(_1264_));
 sky130_fd_sc_hd__mux4_1 _2275_ (.A0(net175),
    .A1(net1218),
    .A2(net183),
    .A3(net129),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1265_));
 sky130_fd_sc_hd__nor2_1 _2276_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .B(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__a311o_1 _2277_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_1262_),
    .A3(_1264_),
    .B1(_1266_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_1267_));
 sky130_fd_sc_hd__nand2_2 _2278_ (.A(_1260_),
    .B(_1267_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__o21ai_1 _2279_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .Y(_1268_));
 sky130_fd_sc_hd__o221a_1 _2280_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .A2(_1244_),
    .B1(_1256_),
    .B2(_1268_),
    .C1(_0128_),
    .X(_1269_));
 sky130_fd_sc_hd__o21ba_4 _2281_ (.A1(_1242_),
    .A2(_0128_),
    .B1_N(_1269_),
    .X(\Tile_X0Y1_DSP_bot.C9 ));
 sky130_fd_sc_hd__nand2b_1 _2282_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ),
    .B(net1064),
    .Y(_1270_));
 sky130_fd_sc_hd__o211a_1 _2283_ (.A1(net1063),
    .A2(\Tile_X0Y1_DSP_bot.C9 ),
    .B1(_1270_),
    .C1(net1057),
    .X(_1271_));
 sky130_fd_sc_hd__xor2_1 _2284_ (.A(_1094_),
    .B(_0994_),
    .X(_1272_));
 sky130_fd_sc_hd__nor3_2 _2285_ (.A(_1271_),
    .B(_1194_),
    .C(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__inv_2 _2286_ (.A(net616),
    .Y(_1274_));
 sky130_fd_sc_hd__o21a_1 _2287_ (.A1(_1194_),
    .A2(_1271_),
    .B1(_1272_),
    .X(_1275_));
 sky130_fd_sc_hd__nor2_2 _2288_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .B(_0529_),
    .Y(_1276_));
 sky130_fd_sc_hd__a211o_1 _2289_ (.A1(_0349_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .B1(_1276_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1277_));
 sky130_fd_sc_hd__mux2_1 _2290_ (.A0(net76),
    .A1(net1067),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1278_));
 sky130_fd_sc_hd__nand2_1 _2291_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__mux4_1 _2292_ (.A0(net176),
    .A1(net184),
    .A2(net1217),
    .A3(net130),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1280_));
 sky130_fd_sc_hd__nor2_1 _2293_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .B(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__a311o_1 _2294_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_1279_),
    .A3(_1277_),
    .B1(_1281_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_1 _2295_ (.A0(net978),
    .A1(net983),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1283_));
 sky130_fd_sc_hd__inv_1 _2296_ (.A(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__mux2_1 _2297_ (.A0(net1019),
    .A1(net1014),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1285_));
 sky130_fd_sc_hd__nand2_1 _2298_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .B(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__o211a_1 _2299_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .A2(_1284_),
    .B1(_1286_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_1287_));
 sky130_fd_sc_hd__mux4_1 _2300_ (.A0(net973),
    .A1(net969),
    .A2(net987),
    .A3(net993),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1288_));
 sky130_fd_sc_hd__o21ai_1 _2301_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_1288_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ),
    .Y(_1289_));
 sky130_fd_sc_hd__o21ai_4 _2302_ (.A1(_1287_),
    .A2(_1289_),
    .B1(_1282_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _2303_ (.A0(net973),
    .A1(net968),
    .A2(net987),
    .A3(net992),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1290_));
 sky130_fd_sc_hd__mux4_1 _2304_ (.A0(net978),
    .A1(net1019),
    .A2(net984),
    .A3(net1014),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1291_));
 sky130_fd_sc_hd__nor2_1 _2305_ (.A(_0135_),
    .B(_1291_),
    .Y(_1292_));
 sky130_fd_sc_hd__o21ai_1 _2306_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_1290_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .Y(_1293_));
 sky130_fd_sc_hd__nor2_1 _2307_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .B(_0529_),
    .Y(_1294_));
 sky130_fd_sc_hd__a211o_1 _2308_ (.A1(_0349_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .B1(_1294_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_1 _2309_ (.A0(net76),
    .A1(net1067),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1296_));
 sky130_fd_sc_hd__nand2_1 _2310_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__and3_1 _2311_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .B(_1297_),
    .C(_1295_),
    .X(_1298_));
 sky130_fd_sc_hd__mux4_1 _2312_ (.A0(net176),
    .A1(net184),
    .A2(net1217),
    .A3(net130),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1299_));
 sky130_fd_sc_hd__nor2_1 _2313_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .B(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__o32a_4 _2314_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ),
    .A2(_1300_),
    .A3(_1298_),
    .B1(_1292_),
    .B2(_1293_),
    .X(_1301_));
 sky130_fd_sc_hd__inv_4 _2315_ (.A(_1301_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__nand2_1 _2316_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .B(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__o211a_1 _2317_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .B1(_1302_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_1303_));
 sky130_fd_sc_hd__nor2_1 _2318_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .Y(_1304_));
 sky130_fd_sc_hd__a211o_1 _2319_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0557_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .C1(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__nand2_2 _2320_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .B(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__mux2_1 _2321_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_1307_));
 sky130_fd_sc_hd__mux4_1 _2322_ (.A0(net973),
    .A1(net968),
    .A2(net987),
    .A3(net992),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_1308_));
 sky130_fd_sc_hd__mux4_1 _2323_ (.A0(net978),
    .A1(net1019),
    .A2(net983),
    .A3(net1002),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_1309_));
 sky130_fd_sc_hd__o21a_1 _2324_ (.A1(_0134_),
    .A2(_1309_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .X(_1310_));
 sky130_fd_sc_hd__o21ai_1 _2325_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_1308_),
    .B1(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hd__mux2_1 _2326_ (.A0(_0349_),
    .A1(_0045_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_1312_));
 sky130_fd_sc_hd__mux2_1 _2327_ (.A0(net210),
    .A1(net1067),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_1313_));
 sky130_fd_sc_hd__nand2_1 _2328_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .B(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__o211a_1 _2329_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_1312_),
    .B1(_1314_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_1315_));
 sky130_fd_sc_hd__mux4_1 _2330_ (.A0(net176),
    .A1(net184),
    .A2(net1217),
    .A3(net130),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_1316_));
 sky130_fd_sc_hd__nor2_1 _2331_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__o31ai_4 _2332_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_1315_),
    .A3(_1317_),
    .B1(_1311_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(_1307_),
    .A1(_1318_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_1319_));
 sky130_fd_sc_hd__o22a_4 _2335_ (.A1(_1306_),
    .A2(_1303_),
    .B1(_1319_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .X(\Tile_X0Y1_DSP_bot.C8 ));
 sky130_fd_sc_hd__mux2_2 _2336_ (.A0(\Tile_X0Y1_DSP_bot.C8 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ),
    .S(net1063),
    .X(_1320_));
 sky130_fd_sc_hd__mux2_4 _2337_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ),
    .A1(_1320_),
    .S(net1057),
    .X(_1321_));
 sky130_fd_sc_hd__a21oi_1 _2338_ (.A1(_1039_),
    .A2(_1091_),
    .B1(_1020_),
    .Y(_1322_));
 sky130_fd_sc_hd__nor2_4 _2339_ (.A(_1093_),
    .B(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__and2_1 _2340_ (.A(_1321_),
    .B(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__nand2_1 _2341_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ),
    .Y(_1325_));
 sky130_fd_sc_hd__mux4_2 _2342_ (.A0(_0112_),
    .A1(_0111_),
    .A2(_0021_),
    .A3(_0557_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_1326_));
 sky130_fd_sc_hd__inv_2 _2343_ (.A(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__nand2_1 _2344_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .B(_1326_),
    .Y(_1328_));
 sky130_fd_sc_hd__mux4_2 _2345_ (.A0(net178),
    .A1(net144),
    .A2(net70),
    .A3(net214),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .X(_1329_));
 sky130_fd_sc_hd__o211a_1 _2346_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_1329_),
    .B1(_1328_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_1330_));
 sky130_fd_sc_hd__nand2_2 _2347_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .B(_1301_),
    .Y(_1331_));
 sky130_fd_sc_hd__o21a_1 _2348_ (.A1(net221),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_1332_));
 sky130_fd_sc_hd__mux2_1 _2349_ (.A0(net185),
    .A1(net131),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .X(_1333_));
 sky130_fd_sc_hd__a221o_1 _2350_ (.A1(_1332_),
    .A2(_1331_),
    .B1(_1333_),
    .B2(_0136_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_1334_));
 sky130_fd_sc_hd__mux2_4 _2351_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A1(net222),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1335_));
 sky130_fd_sc_hd__mux2_1 _2352_ (.A0(net186),
    .A1(net132),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1336_));
 sky130_fd_sc_hd__inv_1 _2353_ (.A(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__o21ai_1 _2354_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .A2(_1337_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .Y(_1338_));
 sky130_fd_sc_hd__a21o_1 _2355_ (.A1(_1335_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ),
    .B1(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__a31o_4 _2356_ (.A1(_0137_),
    .A2(_1334_),
    .A3(_1339_),
    .B1(_1330_),
    .X(\Tile_X0Y1_DSP_bot.C7 ));
 sky130_fd_sc_hd__mux2_4 _2357_ (.A0(\Tile_X0Y1_DSP_bot.C7 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ),
    .S(net1063),
    .X(_1340_));
 sky130_fd_sc_hd__nand2_4 _2358_ (.A(net1057),
    .B(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__xnor2_2 _2359_ (.A(_1090_),
    .B(_1092_),
    .Y(_1342_));
 sky130_fd_sc_hd__a21oi_2 _2360_ (.A1(_1325_),
    .A2(_1341_),
    .B1(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__nand3_4 _2361_ (.A(_1325_),
    .B(_1341_),
    .C(_1342_),
    .Y(_1344_));
 sky130_fd_sc_hd__nand2b_4 _2362_ (.A_N(_1343_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__mux4_2 _2363_ (.A0(net140),
    .A1(net82),
    .A2(net234),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_1346_));
 sky130_fd_sc_hd__mux4_2 _2364_ (.A0(net202),
    .A1(net128),
    .A2(net74),
    .A3(net218),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .X(_1347_));
 sky130_fd_sc_hd__mux2_4 _2365_ (.A0(_1347_),
    .A1(_1346_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_1348_));
 sky130_fd_sc_hd__mux4_2 _2366_ (.A0(net135),
    .A1(net225),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .X(_1349_));
 sky130_fd_sc_hd__mux2_1 _2367_ (.A0(net190),
    .A1(net136),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_1350_));
 sky130_fd_sc_hd__and2b_1 _2368_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .B(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__mux2_4 _2369_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A1(net226),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_1352_));
 sky130_fd_sc_hd__a21bo_1 _2370_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ),
    .A2(_1352_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_1353_));
 sky130_fd_sc_hd__o22a_1 _2371_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1349_),
    .B1(_1351_),
    .B2(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__mux2_4 _2372_ (.A0(_1354_),
    .A1(_1348_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ),
    .X(\Tile_X0Y1_DSP_bot.C6 ));
 sky130_fd_sc_hd__mux2_1 _2373_ (.A0(\Tile_X0Y1_DSP_bot.C6 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ),
    .S(net1063),
    .X(_1355_));
 sky130_fd_sc_hd__mux2_4 _2374_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ),
    .A1(_1355_),
    .S(net1057),
    .X(_1356_));
 sky130_fd_sc_hd__xnor2_2 _2375_ (.A(_1089_),
    .B(_1055_),
    .Y(_1357_));
 sky130_fd_sc_hd__and2b_1 _2376_ (.A_N(_1357_),
    .B(_1356_),
    .X(_1358_));
 sky130_fd_sc_hd__xnor2_2 _2377_ (.A(_1357_),
    .B(_1356_),
    .Y(_1359_));
 sky130_fd_sc_hd__mux4_2 _2378_ (.A0(net187),
    .A1(net223),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_1360_));
 sky130_fd_sc_hd__mux4_2 _2379_ (.A0(net188),
    .A1(net134),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(net224),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .X(_1361_));
 sky130_fd_sc_hd__mux2_2 _2380_ (.A0(_1360_),
    .A1(net1003),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_1362_));
 sky130_fd_sc_hd__mux4_2 _2381_ (.A0(net195),
    .A1(net215),
    .A2(net91),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_1363_));
 sky130_fd_sc_hd__mux4_1 _2382_ (.A0(net180),
    .A1(net126),
    .A2(net89),
    .A3(net216),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_1364_));
 sky130_fd_sc_hd__mux2_4 _2383_ (.A0(_1364_),
    .A1(_1363_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_4 _2384_ (.A0(_1362_),
    .A1(_1365_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .X(\Tile_X0Y1_DSP_bot.C5 ));
 sky130_fd_sc_hd__mux2_2 _2385_ (.A0(\Tile_X0Y1_DSP_bot.C5 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ),
    .S(net1063),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_4 _2386_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ),
    .A1(_1366_),
    .S(net1057),
    .X(_1367_));
 sky130_fd_sc_hd__xnor2_4 _2387_ (.A(_1088_),
    .B(_1070_),
    .Y(_1368_));
 sky130_fd_sc_hd__and2b_1 _2388_ (.A_N(_1368_),
    .B(_1367_),
    .X(_1369_));
 sky130_fd_sc_hd__xnor2_4 _2389_ (.A(_1368_),
    .B(_1367_),
    .Y(_1370_));
 sky130_fd_sc_hd__mux2_1 _2390_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_1371_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(net191),
    .A1(net137),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_1372_));
 sky130_fd_sc_hd__and2b_1 _2392_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .B(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__a211o_1 _2393_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .A2(_1371_),
    .B1(_1373_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_1374_));
 sky130_fd_sc_hd__mux2_1 _2394_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .A1(net228),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_1375_));
 sky130_fd_sc_hd__nand2_1 _2395_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .B(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__mux2_1 _2396_ (.A0(net192),
    .A1(net138),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_1377_));
 sky130_fd_sc_hd__inv_1 _2397_ (.A(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__o211a_1 _2398_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .A2(_1378_),
    .B1(_1376_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_1379_));
 sky130_fd_sc_hd__nor2_1 _2399_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__mux4_1 _2400_ (.A0(net196),
    .A1(net84),
    .A2(net141),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_1381_));
 sky130_fd_sc_hd__mux4_1 _2401_ (.A0(net184),
    .A1(net130),
    .A2(net76),
    .A3(net231),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .X(_1382_));
 sky130_fd_sc_hd__mux2_1 _2402_ (.A0(_1382_),
    .A1(_1381_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_1383_));
 sky130_fd_sc_hd__a22o_1 _2403_ (.A1(_1374_),
    .A2(_1380_),
    .B1(_1383_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .X(\Tile_X0Y1_DSP_bot.C4 ));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(\Tile_X0Y1_DSP_bot.C4 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ),
    .S(net1063),
    .X(_1384_));
 sky130_fd_sc_hd__mux2_1 _2405_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ),
    .A1(_1384_),
    .S(net1057),
    .X(_1385_));
 sky130_fd_sc_hd__a21o_1 _2406_ (.A1(_1079_),
    .A2(_1086_),
    .B1(_1085_),
    .X(_1386_));
 sky130_fd_sc_hd__and3_1 _2407_ (.A(_1087_),
    .B(_1385_),
    .C(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__a21oi_1 _2408_ (.A1(_1087_),
    .A2(_1386_),
    .B1(_1385_),
    .Y(_1388_));
 sky130_fd_sc_hd__nor2_4 _2409_ (.A(_1388_),
    .B(_1387_),
    .Y(_1389_));
 sky130_fd_sc_hd__mux4_1 _2410_ (.A0(net144),
    .A1(net232),
    .A2(net81),
    .A3(_0184_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_1390_));
 sky130_fd_sc_hd__mux4_2 _2411_ (.A0(net203),
    .A1(net124),
    .A2(net70),
    .A3(net214),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .X(_1391_));
 sky130_fd_sc_hd__mux2_1 _2412_ (.A0(_1391_),
    .A1(_1390_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_1392_));
 sky130_fd_sc_hd__mux2_1 _2413_ (.A0(net221),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_1393_));
 sky130_fd_sc_hd__mux2_4 _2414_ (.A0(net131),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_1394_));
 sky130_fd_sc_hd__and2b_1 _2415_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .B(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__a211o_1 _2416_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .A2(_1393_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .C1(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__mux2_1 _2417_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A1(net222),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_1397_));
 sky130_fd_sc_hd__nand2_1 _2418_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .B(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(net186),
    .A1(net132),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_1399_));
 sky130_fd_sc_hd__inv_1 _2420_ (.A(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__o211a_1 _2421_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .A2(_1400_),
    .B1(_1398_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_1401_));
 sky130_fd_sc_hd__nor2_1 _2422_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .B(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__a22o_4 _2423_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .A2(_1392_),
    .B1(_1402_),
    .B2(_1396_),
    .X(\Tile_X0Y1_DSP_bot.C3 ));
 sky130_fd_sc_hd__mux2_4 _2424_ (.A0(\Tile_X0Y1_DSP_bot.C3 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ),
    .S(net1063),
    .X(_1403_));
 sky130_fd_sc_hd__mux2_4 _2425_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ),
    .A1(_1403_),
    .S(net1057),
    .X(_1404_));
 sky130_fd_sc_hd__xnor2_1 _2426_ (.A(_1080_),
    .B(_1084_),
    .Y(_1405_));
 sky130_fd_sc_hd__nand2b_4 _2427_ (.A_N(_1405_),
    .B(_1404_),
    .Y(_1406_));
 sky130_fd_sc_hd__xor2_1 _2428_ (.A(_1404_),
    .B(_1405_),
    .X(_1407_));
 sky130_fd_sc_hd__mux4_1 _2429_ (.A0(net182),
    .A1(net128),
    .A2(net90),
    .A3(net218),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .X(_1408_));
 sky130_fd_sc_hd__mux2_4 _2430_ (.A0(_1408_),
    .A1(_0230_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_1409_));
 sky130_fd_sc_hd__mux4_2 _2431_ (.A0(net189),
    .A1(net225),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1410_));
 sky130_fd_sc_hd__mux4_2 _2432_ (.A0(net190),
    .A1(net136),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A3(net226),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_1 _2433_ (.A0(_1410_),
    .A1(_1411_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_1412_));
 sky130_fd_sc_hd__mux2_4 _2434_ (.A0(_1412_),
    .A1(_1409_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .X(\Tile_X0Y1_DSP_bot.C2 ));
 sky130_fd_sc_hd__mux2_4 _2435_ (.A0(\Tile_X0Y1_DSP_bot.C2 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ),
    .S(net1063),
    .X(_1413_));
 sky130_fd_sc_hd__mux2_4 _2436_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ),
    .A1(_1413_),
    .S(net1057),
    .X(_1414_));
 sky130_fd_sc_hd__xor2_4 _2437_ (.A(_1083_),
    .B(_1082_),
    .X(_1415_));
 sky130_fd_sc_hd__xnor2_2 _2438_ (.A(_1415_),
    .B(_1414_),
    .Y(_1416_));
 sky130_fd_sc_hd__mux2_1 _2439_ (.A0(net83),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1417_));
 sky130_fd_sc_hd__mux2_1 _2440_ (.A0(net203),
    .A1(net125),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1418_));
 sky130_fd_sc_hd__o21a_1 _2441_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_1418_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_1419_));
 sky130_fd_sc_hd__o21ai_1 _2442_ (.A1(_0138_),
    .A2(_1417_),
    .B1(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__mux4_1 _2443_ (.A0(net180),
    .A1(net126),
    .A2(net72),
    .A3(net232),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_1421_));
 sky130_fd_sc_hd__inv_2 _2444_ (.A(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__o211a_1 _2445_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_1422_),
    .B1(_1420_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .X(_1423_));
 sky130_fd_sc_hd__nand2_1 _2446_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .Y(_1424_));
 sky130_fd_sc_hd__or2_4 _2447_ (.A(_0632_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_1425_));
 sky130_fd_sc_hd__mux2_1 _2448_ (.A0(net187),
    .A1(net133),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_1426_));
 sky130_fd_sc_hd__nor2_1 _2449_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .B(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__a311o_1 _2450_ (.A1(_1425_),
    .A2(_1424_),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .B1(_1427_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_1428_));
 sky130_fd_sc_hd__mux4_2 _2451_ (.A0(net188),
    .A1(net134),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(net224),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_1429_));
 sky130_fd_sc_hd__a21oi_1 _2452_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_1429_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_1430_));
 sky130_fd_sc_hd__a21oi_2 _2453_ (.A1(_1430_),
    .A2(_1428_),
    .B1(_1423_),
    .Y(\Tile_X0Y1_DSP_bot.C1 ));
 sky130_fd_sc_hd__mux2_2 _2454_ (.A0(\Tile_X0Y1_DSP_bot.C1 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ),
    .S(net1063),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_4 _2455_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ),
    .A1(_1431_),
    .S(net1057),
    .X(_1432_));
 sky130_fd_sc_hd__o22a_1 _2456_ (.A1(net624),
    .A2(_0944_),
    .B1(_0981_),
    .B2(_0785_),
    .X(_1433_));
 sky130_fd_sc_hd__a21o_1 _2457_ (.A1(_1073_),
    .A2(_1081_),
    .B1(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__inv_1 _2458_ (.A(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__mux4_1 _2459_ (.A0(net196),
    .A1(net126),
    .A2(net216),
    .A3(net658),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_1436_));
 sky130_fd_sc_hd__mux4_1 _2460_ (.A0(net184),
    .A1(net143),
    .A2(net76),
    .A3(net220),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_1437_));
 sky130_fd_sc_hd__mux2_1 _2461_ (.A0(_1437_),
    .A1(_1436_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_1438_));
 sky130_fd_sc_hd__mux4_2 _2462_ (.A0(net191),
    .A1(net227),
    .A2(net137),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .X(_1439_));
 sky130_fd_sc_hd__mux2_4 _2463_ (.A0(_1439_),
    .A1(_0216_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_1440_));
 sky130_fd_sc_hd__mux2_4 _2464_ (.A0(_1440_),
    .A1(_1438_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .X(\Tile_X0Y1_DSP_bot.C0 ));
 sky130_fd_sc_hd__mux2_2 _2465_ (.A0(\Tile_X0Y1_DSP_bot.C0 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ),
    .S(net1063),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_4 _2466_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ),
    .A1(_1441_),
    .S(net1057),
    .X(_1442_));
 sky130_fd_sc_hd__and2_4 _2467_ (.A(_1081_),
    .B(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__xor2_4 _2468_ (.A(_1434_),
    .B(_1432_),
    .X(_1444_));
 sky130_fd_sc_hd__nor4b_4 _2469_ (.A(_1444_),
    .B(_0981_),
    .C(_0878_),
    .D_N(_1442_),
    .Y(_1445_));
 sky130_fd_sc_hd__a21oi_2 _2470_ (.A1(_1432_),
    .A2(_1435_),
    .B1(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__or2_4 _2471_ (.A(_1416_),
    .B(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__a21boi_4 _2472_ (.A1(_1414_),
    .A2(_1415_),
    .B1_N(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__o21a_4 _2473_ (.A1(_1407_),
    .A2(_1448_),
    .B1(_1406_),
    .X(_1449_));
 sky130_fd_sc_hd__o21bai_4 _2474_ (.A1(_1388_),
    .A2(_1449_),
    .B1_N(_1387_),
    .Y(_1450_));
 sky130_fd_sc_hd__a21o_1 _2475_ (.A1(_1370_),
    .A2(_1450_),
    .B1(_1369_),
    .X(_1451_));
 sky130_fd_sc_hd__a21o_1 _2476_ (.A1(_1451_),
    .A2(_1359_),
    .B1(_1358_),
    .X(_1452_));
 sky130_fd_sc_hd__a21o_1 _2477_ (.A1(_1452_),
    .A2(_1344_),
    .B1(_1343_),
    .X(_1453_));
 sky130_fd_sc_hd__xor2_2 _2478_ (.A(_1323_),
    .B(_1321_),
    .X(_1454_));
 sky130_fd_sc_hd__a21o_1 _2479_ (.A1(_1454_),
    .A2(_1453_),
    .B1(_1324_),
    .X(_1455_));
 sky130_fd_sc_hd__a211o_4 _2480_ (.A1(_1453_),
    .A2(_1454_),
    .B1(_1324_),
    .C1(_1275_),
    .X(_1456_));
 sky130_fd_sc_hd__and3_1 _2481_ (.A(_1193_),
    .B(_1456_),
    .C(_1274_),
    .X(_1457_));
 sky130_fd_sc_hd__a31o_4 _2482_ (.A1(_1193_),
    .A2(_1456_),
    .A3(_1274_),
    .B1(_1192_),
    .X(_1458_));
 sky130_fd_sc_hd__a21o_1 _2483_ (.A1(_1458_),
    .A2(_1173_),
    .B1(_1172_),
    .X(_1459_));
 sky130_fd_sc_hd__a21o_1 _2484_ (.A1(_1459_),
    .A2(_1157_),
    .B1(_1156_),
    .X(_1460_));
 sky130_fd_sc_hd__a21oi_4 _2485_ (.A1(_1460_),
    .A2(_1144_),
    .B1(_1146_),
    .Y(_1461_));
 sky130_fd_sc_hd__xor2_1 _2486_ (.A(_1118_),
    .B(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_4 _2487_ (.A0(_1462_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ));
 sky130_fd_sc_hd__nand2_1 _2488_ (.A(_1416_),
    .B(_1446_),
    .Y(_1463_));
 sky130_fd_sc_hd__and2_4 _2489_ (.A(_1447_),
    .B(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__mux2_4 _2490_ (.A0(_1464_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ));
 sky130_fd_sc_hd__nor2_1 _2491_ (.A(_1081_),
    .B(_1442_),
    .Y(_1465_));
 sky130_fd_sc_hd__nor2_1 _2492_ (.A(_1443_),
    .B(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__mux2_2 _2493_ (.A0(_1466_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ));
 sky130_fd_sc_hd__xnor2_2 _2494_ (.A(_1389_),
    .B(_1449_),
    .Y(_1467_));
 sky130_fd_sc_hd__mux2_4 _2495_ (.A0(_1467_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ));
 sky130_fd_sc_hd__xor2_1 _2496_ (.A(_1407_),
    .B(_1448_),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_4 _2497_ (.A0(_1468_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ));
 sky130_fd_sc_hd__xor2_1 _2498_ (.A(_1450_),
    .B(_1370_),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_4 _2499_ (.A0(_1469_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ));
 sky130_fd_sc_hd__xor2_1 _2500_ (.A(_1451_),
    .B(_1359_),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_4 _2501_ (.A0(_1470_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ));
 sky130_fd_sc_hd__xnor2_2 _2502_ (.A(_1345_),
    .B(_1452_),
    .Y(_1471_));
 sky130_fd_sc_hd__mux2_4 _2503_ (.A0(_1471_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ));
 sky130_fd_sc_hd__nor2_2 _2504_ (.A(_1273_),
    .B(_1275_),
    .Y(_1472_));
 sky130_fd_sc_hd__xor2_1 _2505_ (.A(_1455_),
    .B(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_4 _2506_ (.A0(_1473_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ));
 sky130_fd_sc_hd__mux4_2 _2507_ (.A0(net977),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .A2(net1003),
    .A3(_1327_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ));
 sky130_fd_sc_hd__a21oi_1 _2508_ (.A1(_1274_),
    .A2(_1456_),
    .B1(_1193_),
    .Y(_1474_));
 sky130_fd_sc_hd__nor2_2 _2509_ (.A(_1474_),
    .B(_1457_),
    .Y(_1475_));
 sky130_fd_sc_hd__mux2_4 _2510_ (.A0(_1475_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ));
 sky130_fd_sc_hd__xor2_2 _2511_ (.A(_1174_),
    .B(_1458_),
    .X(_1476_));
 sky130_fd_sc_hd__inv_2 _2512_ (.A(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__mux2_4 _2513_ (.A0(_1477_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ));
 sky130_fd_sc_hd__xor2_1 _2514_ (.A(_1459_),
    .B(_1157_),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_4 _2515_ (.A0(_1478_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ));
 sky130_fd_sc_hd__o21a_1 _2516_ (.A1(_1118_),
    .A2(_1461_),
    .B1(_1117_),
    .X(_1479_));
 sky130_fd_sc_hd__o21bai_2 _2517_ (.A1(_0843_),
    .A2(_1113_),
    .B1_N(_1103_),
    .Y(_1480_));
 sky130_fd_sc_hd__nand2_1 _2518_ (.A(_1115_),
    .B(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__and2_1 _2519_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ),
    .X(_1482_));
 sky130_fd_sc_hd__mux4_1 _2520_ (.A0(net1012),
    .A1(net1047),
    .A2(net1027),
    .A3(net1051),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1483_));
 sky130_fd_sc_hd__and2_1 _2521_ (.A(_0094_),
    .B(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__mux4_2 _2522_ (.A0(net1043),
    .A1(net1032),
    .A2(net1038),
    .A3(net1022),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1485_));
 sky130_fd_sc_hd__a21bo_1 _2523_ (.A1(_1485_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(net675),
    .A1(net192),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1487_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(net1257),
    .A1(net12),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1488_));
 sky130_fd_sc_hd__or2_1 _2526_ (.A(_0093_),
    .B(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__o211a_1 _2527_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .A2(_1487_),
    .B1(_1489_),
    .C1(_0094_),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(net58),
    .A1(net60),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1491_));
 sky130_fd_sc_hd__or2_1 _2529_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .B(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(net68),
    .A1(net1219),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_1493_));
 sky130_fd_sc_hd__o211a_1 _2531_ (.A1(_0093_),
    .A2(_1493_),
    .B1(_1492_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_1494_));
 sky130_fd_sc_hd__o32a_4 _2532_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_1490_),
    .A3(_1494_),
    .B1(_1486_),
    .B2(_1484_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _2533_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A1(net107),
    .A2(net71),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_4 _2534_ (.A0(_1495_),
    .A1(_0299_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_1496_));
 sky130_fd_sc_hd__mux4_1 _2535_ (.A0(net199),
    .A1(net87),
    .A2(net99),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_1497_));
 sky130_fd_sc_hd__mux4_2 _2536_ (.A0(net188),
    .A1(net8),
    .A2(net85),
    .A3(net100),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(_1498_),
    .A1(_1497_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_4 _2538_ (.A0(_1496_),
    .A1(_1499_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ));
 sky130_fd_sc_hd__mux2_4 _2539_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ),
    .S(net1064),
    .X(_1500_));
 sky130_fd_sc_hd__a21oi_2 _2540_ (.A1(_1500_),
    .A2(net1058),
    .B1(_1482_),
    .Y(_1501_));
 sky130_fd_sc_hd__and3_4 _2541_ (.A(_1115_),
    .B(_1480_),
    .C(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__a21o_1 _2542_ (.A1(_1115_),
    .A2(_1480_),
    .B1(_1501_),
    .X(_1503_));
 sky130_fd_sc_hd__and2b_1 _2543_ (.A_N(_1502_),
    .B(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__xnor2_2 _2544_ (.A(_1504_),
    .B(_1479_),
    .Y(_1505_));
 sky130_fd_sc_hd__mux2_4 _2545_ (.A0(_1505_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ));
 sky130_fd_sc_hd__a21bo_2 _2546_ (.A1(_1115_),
    .A2(_1480_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ),
    .X(_1506_));
 sky130_fd_sc_hd__and2_1 _2547_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ),
    .X(_1507_));
 sky130_fd_sc_hd__mux4_1 _2548_ (.A0(net22),
    .A1(net78),
    .A2(net118),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_1508_));
 sky130_fd_sc_hd__mux4_1 _2549_ (.A0(net206),
    .A1(net66),
    .A2(net10),
    .A3(net102),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(_1509_),
    .A1(_1508_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_1510_));
 sky130_fd_sc_hd__mux4_2 _2551_ (.A0(net710),
    .A1(net74),
    .A2(net18),
    .A3(net110),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_1511_));
 sky130_fd_sc_hd__mux4_2 _2552_ (.A0(net17),
    .A1(net109),
    .A2(net73),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_4 _2553_ (.A0(_1512_),
    .A1(_1511_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_4 _2554_ (.A0(_1513_),
    .A1(_1510_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ));
 sky130_fd_sc_hd__mux2_4 _2555_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ),
    .S(net1064),
    .X(_1514_));
 sky130_fd_sc_hd__a21oi_4 _2556_ (.A1(net1058),
    .A2(_1514_),
    .B1(_1507_),
    .Y(_1515_));
 sky130_fd_sc_hd__or2_1 _2557_ (.A(_1506_),
    .B(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__xnor2_2 _2558_ (.A(_1506_),
    .B(_1515_),
    .Y(_1517_));
 sky130_fd_sc_hd__o211a_4 _2559_ (.A1(_1118_),
    .A2(_1461_),
    .B1(_1117_),
    .C1(_1503_),
    .X(_1518_));
 sky130_fd_sc_hd__nor2_2 _2560_ (.A(_1502_),
    .B(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__xnor2_1 _2561_ (.A(_1517_),
    .B(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__mux2_4 _2562_ (.A0(_1520_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ));
 sky130_fd_sc_hd__o31a_1 _2563_ (.A1(_1502_),
    .A2(_1517_),
    .A3(_1518_),
    .B1(_1516_),
    .X(_1521_));
 sky130_fd_sc_hd__mux4_2 _2564_ (.A0(net186),
    .A1(net62),
    .A2(net26),
    .A3(net98),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_1522_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(_1522_),
    .A1(_0278_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_1523_));
 sky130_fd_sc_hd__mux4_1 _2566_ (.A0(net1011),
    .A1(net1047),
    .A2(net1026),
    .A3(net1052),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1524_));
 sky130_fd_sc_hd__and2_1 _2567_ (.A(_0098_),
    .B(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__mux4_1 _2568_ (.A0(net1042),
    .A1(net1033),
    .A2(net1037),
    .A3(net1021),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1526_));
 sky130_fd_sc_hd__a21bo_1 _2569_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_1526_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ),
    .X(_1527_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(net674),
    .A1(net192),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(net1257),
    .A1(net12),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1529_));
 sky130_fd_sc_hd__or2_1 _2572_ (.A(_0097_),
    .B(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__o211a_1 _2573_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .A2(_1528_),
    .B1(_1530_),
    .C1(_0098_),
    .X(_1531_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(net58),
    .A1(net60),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1532_));
 sky130_fd_sc_hd__or2_1 _2575_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .B(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(net68),
    .A1(net1219),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_1534_));
 sky130_fd_sc_hd__o211a_1 _2577_ (.A1(_0097_),
    .A2(_1534_),
    .B1(_1533_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ),
    .X(_1535_));
 sky130_fd_sc_hd__o32a_2 _2578_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ),
    .A2(_1531_),
    .A3(_1535_),
    .B1(_1525_),
    .B2(_1527_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _2579_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .A1(net105),
    .A2(net13),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(net690),
    .A1(net14),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1537_));
 sky130_fd_sc_hd__and2b_1 _2581_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ),
    .B(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(net70),
    .A1(net106),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1539_));
 sky130_fd_sc_hd__a21bo_1 _2583_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ),
    .A2(_1539_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_1540_));
 sky130_fd_sc_hd__o22a_1 _2584_ (.A1(_1536_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .B1(_1538_),
    .B2(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__mux2_4 _2585_ (.A0(_1541_),
    .A1(_1523_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ));
 sky130_fd_sc_hd__mux2_4 _2586_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ),
    .S(net1064),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_4 _2587_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ),
    .A1(_1542_),
    .S(net1058),
    .X(_1543_));
 sky130_fd_sc_hd__and3_1 _2588_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ),
    .B(_1543_),
    .C(_1481_),
    .X(_1544_));
 sky130_fd_sc_hd__nand2b_1 _2589_ (.A_N(_1506_),
    .B(_1543_),
    .Y(_1545_));
 sky130_fd_sc_hd__a21oi_1 _2590_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ),
    .A2(_1481_),
    .B1(_1543_),
    .Y(_1546_));
 sky130_fd_sc_hd__nor2_4 _2591_ (.A(_1546_),
    .B(_1544_),
    .Y(_1547_));
 sky130_fd_sc_hd__xnor2_2 _2592_ (.A(_1547_),
    .B(_1521_),
    .Y(_1548_));
 sky130_fd_sc_hd__mux2_4 _2593_ (.A0(_1548_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ));
 sky130_fd_sc_hd__a21bo_1 _2594_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1549_));
 sky130_fd_sc_hd__a21o_1 _2595_ (.A1(_0139_),
    .A2(_0274_),
    .B1(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__mux2_1 _2596_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_1551_));
 sky130_fd_sc_hd__o21a_1 _2597_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .A2(_1551_),
    .B1(_1550_),
    .X(_1552_));
 sky130_fd_sc_hd__mux2_4 _2598_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_1553_));
 sky130_fd_sc_hd__nand2_1 _2599_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .Y(_1554_));
 sky130_fd_sc_hd__o211a_1 _2600_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(_0696_),
    .B1(_1554_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1555_));
 sky130_fd_sc_hd__o21ba_1 _2601_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .A2(_1553_),
    .B1_N(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_4 _2602_ (.A0(_1556_),
    .A1(_1552_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ));
 sky130_fd_sc_hd__mux2_2 _2603_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ),
    .S(net1064),
    .X(_1557_));
 sky130_fd_sc_hd__mux2_4 _2604_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ),
    .A1(_1557_),
    .S(net1058),
    .X(_1558_));
 sky130_fd_sc_hd__nand2b_1 _2605_ (.A_N(_1506_),
    .B(_1558_),
    .Y(_1559_));
 sky130_fd_sc_hd__xor2_2 _2606_ (.A(_1506_),
    .B(_1558_),
    .X(_1560_));
 sky130_fd_sc_hd__o311a_1 _2607_ (.A1(_1502_),
    .A2(_1517_),
    .A3(_1518_),
    .B1(_1545_),
    .C1(_1516_),
    .X(_1561_));
 sky130_fd_sc_hd__nor2_1 _2608_ (.A(_1546_),
    .B(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__o31a_1 _2609_ (.A1(_1546_),
    .A2(_1560_),
    .A3(_1561_),
    .B1(_1559_),
    .X(_1563_));
 sky130_fd_sc_hd__mux2_1 _2610_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_1564_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(net744),
    .A1(net185),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_2 _2612_ (.A0(net1),
    .A1(net5),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1566_));
 sky130_fd_sc_hd__or2_4 _2613_ (.A(_0145_),
    .B(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__o211a_1 _2614_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .A2(_1565_),
    .B1(_1567_),
    .C1(_0146_),
    .X(_1568_));
 sky130_fd_sc_hd__mux2_2 _2615_ (.A0(net57),
    .A1(net59),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1569_));
 sky130_fd_sc_hd__or2_4 _2616_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .B(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(net61),
    .A1(net93),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1571_));
 sky130_fd_sc_hd__o211a_1 _2618_ (.A1(_0145_),
    .A2(_1571_),
    .B1(_1570_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .X(_1572_));
 sky130_fd_sc_hd__mux4_1 _2619_ (.A0(net1012),
    .A1(net1048),
    .A2(net1027),
    .A3(net1051),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1573_));
 sky130_fd_sc_hd__mux4_1 _2620_ (.A0(net1044),
    .A1(net1008),
    .A2(net1038),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_1574_));
 sky130_fd_sc_hd__a21bo_1 _2621_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(_1574_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_1575_));
 sky130_fd_sc_hd__a21o_1 _2622_ (.A1(_0146_),
    .A2(_1573_),
    .B1(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__o311a_1 _2623_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ),
    .A2(_1572_),
    .A3(_1568_),
    .B1(_1576_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_1577_));
 sky130_fd_sc_hd__o21ai_1 _2624_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_1127_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .Y(_1578_));
 sky130_fd_sc_hd__o221a_1 _2625_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(_1564_),
    .B1(_1578_),
    .B2(_1577_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_1579_));
 sky130_fd_sc_hd__mux4_1 _2626_ (.A0(net1012),
    .A1(net1047),
    .A2(net1027),
    .A3(net1051),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1580_));
 sky130_fd_sc_hd__and2_1 _2627_ (.A(_0143_),
    .B(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__mux4_1 _2628_ (.A0(net1043),
    .A1(net740),
    .A2(net1038),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1582_));
 sky130_fd_sc_hd__a21bo_1 _2629_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_1582_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_1583_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(_0199_),
    .A1(net185),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1584_));
 sky130_fd_sc_hd__mux2_1 _2631_ (.A0(net1),
    .A1(net5),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1585_));
 sky130_fd_sc_hd__or2_1 _2632_ (.A(_0142_),
    .B(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__o211a_1 _2633_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .A2(_1584_),
    .B1(_1586_),
    .C1(_0143_),
    .X(_1587_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(net57),
    .A1(net59),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1588_));
 sky130_fd_sc_hd__or2_1 _2635_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .B(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(net85),
    .A1(net115),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1590_));
 sky130_fd_sc_hd__o211a_1 _2637_ (.A1(_0142_),
    .A2(_1590_),
    .B1(_1589_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_1591_));
 sky130_fd_sc_hd__o32a_1 _2638_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_1587_),
    .A3(_1591_),
    .B1(_1581_),
    .B2(_1583_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__mux2_1 _2639_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_1592_));
 sky130_fd_sc_hd__or2_1 _2640_ (.A(_0144_),
    .B(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__mux4_1 _2641_ (.A0(net1011),
    .A1(net1047),
    .A2(net1026),
    .A3(net1052),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_1594_));
 sky130_fd_sc_hd__and2_1 _2642_ (.A(_0141_),
    .B(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__mux4_1 _2643_ (.A0(net1042),
    .A1(net1007),
    .A2(net1037),
    .A3(net1021),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1596_));
 sky130_fd_sc_hd__a21bo_1 _2644_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_1596_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_1597_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(_0199_),
    .A1(net185),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1598_));
 sky130_fd_sc_hd__mux2_1 _2646_ (.A0(net1),
    .A1(net23),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1599_));
 sky130_fd_sc_hd__or2_1 _2647_ (.A(_0140_),
    .B(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__o211a_1 _2648_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_1598_),
    .B1(_1600_),
    .C1(_0141_),
    .X(_1601_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(net57),
    .A1(net61),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1602_));
 sky130_fd_sc_hd__or2_1 _2650_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .B(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _2651_ (.A0(net93),
    .A1(net1220),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_1604_));
 sky130_fd_sc_hd__o211a_1 _2652_ (.A1(_0140_),
    .A2(_1604_),
    .B1(_1603_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_1605_));
 sky130_fd_sc_hd__o32a_1 _2653_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ),
    .A2(_1601_),
    .A3(_1605_),
    .B1(_1595_),
    .B2(_1597_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ));
 sky130_fd_sc_hd__nor2_1 _2654_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .B(_1186_),
    .Y(_1606_));
 sky130_fd_sc_hd__a211o_1 _2655_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ),
    .B1(_1606_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_1607_));
 sky130_fd_sc_hd__a31o_1 _2656_ (.A1(_0147_),
    .A2(_1593_),
    .A3(_1607_),
    .B1(_1579_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ));
 sky130_fd_sc_hd__mux2_4 _2657_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ),
    .S(net1064),
    .X(_1608_));
 sky130_fd_sc_hd__mux2_4 _2658_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ),
    .A1(_1608_),
    .S(net1058),
    .X(_1609_));
 sky130_fd_sc_hd__xnor2_2 _2659_ (.A(_1609_),
    .B(_1506_),
    .Y(_1610_));
 sky130_fd_sc_hd__xnor2_1 _2660_ (.A(_1563_),
    .B(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__mux2_4 _2661_ (.A0(_1611_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ));
 sky130_fd_sc_hd__nor2_2 _2662_ (.A(_1146_),
    .B(_1145_),
    .Y(_1612_));
 sky130_fd_sc_hd__xor2_1 _2663_ (.A(_1460_),
    .B(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_4 _2664_ (.A0(_1613_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ));
 sky130_fd_sc_hd__xnor2_1 _2665_ (.A(_1562_),
    .B(_1560_),
    .Y(_1614_));
 sky130_fd_sc_hd__mux2_4 _2666_ (.A0(_1614_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ),
    .S(net1066),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ));
 sky130_fd_sc_hd__xnor2_2 _2667_ (.A(_1443_),
    .B(_1444_),
    .Y(_1615_));
 sky130_fd_sc_hd__mux2_4 _2668_ (.A0(_1615_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ));
 sky130_fd_sc_hd__xor2_1 _2669_ (.A(_1453_),
    .B(_1454_),
    .X(_1616_));
 sky130_fd_sc_hd__mux2_4 _2670_ (.A0(_1616_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ),
    .S(net1065),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ));
 sky130_fd_sc_hd__mux4_1 _2671_ (.A0(net1012),
    .A1(net1048),
    .A2(net1027),
    .A3(net1051),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1617_));
 sky130_fd_sc_hd__mux4_2 _2672_ (.A0(net1043),
    .A1(net1032),
    .A2(net1008),
    .A3(net1022),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1618_));
 sky130_fd_sc_hd__mux2_4 _2673_ (.A0(_1617_),
    .A1(_1618_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_1619_));
 sky130_fd_sc_hd__mux4_2 _2674_ (.A0(net619),
    .A1(net1258),
    .A2(net191),
    .A3(net11),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1620_));
 sky130_fd_sc_hd__mux4_1 _2675_ (.A0(net59),
    .A1(net67),
    .A2(net93),
    .A3(net1220),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1621_));
 sky130_fd_sc_hd__mux2_4 _2676_ (.A0(_1620_),
    .A1(_1621_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_1622_));
 sky130_fd_sc_hd__mux2_4 _2677_ (.A0(_1622_),
    .A1(_1619_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__or2_1 _2678_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .B(net673),
    .X(_1623_));
 sky130_fd_sc_hd__a21oi_1 _2679_ (.A1(_0024_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_1624_));
 sky130_fd_sc_hd__mux2_1 _2680_ (.A0(net6),
    .A1(net22),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_1625_));
 sky130_fd_sc_hd__a221o_1 _2681_ (.A1(_1623_),
    .A2(_1624_),
    .B1(_1625_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_1626_));
 sky130_fd_sc_hd__mux2_1 _2682_ (.A0(net62),
    .A1(net78),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_1627_));
 sky130_fd_sc_hd__and2b_1 _2683_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .B(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(net98),
    .A1(net114),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_1629_));
 sky130_fd_sc_hd__a211o_1 _2685_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .A2(_1629_),
    .B1(_1628_),
    .C1(_0047_),
    .X(_1630_));
 sky130_fd_sc_hd__mux4_1 _2686_ (.A0(net1046),
    .A1(net1026),
    .A2(net1050),
    .A3(net1042),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_1631_));
 sky130_fd_sc_hd__or2_1 _2687_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .B(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__mux4_1 _2688_ (.A0(net1037),
    .A1(net1007),
    .A2(net1031),
    .A3(net1021),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_1633_));
 sky130_fd_sc_hd__o211a_1 _2689_ (.A1(_0047_),
    .A2(_1633_),
    .B1(_1632_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_1634_));
 sky130_fd_sc_hd__a31o_1 _2690_ (.A1(_0048_),
    .A2(_1626_),
    .A3(_1630_),
    .B1(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_1 _2691_ (.A0(_1635_),
    .A1(_0520_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ),
    .X(_1636_));
 sky130_fd_sc_hd__mux2_4 _2692_ (.A0(net1050),
    .A1(_0526_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ),
    .X(_1637_));
 sky130_fd_sc_hd__mux2_4 _2693_ (.A0(_1637_),
    .A1(_1636_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .A1(_0278_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ),
    .X(_1638_));
 sky130_fd_sc_hd__mux2_1 _2695_ (.A0(net1039),
    .A1(net965),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ),
    .X(_1639_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(_1639_),
    .A1(_1638_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2697_ (.A0(net1035),
    .A1(_0322_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .A3(_0346_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2698_ (.A0(net187),
    .A1(net198),
    .A2(net1255),
    .A3(net1042),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2699_ (.A0(net188),
    .A1(net199),
    .A2(net21),
    .A3(net1036),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2700_ (.A0(net185),
    .A1(net200),
    .A2(net114),
    .A3(net1006),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2701_ (.A0(net186),
    .A1(net113),
    .A2(net197),
    .A3(net695),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2702_ (.A0(net1053),
    .A1(_0407_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .A3(_0398_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2703_ (.A0(net1046),
    .A1(net1026),
    .A2(net1050),
    .A3(net1042),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_1640_));
 sky130_fd_sc_hd__mux4_1 _2704_ (.A0(net1036),
    .A1(net1006),
    .A2(net1031),
    .A3(net1054),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_1641_));
 sky130_fd_sc_hd__or2_1 _2705_ (.A(_0068_),
    .B(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__o21a_1 _2706_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_1640_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_1643_));
 sky130_fd_sc_hd__mux4_1 _2707_ (.A0(net1255),
    .A1(net98),
    .A2(net86),
    .A3(net114),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_1644_));
 sky130_fd_sc_hd__mux4_1 _2708_ (.A0(net186),
    .A1(net198),
    .A2(net4),
    .A3(net6),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_1645_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(_1644_),
    .A1(_1645_),
    .S(_0068_),
    .X(_1646_));
 sky130_fd_sc_hd__a22o_1 _2710_ (.A1(_1642_),
    .A2(_1643_),
    .B1(_1646_),
    .B2(_0069_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ));
 sky130_fd_sc_hd__mux4_2 _2711_ (.A0(net1042),
    .A1(_0526_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ),
    .A3(_0520_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2712_ (.A0(net1035),
    .A1(net965),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .A3(_0278_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2713_ (.A0(net1005),
    .A1(_0322_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .A3(_0346_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2714_ (.A0(net1255),
    .A1(net78),
    .A2(net63),
    .A3(net1010),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2715_ (.A0(net1256),
    .A1(net79),
    .A2(net64),
    .A3(net1048),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2716_ (.A0(net61),
    .A1(net114),
    .A2(net80),
    .A3(net1025),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2717_ (.A0(net62),
    .A1(net77),
    .A2(net113),
    .A3(net1053),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2718_ (.A0(net737),
    .A1(_0407_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(_0398_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2719_ (.A0(net1004),
    .A1(_0526_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .A3(_0520_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2720_ (.A0(net695),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A2(net965),
    .A3(_0278_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2721_ (.A0(net708),
    .A1(_0322_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .A3(_0346_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2722_ (.A0(net619),
    .A1(net1258),
    .A2(net1220),
    .A3(net1026),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_1647_));
 sky130_fd_sc_hd__mux4_1 _2723_ (.A0(net1006),
    .A1(_0704_),
    .A2(_0733_),
    .A3(_1498_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_1 _2724_ (.A0(_1647_),
    .A1(_1648_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2725_ (.A0(net618),
    .A1(net1219),
    .A2(net1257),
    .A3(net1050),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_1649_));
 sky130_fd_sc_hd__mux4_1 _2726_ (.A0(net1031),
    .A1(net721),
    .A2(_0652_),
    .A3(_1166_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_1650_));
 sky130_fd_sc_hd__mux2_1 _2727_ (.A0(_1649_),
    .A1(_1650_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _2728_ (.A0(net1022),
    .A1(net657),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_1651_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(net965),
    .A1(_0706_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_1652_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(_1651_),
    .A1(_1652_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .X(_1653_));
 sky130_fd_sc_hd__mux4_1 _2731_ (.A0(_0199_),
    .A1(net93),
    .A2(net1),
    .A3(net1043),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(_1654_),
    .A1(_1653_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ));
 sky130_fd_sc_hd__nor2_1 _2733_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .B(net1054),
    .Y(_1655_));
 sky130_fd_sc_hd__a211oi_1 _2734_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .A2(_1149_),
    .B1(_1655_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .Y(_1656_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(_1512_),
    .A1(_0737_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .X(_1657_));
 sky130_fd_sc_hd__a21bo_1 _2736_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .A2(_1657_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ),
    .X(_1658_));
 sky130_fd_sc_hd__mux4_1 _2737_ (.A0(_0243_),
    .A1(net94),
    .A2(net2),
    .A3(net1037),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .X(_1659_));
 sky130_fd_sc_hd__o22a_1 _2738_ (.A1(_1656_),
    .A2(_1658_),
    .B1(_1659_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2739_ (.A0(net621),
    .A1(net59),
    .A2(net1258),
    .A3(net1027),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_1660_));
 sky130_fd_sc_hd__mux4_1 _2740_ (.A0(net740),
    .A1(_0704_),
    .A2(_0733_),
    .A3(_0253_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_1661_));
 sky130_fd_sc_hd__mux2_1 _2741_ (.A0(_1660_),
    .A1(_1661_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2742_ (.A0(net1032),
    .A1(net721),
    .A2(_0652_),
    .A3(_1176_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_1662_));
 sky130_fd_sc_hd__mux4_1 _2743_ (.A0(net618),
    .A1(net1257),
    .A2(net60),
    .A3(net1051),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(_1663_),
    .A1(_1662_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2745_ (.A0(net744),
    .A1(net57),
    .A2(net1),
    .A3(net1043),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1664_));
 sky130_fd_sc_hd__mux2_1 _2746_ (.A0(net965),
    .A1(_0441_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1665_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(net1022),
    .A1(net657),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1666_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(_1666_),
    .A1(_1665_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ),
    .X(_1667_));
 sky130_fd_sc_hd__mux2_1 _2749_ (.A0(_1664_),
    .A1(_1667_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__nor2_1 _2750_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .B(net1055),
    .Y(_1668_));
 sky130_fd_sc_hd__a211oi_1 _2751_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .A2(_1149_),
    .B1(_1668_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .Y(_1669_));
 sky130_fd_sc_hd__mux2_1 _2752_ (.A0(_1512_),
    .A1(_0710_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1670_));
 sky130_fd_sc_hd__a21bo_1 _2753_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_1670_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ),
    .X(_1671_));
 sky130_fd_sc_hd__mux4_1 _2754_ (.A0(_0243_),
    .A1(net58),
    .A2(net2),
    .A3(net1038),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1672_));
 sky130_fd_sc_hd__o22a_1 _2755_ (.A1(_1669_),
    .A2(_1671_),
    .B1(_1672_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2756_ (.A0(_0733_),
    .A1(net622),
    .A2(_0704_),
    .A3(net965),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1673_));
 sky130_fd_sc_hd__nand2b_1 _2757_ (.A_N(_1673_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .Y(_1674_));
 sky130_fd_sc_hd__mux4_1 _2758_ (.A0(net740),
    .A1(net1032),
    .A2(net1022),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1675_));
 sky130_fd_sc_hd__o211a_1 _2759_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_1675_),
    .B1(_1674_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ),
    .X(_1676_));
 sky130_fd_sc_hd__nand2b_1 _2760_ (.A_N(net1219),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .Y(_1677_));
 sky130_fd_sc_hd__o21ba_1 _2761_ (.A1(net1257),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1678_));
 sky130_fd_sc_hd__mux2_1 _2762_ (.A0(net1012),
    .A1(net1047),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1679_));
 sky130_fd_sc_hd__a221o_1 _2763_ (.A1(_1677_),
    .A2(_1678_),
    .B1(_1679_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_1680_));
 sky130_fd_sc_hd__mux2_1 _2764_ (.A0(net1027),
    .A1(net1051),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1681_));
 sky130_fd_sc_hd__inv_1 _2765_ (.A(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__mux2_1 _2766_ (.A0(net1043),
    .A1(net1038),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1683_));
 sky130_fd_sc_hd__o21ai_1 _2767_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .A2(_1682_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .Y(_1684_));
 sky130_fd_sc_hd__a21o_1 _2768_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .A2(_1683_),
    .B1(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__a31o_1 _2769_ (.A1(_0148_),
    .A2(_1680_),
    .A3(_1685_),
    .B1(_1676_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux2_1 _2770_ (.A0(net721),
    .A1(_0652_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_1686_));
 sky130_fd_sc_hd__and2b_1 _2771_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .B(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__mux2_1 _2772_ (.A0(_1150_),
    .A1(_1512_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_1688_));
 sky130_fd_sc_hd__a21bo_1 _2773_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .A2(_1688_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .X(_1689_));
 sky130_fd_sc_hd__mux4_1 _2774_ (.A0(net1007),
    .A1(net1032),
    .A2(net1021),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_1690_));
 sky130_fd_sc_hd__o221a_1 _2775_ (.A1(_1687_),
    .A2(_1689_),
    .B1(_1690_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ),
    .X(_1691_));
 sky130_fd_sc_hd__mux4_1 _2776_ (.A0(net1258),
    .A1(net1012),
    .A2(net1220),
    .A3(net1047),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_1692_));
 sky130_fd_sc_hd__mux4_1 _2777_ (.A0(net1028),
    .A1(net1051),
    .A2(net1043),
    .A3(net1038),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_1693_));
 sky130_fd_sc_hd__inv_1 _2778_ (.A(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__a21oi_1 _2779_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_1694_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ),
    .Y(_1695_));
 sky130_fd_sc_hd__o21a_1 _2780_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_1692_),
    .B1(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__or2_1 _2781_ (.A(_1691_),
    .B(_1696_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2782_ (.A0(net621),
    .A1(net1258),
    .A2(net1220),
    .A3(net1025),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_1697_));
 sky130_fd_sc_hd__mux2_1 _2783_ (.A0(net1005),
    .A1(_0733_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_1698_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(_0704_),
    .A1(_1522_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_1699_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(_1698_),
    .A1(_1699_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_1700_));
 sky130_fd_sc_hd__mux2_2 _2786_ (.A0(_1697_),
    .A1(_1700_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2787_ (.A0(net618),
    .A1(net96),
    .A2(net1257),
    .A3(net1049),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_1701_));
 sky130_fd_sc_hd__mux4_1 _2788_ (.A0(net1030),
    .A1(net721),
    .A2(_0652_),
    .A3(_1139_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ),
    .X(_1702_));
 sky130_fd_sc_hd__mux2_2 _2789_ (.A0(_1701_),
    .A1(_1702_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2790_ (.A0(_0199_),
    .A1(net93),
    .A2(net1),
    .A3(net1041),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_1703_));
 sky130_fd_sc_hd__mux2_1 _2791_ (.A0(net676),
    .A1(net623),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_1704_));
 sky130_fd_sc_hd__mux2_1 _2792_ (.A0(net965),
    .A1(_0615_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_1705_));
 sky130_fd_sc_hd__mux2_1 _2793_ (.A0(_1704_),
    .A1(_1705_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .X(_1706_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(_1703_),
    .A1(_1706_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ));
 sky130_fd_sc_hd__nor2_1 _2795_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .B(net1054),
    .Y(_1707_));
 sky130_fd_sc_hd__a211oi_1 _2796_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .A2(_1149_),
    .B1(_1707_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .Y(_1708_));
 sky130_fd_sc_hd__mux2_1 _2797_ (.A0(_1512_),
    .A1(_0489_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .X(_1709_));
 sky130_fd_sc_hd__a21bo_1 _2798_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_1709_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ),
    .X(_1710_));
 sky130_fd_sc_hd__mux4_1 _2799_ (.A0(_0243_),
    .A1(net94),
    .A2(net2),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .X(_1711_));
 sky130_fd_sc_hd__o22a_1 _2800_ (.A1(_1708_),
    .A2(_1710_),
    .B1(_1711_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2801_ (.A0(net621),
    .A1(net59),
    .A2(net1220),
    .A3(net1028),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .X(_1712_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(_0704_),
    .A1(_1509_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_1713_));
 sky130_fd_sc_hd__nand2_1 _2803_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .B(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__mux2_1 _2804_ (.A0(net740),
    .A1(_0733_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_1715_));
 sky130_fd_sc_hd__inv_1 _2805_ (.A(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__o211a_1 _2806_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .A2(_1716_),
    .B1(_1714_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_1717_));
 sky130_fd_sc_hd__o21ba_1 _2807_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_1712_),
    .B1_N(_1717_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2808_ (.A0(net1031),
    .A1(net721),
    .A2(_0652_),
    .A3(_1147_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .X(_1718_));
 sky130_fd_sc_hd__mux4_1 _2809_ (.A0(net618),
    .A1(net1219),
    .A2(net60),
    .A3(net1050),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .X(_1719_));
 sky130_fd_sc_hd__mux2_1 _2810_ (.A0(_1719_),
    .A1(_1718_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _2811_ (.A0(net676),
    .A1(net623),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_1720_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(net965),
    .A1(_0634_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_1721_));
 sky130_fd_sc_hd__mux2_1 _2813_ (.A0(_1720_),
    .A1(_1721_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .X(_1722_));
 sky130_fd_sc_hd__mux4_1 _2814_ (.A0(net744),
    .A1(net93),
    .A2(net57),
    .A3(net1039),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_1723_));
 sky130_fd_sc_hd__mux2_1 _2815_ (.A0(_1723_),
    .A1(_1722_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__nor2_1 _2816_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .B(net1054),
    .Y(_1724_));
 sky130_fd_sc_hd__a211oi_1 _2817_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_1149_),
    .B1(_1724_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .Y(_1725_));
 sky130_fd_sc_hd__mux2_1 _2818_ (.A0(_1512_),
    .A1(_0540_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_1726_));
 sky130_fd_sc_hd__a21bo_1 _2819_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_1726_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_1727_));
 sky130_fd_sc_hd__mux4_1 _2820_ (.A0(_0243_),
    .A1(net94),
    .A2(net58),
    .A3(net1037),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_1728_));
 sky130_fd_sc_hd__o22a_1 _2821_ (.A1(_1725_),
    .A2(_1727_),
    .B1(_1728_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__nand2b_1 _2822_ (.A_N(net1219),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .Y(_1729_));
 sky130_fd_sc_hd__o21ba_1 _2823_ (.A1(net1257),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_1730_));
 sky130_fd_sc_hd__mux2_1 _2824_ (.A0(net1011),
    .A1(net1046),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_1731_));
 sky130_fd_sc_hd__a221o_1 _2825_ (.A1(_1729_),
    .A2(_1730_),
    .B1(_1731_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .X(_1732_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(net1026),
    .A1(net1050),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_1733_));
 sky130_fd_sc_hd__inv_1 _2827_ (.A(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__mux2_1 _2828_ (.A0(net1044),
    .A1(net1036),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_1735_));
 sky130_fd_sc_hd__o21ai_1 _2829_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .A2(_1734_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .Y(_1736_));
 sky130_fd_sc_hd__a21o_1 _2830_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .A2(_1735_),
    .B1(_1736_),
    .X(_1737_));
 sky130_fd_sc_hd__mux4_1 _2831_ (.A0(_0733_),
    .A1(net622),
    .A2(_0704_),
    .A3(net965),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_1738_));
 sky130_fd_sc_hd__nand2b_1 _2832_ (.A_N(_1738_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .Y(_1739_));
 sky130_fd_sc_hd__mux4_1 _2833_ (.A0(net1006),
    .A1(net1033),
    .A2(net1021),
    .A3(net1054),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_1740_));
 sky130_fd_sc_hd__o211a_1 _2834_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_1740_),
    .B1(_1739_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ),
    .X(_1741_));
 sky130_fd_sc_hd__a31o_1 _2835_ (.A1(_0149_),
    .A2(_1732_),
    .A3(_1737_),
    .B1(_1741_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux2_1 _2836_ (.A0(net721),
    .A1(_0652_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_1742_));
 sky130_fd_sc_hd__and2b_1 _2837_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .B(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__mux2_1 _2838_ (.A0(_1150_),
    .A1(_1512_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_1744_));
 sky130_fd_sc_hd__a21bo_1 _2839_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .A2(_1744_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .X(_1745_));
 sky130_fd_sc_hd__mux4_1 _2840_ (.A0(net1006),
    .A1(net1031),
    .A2(net1021),
    .A3(net1054),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .X(_1746_));
 sky130_fd_sc_hd__o221a_1 _2841_ (.A1(_1743_),
    .A2(_1745_),
    .B1(_1746_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ),
    .X(_1747_));
 sky130_fd_sc_hd__mux4_1 _2842_ (.A0(net1258),
    .A1(net1011),
    .A2(net1220),
    .A3(net1046),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_1748_));
 sky130_fd_sc_hd__mux4_1 _2843_ (.A0(net1026),
    .A1(net1050),
    .A2(net1042),
    .A3(net1036),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .X(_1749_));
 sky130_fd_sc_hd__inv_1 _2844_ (.A(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__a21oi_1 _2845_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_1750_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ),
    .Y(_1751_));
 sky130_fd_sc_hd__o21a_1 _2846_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_1748_),
    .B1(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__or2_1 _2847_ (.A(_1747_),
    .B(_1752_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2848_ (.A0(net1025),
    .A1(_0407_),
    .A2(_0468_),
    .A3(_0398_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2849_ (.A0(net179),
    .A1(net1215),
    .A2(net194),
    .A3(net743),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__mux4_1 _2850_ (.A0(net180),
    .A1(net139),
    .A2(net195),
    .A3(net983),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__mux4_1 _2851_ (.A0(net177),
    .A1(net196),
    .A2(net230),
    .A3(net997),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__mux4_1 _2852_ (.A0(net178),
    .A1(net193),
    .A2(net229),
    .A3(net1016),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__mux4_1 _2853_ (.A0(net990),
    .A1(_0196_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A3(_0173_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2854_ (.A0(net976),
    .A1(_0216_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .A3(_0230_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2855_ (.A0(net692),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .A2(net1003),
    .A3(_1327_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2856_ (.A0(net747),
    .A1(_0382_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A3(net688),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2857_ (.A0(net743),
    .A1(_0196_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .A3(_0173_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2858_ (.A0(net980),
    .A1(net995),
    .A2(net1016),
    .A3(net709),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_1753_));
 sky130_fd_sc_hd__mux4_1 _2859_ (.A0(net691),
    .A1(net985),
    .A2(net716),
    .A3(net743),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_1754_));
 sky130_fd_sc_hd__or2_1 _2860_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .B(_1754_),
    .X(_1755_));
 sky130_fd_sc_hd__o21a_1 _2861_ (.A1(_0150_),
    .A2(_1753_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_1756_));
 sky130_fd_sc_hd__mux4_1 _2862_ (.A0(net176),
    .A1(net178),
    .A2(net194),
    .A3(net142),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_1757_));
 sky130_fd_sc_hd__mux4_1 _2863_ (.A0(net1215),
    .A1(net214),
    .A2(net70),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_1758_));
 sky130_fd_sc_hd__mux2_1 _2864_ (.A0(_1757_),
    .A1(_1758_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_1759_));
 sky130_fd_sc_hd__a22o_1 _2865_ (.A1(_1755_),
    .A2(_1756_),
    .B1(_1759_),
    .B2(_0151_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2866_ (.A0(net715),
    .A1(_0216_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ),
    .A3(_0230_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ));
 sky130_fd_sc_hd__mux2_1 _2867_ (.A0(net747),
    .A1(_1361_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ),
    .X(_1760_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .A1(_1327_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ),
    .X(_1761_));
 sky130_fd_sc_hd__mux2_1 _2869_ (.A0(_1760_),
    .A1(_1761_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2870_ (.A0(net1016),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .A2(_0382_),
    .A3(net688),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2871_ (.A0(net1215),
    .A1(net82),
    .A2(net71),
    .A3(net972),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2872_ (.A0(net1216),
    .A1(net72),
    .A2(net83),
    .A3(net967),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2873_ (.A0(net69),
    .A1(net84),
    .A2(net230),
    .A3(net986),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2874_ (.A0(net70),
    .A1(net81),
    .A2(net229),
    .A3(net990),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2875_ (.A0(net715),
    .A1(_0196_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .A3(_0173_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2876_ (.A0(net729),
    .A1(net985),
    .A2(net716),
    .A3(net975),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_1762_));
 sky130_fd_sc_hd__or2_1 _2877_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .B(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__mux4_1 _2878_ (.A0(net981),
    .A1(net995),
    .A2(net1017),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_1764_));
 sky130_fd_sc_hd__o21a_1 _2879_ (.A1(_0152_),
    .A2(_1764_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_1765_));
 sky130_fd_sc_hd__mux4_1 _2880_ (.A0(net70),
    .A1(net82),
    .A2(net214),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_1766_));
 sky130_fd_sc_hd__mux4_1 _2881_ (.A0(net202),
    .A1(net1217),
    .A2(net124),
    .A3(net1215),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_1767_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(_1766_),
    .A1(_1767_),
    .S(_0152_),
    .X(_1768_));
 sky130_fd_sc_hd__a22o_1 _2883_ (.A1(_1763_),
    .A2(_1765_),
    .B1(_1768_),
    .B2(_0153_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2884_ (.A0(net995),
    .A1(_0216_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ),
    .A3(_0230_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(net1017),
    .A1(net1003),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ),
    .X(_1769_));
 sky130_fd_sc_hd__mux2_1 _2886_ (.A0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .A1(_1327_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ),
    .X(_1770_));
 sky130_fd_sc_hd__mux2_1 _2887_ (.A0(_1769_),
    .A1(_1770_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2888_ (.A0(net971),
    .A1(_0382_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .A3(net688),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _2889_ (.A0(net175),
    .A1(net1218),
    .A2(net1068),
    .A3(net987),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ),
    .X(_1771_));
 sky130_fd_sc_hd__mux2_1 _2890_ (.A0(net997),
    .A1(_0767_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .X(_1772_));
 sky130_fd_sc_hd__and2b_1 _2891_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ),
    .B(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__mux2_1 _2892_ (.A0(_0940_),
    .A1(_1364_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .X(_1774_));
 sky130_fd_sc_hd__a21bo_1 _2893_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ),
    .A2(_1774_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ),
    .X(_1775_));
 sky130_fd_sc_hd__o22a_1 _2894_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ),
    .A2(_1771_),
    .B1(_1773_),
    .B2(_1775_),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__mux4_1 _2895_ (.A0(net176),
    .A1(net1217),
    .A2(net1067),
    .A3(net716),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_1776_));
 sky130_fd_sc_hd__mux2_1 _2896_ (.A0(_0818_),
    .A1(_1421_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .X(_1777_));
 sky130_fd_sc_hd__nor2_1 _2897_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .B(net733),
    .Y(_1778_));
 sky130_fd_sc_hd__a211o_1 _2898_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .A2(_0662_),
    .B1(_1778_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_1779_));
 sky130_fd_sc_hd__a21bo_1 _2899_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_1777_),
    .B1_N(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__mux2_1 _2900_ (.A0(_1776_),
    .A1(_1780_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__mux4_1 _2901_ (.A0(net173),
    .A1(net119),
    .A2(net209),
    .A3(net979),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_1781_));
 sky130_fd_sc_hd__mux2_1 _2902_ (.A0(net1003),
    .A1(_0921_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .X(_1782_));
 sky130_fd_sc_hd__mux2_1 _2903_ (.A0(net1001),
    .A1(_1429_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .X(_1783_));
 sky130_fd_sc_hd__mux2_1 _2904_ (.A0(_1783_),
    .A1(_1782_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_1784_));
 sky130_fd_sc_hd__mux2_1 _2905_ (.A0(_1781_),
    .A1(_1784_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__mux4_1 _2906_ (.A0(net174),
    .A1(net210),
    .A2(net120),
    .A3(net983),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ),
    .X(_1785_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(_1349_),
    .A1(_0781_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ),
    .X(_1786_));
 sky130_fd_sc_hd__mux2_1 _2908_ (.A0(net1014),
    .A1(_1410_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ),
    .X(_1787_));
 sky130_fd_sc_hd__inv_1 _2909_ (.A(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__o21ai_1 _2910_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_1788_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ),
    .Y(_1789_));
 sky130_fd_sc_hd__a21o_1 _2911_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_1786_),
    .B1(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__o21a_1 _2912_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ),
    .A2(_1785_),
    .B1(_1790_),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__mux4_1 _2913_ (.A0(net175),
    .A1(net1218),
    .A2(_0302_),
    .A3(net989),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .X(_1791_));
 sky130_fd_sc_hd__mux4_1 _2914_ (.A0(net998),
    .A1(_0767_),
    .A2(_0940_),
    .A3(_1382_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .X(_1792_));
 sky130_fd_sc_hd__mux2_1 _2915_ (.A0(_1791_),
    .A1(_1792_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(_0818_),
    .A1(_1437_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .X(_1793_));
 sky130_fd_sc_hd__nand2_1 _2917_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .B(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__nor2_1 _2918_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .B(net733),
    .Y(_1795_));
 sky130_fd_sc_hd__a211o_1 _2919_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .A2(_0662_),
    .B1(_1795_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_1796_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(_0350_),
    .A1(net990),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .X(_1797_));
 sky130_fd_sc_hd__mux2_1 _2921_ (.A0(net176),
    .A1(net1217),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .X(_1798_));
 sky130_fd_sc_hd__a21o_1 _2922_ (.A1(_0154_),
    .A2(_1798_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_1799_));
 sky130_fd_sc_hd__a21oi_1 _2923_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(_1797_),
    .B1(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__a31oi_1 _2924_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ),
    .A2(_1794_),
    .A3(_1796_),
    .B1(_1800_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__mux4_2 _2925_ (.A0(net173),
    .A1(net119),
    .A2(_0410_),
    .A3(net979),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ),
    .X(_1801_));
 sky130_fd_sc_hd__mux2_1 _2926_ (.A0(net1003),
    .A1(_0968_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .X(_1802_));
 sky130_fd_sc_hd__mux2_1 _2927_ (.A0(net1000),
    .A1(_1429_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .X(_1803_));
 sky130_fd_sc_hd__mux2_1 _2928_ (.A0(_1803_),
    .A1(_1802_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ),
    .X(_1804_));
 sky130_fd_sc_hd__mux2_2 _2929_ (.A0(_1801_),
    .A1(_1804_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__nand2b_1 _2930_ (.A_N(_0860_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .Y(_1805_));
 sky130_fd_sc_hd__o211a_1 _2931_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(_1349_),
    .B1(_1805_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1806_));
 sky130_fd_sc_hd__mux2_4 _2932_ (.A0(net1015),
    .A1(_1410_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .X(_1807_));
 sky130_fd_sc_hd__inv_1 _2933_ (.A(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__o21ai_1 _2934_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_1808_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ),
    .Y(_1809_));
 sky130_fd_sc_hd__mux4_2 _2935_ (.A0(net174),
    .A1(net120),
    .A2(_0529_),
    .A3(net984),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_1810_));
 sky130_fd_sc_hd__o22a_4 _2936_ (.A1(_1806_),
    .A2(_1809_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ),
    .B2(_1810_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__nand2b_1 _2937_ (.A_N(net212),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .Y(_1811_));
 sky130_fd_sc_hd__o21ba_1 _2938_ (.A1(net1217),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1812_));
 sky130_fd_sc_hd__mux2_1 _2939_ (.A0(net972),
    .A1(net967),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_1813_));
 sky130_fd_sc_hd__a221o_1 _2940_ (.A1(_1811_),
    .A2(_1812_),
    .B1(_1813_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_1814_));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(net986),
    .A1(net990),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_1815_));
 sky130_fd_sc_hd__inv_1 _2942_ (.A(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__mux2_1 _2943_ (.A0(net976),
    .A1(net692),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_1817_));
 sky130_fd_sc_hd__o21ai_1 _2944_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .A2(_1816_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .Y(_1818_));
 sky130_fd_sc_hd__a21o_1 _2945_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .A2(_1817_),
    .B1(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__mux4_1 _2946_ (.A0(_0767_),
    .A1(_0940_),
    .A2(_1429_),
    .A3(net1003),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1820_));
 sky130_fd_sc_hd__nand2b_1 _2947_ (.A_N(_1820_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .Y(_1821_));
 sky130_fd_sc_hd__mux4_1 _2948_ (.A0(net999),
    .A1(net1018),
    .A2(net693),
    .A3(net709),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_1822_));
 sky130_fd_sc_hd__o211a_1 _2949_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_1822_),
    .B1(_1821_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ),
    .X(_1823_));
 sky130_fd_sc_hd__a31o_1 _2950_ (.A1(_0155_),
    .A2(_1814_),
    .A3(_1819_),
    .B1(_1823_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(_0662_),
    .A1(_0819_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1824_));
 sky130_fd_sc_hd__mux2_1 _2952_ (.A0(_1410_),
    .A1(_1349_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1825_));
 sky130_fd_sc_hd__nand2_1 _2953_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__o211a_1 _2954_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .A2(_1824_),
    .B1(_1826_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_1827_));
 sky130_fd_sc_hd__mux4_1 _2955_ (.A0(net747),
    .A1(net733),
    .A2(net693),
    .A3(net709),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1828_));
 sky130_fd_sc_hd__o21ai_1 _2956_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_1828_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ),
    .Y(_1829_));
 sky130_fd_sc_hd__mux4_1 _2957_ (.A0(net1218),
    .A1(net1068),
    .A2(net972),
    .A3(net967),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_1830_));
 sky130_fd_sc_hd__nor2_1 _2958_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .B(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__mux4_1 _2959_ (.A0(net986),
    .A1(net976),
    .A2(net990),
    .A3(net692),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_1832_));
 sky130_fd_sc_hd__inv_1 _2960_ (.A(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__a211o_1 _2961_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_1833_),
    .B1(_1831_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ),
    .X(_1834_));
 sky130_fd_sc_hd__o21ai_1 _2962_ (.A1(_1827_),
    .A2(_1829_),
    .B1(_1834_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2963_ (.A0(net175),
    .A1(net1218),
    .A2(net1068),
    .A3(net986),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_1 _2964_ (.A0(net996),
    .A1(_0767_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(_0940_),
    .A1(_1329_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .X(_1837_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(_1836_),
    .A1(_1837_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ),
    .X(_1838_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(_1835_),
    .A1(_1838_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _2968_ (.A0(net176),
    .A1(net1217),
    .A2(net1067),
    .A3(net994),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_1839_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(_0818_),
    .A1(_1391_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .X(_1840_));
 sky130_fd_sc_hd__nor2_1 _2970_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .B(net734),
    .Y(_1841_));
 sky130_fd_sc_hd__a211o_1 _2971_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .A2(_0662_),
    .B1(_1841_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_1842_));
 sky130_fd_sc_hd__a21bo_1 _2972_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_1840_),
    .B1_N(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(_1839_),
    .A1(_1843_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _2974_ (.A0(net173),
    .A1(net119),
    .A2(net209),
    .A3(net976),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_1844_));
 sky130_fd_sc_hd__mux2_1 _2975_ (.A0(net1003),
    .A1(_0571_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .X(_1845_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(net693),
    .A1(_1429_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_1 _2977_ (.A0(_1846_),
    .A1(_1845_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_1847_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(_1844_),
    .A1(_1847_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _2979_ (.A0(net174),
    .A1(net210),
    .A2(net120),
    .A3(net692),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_1848_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(_1349_),
    .A1(_0598_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_1849_));
 sky130_fd_sc_hd__mux2_1 _2981_ (.A0(net709),
    .A1(_1410_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_1850_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(_1850_),
    .A1(_1849_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_1851_));
 sky130_fd_sc_hd__mux2_1 _2983_ (.A0(_1848_),
    .A1(_1851_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(net997),
    .A1(_0767_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .X(_1852_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(_0940_),
    .A1(_1347_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .X(_1853_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(_1852_),
    .A1(_1853_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .X(_1854_));
 sky130_fd_sc_hd__mux4_1 _2987_ (.A0(net175),
    .A1(net1068),
    .A2(_0302_),
    .A3(net988),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .X(_1855_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(_1855_),
    .A1(_1854_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(_0818_),
    .A1(_1408_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .X(_1856_));
 sky130_fd_sc_hd__nand2_1 _2990_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .B(_0662_),
    .Y(_1857_));
 sky130_fd_sc_hd__o21ba_1 _2991_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .A2(net733),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_1858_));
 sky130_fd_sc_hd__a221o_1 _2992_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_1856_),
    .B1(_1857_),
    .B2(_1858_),
    .C1(_0156_),
    .X(_1859_));
 sky130_fd_sc_hd__mux4_1 _2993_ (.A0(net176),
    .A1(net1067),
    .A2(_0350_),
    .A3(net990),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .X(_1860_));
 sky130_fd_sc_hd__o21a_1 _2994_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ),
    .A2(_1860_),
    .B1(_1859_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _2995_ (.A0(net1003),
    .A1(_0802_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_1861_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(net714),
    .A1(_1429_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_1862_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(_1862_),
    .A1(_1861_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .X(_1863_));
 sky130_fd_sc_hd__mux4_1 _2998_ (.A0(net173),
    .A1(net209),
    .A2(_0410_),
    .A3(net977),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_1864_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(_1864_),
    .A1(_1863_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux4_2 _3000_ (.A0(net174),
    .A1(net210),
    .A2(_0529_),
    .A3(net983),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .X(_1865_));
 sky130_fd_sc_hd__mux2_2 _3001_ (.A0(_1349_),
    .A1(_0672_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .X(_1866_));
 sky130_fd_sc_hd__mux2_4 _3002_ (.A0(net1014),
    .A1(_1410_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .X(_1867_));
 sky130_fd_sc_hd__inv_1 _3003_ (.A(_1867_),
    .Y(_1868_));
 sky130_fd_sc_hd__o21ai_1 _3004_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_1868_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ),
    .Y(_1869_));
 sky130_fd_sc_hd__a21o_1 _3005_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_1866_),
    .B1(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__o21a_1 _3006_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_1865_),
    .B1(_1870_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__nand2b_1 _3007_ (.A_N(net1067),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .Y(_1871_));
 sky130_fd_sc_hd__o21ba_1 _3008_ (.A1(net122),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_1872_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(net974),
    .A1(net969),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_1873_));
 sky130_fd_sc_hd__a221o_1 _3010_ (.A1(_1871_),
    .A2(_1872_),
    .B1(_1873_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_1874_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(net988),
    .A1(net993),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_1875_));
 sky130_fd_sc_hd__inv_1 _3012_ (.A(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__mux2_1 _3013_ (.A0(net978),
    .A1(net983),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_1877_));
 sky130_fd_sc_hd__o21ai_1 _3014_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_1876_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .Y(_1878_));
 sky130_fd_sc_hd__a21o_1 _3015_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_1877_),
    .B1(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__mux4_1 _3016_ (.A0(_0767_),
    .A1(_0940_),
    .A2(_1429_),
    .A3(net1003),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_1880_));
 sky130_fd_sc_hd__nand2b_1 _3017_ (.A_N(_1880_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .Y(_1881_));
 sky130_fd_sc_hd__mux4_1 _3018_ (.A0(net997),
    .A1(net1019),
    .A2(net1002),
    .A3(net1014),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_1882_));
 sky130_fd_sc_hd__o211a_1 _3019_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_1882_),
    .B1(_1881_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_1883_));
 sky130_fd_sc_hd__a31o_1 _3020_ (.A1(_0157_),
    .A2(_1874_),
    .A3(_1879_),
    .B1(_1883_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux2_2 _3021_ (.A0(_0662_),
    .A1(_0819_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_1884_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(_1410_),
    .A1(_1349_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_1885_));
 sky130_fd_sc_hd__nand2_1 _3023_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .B(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__o211a_1 _3024_ (.A1(_1884_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .B1(_1886_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .X(_1887_));
 sky130_fd_sc_hd__mux4_1 _3025_ (.A0(net995),
    .A1(net1016),
    .A2(net714),
    .A3(net709),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_1888_));
 sky130_fd_sc_hd__o21ai_1 _3026_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_1888_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ),
    .Y(_1889_));
 sky130_fd_sc_hd__mux4_1 _3027_ (.A0(net1218),
    .A1(net1068),
    .A2(net971),
    .A3(net691),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_1890_));
 sky130_fd_sc_hd__nor2_1 _3028_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .B(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__mux4_1 _3029_ (.A0(net707),
    .A1(net743),
    .A2(net716),
    .A3(net980),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_1892_));
 sky130_fd_sc_hd__inv_1 _3030_ (.A(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__a211o_1 _3031_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_1893_),
    .B1(_1891_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ),
    .X(_1894_));
 sky130_fd_sc_hd__o21ai_2 _3032_ (.A1(_1889_),
    .A2(_1887_),
    .B1(_1894_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__nor2_1 _3033_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .Y(_1895_));
 sky130_fd_sc_hd__mux4_1 _3034_ (.A0(net191),
    .A1(net131),
    .A2(net137),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_1896_));
 sky130_fd_sc_hd__mux4_1 _3035_ (.A0(net221),
    .A1(net658),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .X(_1897_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(_1896_),
    .A1(_1897_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_1898_));
 sky130_fd_sc_hd__o21ai_1 _3037_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .Y(_1899_));
 sky130_fd_sc_hd__o31a_1 _3038_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .A3(_0183_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_1900_));
 sky130_fd_sc_hd__nand2_1 _3039_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .B(net703),
    .Y(_1901_));
 sky130_fd_sc_hd__o211a_1 _3040_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .B1(_1901_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_1902_));
 sky130_fd_sc_hd__and3b_1 _3041_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .X(_1903_));
 sky130_fd_sc_hd__a211o_1 _3042_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .A2(_1895_),
    .B1(_1902_),
    .C1(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__o2bb2a_1 _3043_ (.A1_N(_1899_),
    .A2_N(_1900_),
    .B1(_1904_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_1905_));
 sky130_fd_sc_hd__mux2_1 _3044_ (.A0(_1898_),
    .A1(_1905_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ));
 sky130_fd_sc_hd__and2b_1 _3045_ (.A_N(net963),
    .B(_1466_),
    .X(_0000_));
 sky130_fd_sc_hd__and2b_1 _3046_ (.A_N(net963),
    .B(_1615_),
    .X(_0001_));
 sky130_fd_sc_hd__and2b_1 _3047_ (.A_N(net963),
    .B(_1464_),
    .X(_0002_));
 sky130_fd_sc_hd__and2b_1 _3048_ (.A_N(net963),
    .B(_1468_),
    .X(_0003_));
 sky130_fd_sc_hd__and2b_1 _3049_ (.A_N(net963),
    .B(_1467_),
    .X(_0004_));
 sky130_fd_sc_hd__and2b_1 _3050_ (.A_N(net963),
    .B(_1469_),
    .X(_0005_));
 sky130_fd_sc_hd__and2b_1 _3051_ (.A_N(net963),
    .B(_1470_),
    .X(_0006_));
 sky130_fd_sc_hd__and2b_1 _3052_ (.A_N(net963),
    .B(_1471_),
    .X(_0007_));
 sky130_fd_sc_hd__and2b_1 _3053_ (.A_N(net963),
    .B(_1616_),
    .X(_0008_));
 sky130_fd_sc_hd__and2b_1 _3054_ (.A_N(net963),
    .B(_1473_),
    .X(_0009_));
 sky130_fd_sc_hd__and2b_1 _3055_ (.A_N(net964),
    .B(_1475_),
    .X(_0010_));
 sky130_fd_sc_hd__nor2_1 _3056_ (.A(net964),
    .B(_1476_),
    .Y(_0011_));
 sky130_fd_sc_hd__and2b_1 _3057_ (.A_N(net964),
    .B(_1478_),
    .X(_0012_));
 sky130_fd_sc_hd__and2b_1 _3058_ (.A_N(net964),
    .B(_1613_),
    .X(_0013_));
 sky130_fd_sc_hd__and2b_1 _3059_ (.A_N(net964),
    .B(_1462_),
    .X(_0014_));
 sky130_fd_sc_hd__and2b_1 _3060_ (.A_N(net964),
    .B(_1505_),
    .X(_0015_));
 sky130_fd_sc_hd__and2b_1 _3061_ (.A_N(net964),
    .B(_1520_),
    .X(_0016_));
 sky130_fd_sc_hd__and2b_1 _3062_ (.A_N(net964),
    .B(_1548_),
    .X(_0017_));
 sky130_fd_sc_hd__and2b_1 _3063_ (.A_N(net964),
    .B(_1614_),
    .X(_0018_));
 sky130_fd_sc_hd__and2b_1 _3064_ (.A_N(net964),
    .B(_1611_),
    .X(_0019_));
 sky130_fd_sc_hd__inv_2 _3065_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_1 _3066_ (.A(net139),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_1 _3068_ (.A(net189),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _3069_ (.A(net186),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_1 _3070_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _3071_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_1 _3072_ (.A(net222),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _3073_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _3074_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_1 _3075_ (.A(net73),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _3076_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_1 _3077_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _3078_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _3079_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _3080_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_1 _3081_ (.A(net185),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _3082_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _3083_ (.A(net228),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _3084_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _3085_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _3086_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _3087_ (.A(net188),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _3088_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _3089_ (.A(net20),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _3090_ (.A(net76),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_1 _3091_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _3092_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_1 _3093_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_1 _3094_ (.A(net187),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _3095_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_1 _3096_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _3097_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _3098_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _3099_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _3100_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _3101_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _3102_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _3103_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _3104_ (.A(net75),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _3105_ (.A(net18),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _3106_ (.A(net74),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _3107_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_1 _3108_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _3109_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_1 _3110_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_1 _3111_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_1 _3112_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _3113_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_1 _3114_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _3115_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_1 _3116_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _3117_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _3118_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _3119_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _3120_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _3121_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _3122_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_1 _3123_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _3124_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_1 _3125_ (.A(net17),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_1 _3126_ (.A(net109),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _3127_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_1 _3128_ (.A(net19),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _3129_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _3130_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_1 _3131_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _3132_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _3133_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_1 _3134_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_1 _3135_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _3136_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _3137_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _3138_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _3139_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _3140_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _3141_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _3142_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _3143_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _3144_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_1 _3145_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_1 _3146_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_1 _3147_ (.A(net135),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_1 _3148_ (.A(net225),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_1 _3149_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_1 _3150_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _3151_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _3152_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _3153_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_1 _3154_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _3155_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_1 _3156_ (.A(net213),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_1 _3157_ (.A(net201),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_1 _3158_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_1 _3159_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _3160_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _3161_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _3162_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_1 _3163_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_1 _3164_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _3165_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _3166_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _3167_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _3168_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_1 _3169_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _3170_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_1 _3171_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_1 _3172_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _3173_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_1 _3174_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_1 _3175_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _3176_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_1 _3177_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_1 _3178_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_1 _3179_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_1 _3180_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_1 _3181_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_1 _3182_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_1 _3183_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_1 _3184_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _3185_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _3186_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _3187_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _3188_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_1 _3189_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _3190_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _3191_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_1 _3192_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_1 _3193_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_1 _3194_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_1 _3195_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_1 _3196_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _3197_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_1 _3198_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_1 _3199_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_1 _3200_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_1 _3201_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_1 _3202_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_1 _3203_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .Y(_0158_));
 sky130_fd_sc_hd__mux4_1 _3204_ (.A0(net1011),
    .A1(net1046),
    .A2(net1026),
    .A3(net1050),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _3205_ (.A(_0085_),
    .B(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__mux4_1 _3206_ (.A0(net1036),
    .A1(net1006),
    .A2(net1031),
    .A3(net1054),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0161_));
 sky130_fd_sc_hd__a21bo_1 _3207_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0161_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0162_));
 sky130_fd_sc_hd__mux4_2 _3208_ (.A0(net971),
    .A1(net966),
    .A2(net991),
    .A3(net977),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0163_));
 sky130_fd_sc_hd__or2_4 _3209_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .B(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__mux4_2 _3210_ (.A0(net981),
    .A1(net730),
    .A2(net1017),
    .A3(net1013),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0165_));
 sky130_fd_sc_hd__o21a_1 _3211_ (.A1(_0165_),
    .A2(_0033_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0166_));
 sky130_fd_sc_hd__mux4_1 _3212_ (.A0(net140),
    .A1(net72),
    .A2(net216),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0167_));
 sky130_fd_sc_hd__mux4_1 _3213_ (.A0(net174),
    .A1(net180),
    .A2(net196),
    .A3(net126),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _3214_ (.A0(_0167_),
    .A1(_0168_),
    .S(_0033_),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _3215_ (.A1(_0164_),
    .A2(_0166_),
    .B1(_0169_),
    .B2(_0034_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__a221o_1 _3216_ (.A1(_0166_),
    .A2(_0164_),
    .B1(_0169_),
    .B2(_0034_),
    .C1(_0032_),
    .X(_0170_));
 sky130_fd_sc_hd__o21a_1 _3217_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .A2(net220),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(net195),
    .A1(net125),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_0172_));
 sky130_fd_sc_hd__a22o_4 _3219_ (.A1(_0171_),
    .A2(_0170_),
    .B1(_0172_),
    .B2(_0035_),
    .X(_0173_));
 sky130_fd_sc_hd__a221o_1 _3220_ (.A1(_0170_),
    .A2(_0171_),
    .B1(_0172_),
    .B2(_0035_),
    .C1(_0029_),
    .X(_0174_));
 sky130_fd_sc_hd__mux4_2 _3221_ (.A0(net981),
    .A1(net995),
    .A2(net1017),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0175_));
 sky130_fd_sc_hd__nor2_2 _3222_ (.A(_0031_),
    .B(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__mux4_2 _3223_ (.A0(net971),
    .A1(net727),
    .A2(net707),
    .A3(net977),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0177_));
 sky130_fd_sc_hd__o21ai_2 _3224_ (.A1(_0177_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .Y(_0178_));
 sky130_fd_sc_hd__mux4_1 _3225_ (.A0(net175),
    .A1(net181),
    .A2(net127),
    .A3(net1216),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0179_));
 sky130_fd_sc_hd__nor2_1 _3226_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .B(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__mux4_1 _3227_ (.A0(net73),
    .A1(net81),
    .A2(net217),
    .A3(net229),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0181_));
 sky130_fd_sc_hd__nor2_1 _3228_ (.A(_0031_),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__o32a_4 _3229_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .A2(_0180_),
    .A3(_0182_),
    .B1(_0178_),
    .B2(_0176_),
    .X(_0183_));
 sky130_fd_sc_hd__inv_1 _3230_ (.A(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__a21boi_4 _3231_ (.A1(_0183_),
    .A2(_0029_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ),
    .Y(_0185_));
 sky130_fd_sc_hd__mux4_2 _3232_ (.A0(net1009),
    .A1(net1024),
    .A2(net713),
    .A3(net1039),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0186_));
 sky130_fd_sc_hd__or2_4 _3233_ (.A(_0186_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0187_));
 sky130_fd_sc_hd__mux4_1 _3234_ (.A0(net1034),
    .A1(net1004),
    .A2(net1029),
    .A3(net1023),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0188_));
 sky130_fd_sc_hd__o21a_1 _3235_ (.A1(_0025_),
    .A2(_0188_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0189_));
 sky130_fd_sc_hd__mux4_1 _3236_ (.A0(net207),
    .A1(net1),
    .A2(net25),
    .A3(net1256),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0190_));
 sky130_fd_sc_hd__mux4_1 _3237_ (.A0(net79),
    .A1(net87),
    .A2(net99),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _3238_ (.A0(_0190_),
    .A1(_0191_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0192_));
 sky130_fd_sc_hd__a22o_4 _3239_ (.A1(_0189_),
    .A2(_0187_),
    .B1(_0192_),
    .B2(_0026_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ));
 sky130_fd_sc_hd__a221o_1 _3240_ (.A1(_0187_),
    .A2(_0189_),
    .B1(_0192_),
    .B2(_0026_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .X(_0193_));
 sky130_fd_sc_hd__a21oi_1 _3241_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .A2(_0027_),
    .B1(_0028_),
    .Y(_0194_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(net186),
    .A1(net132),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_2 _3243_ (.A1(_0193_),
    .A2(_0194_),
    .B1(_0195_),
    .B2(_0028_),
    .X(_0196_));
 sky130_fd_sc_hd__a221o_1 _3244_ (.A1(_0193_),
    .A2(_0194_),
    .B1(_0195_),
    .B2(_0028_),
    .C1(_0029_),
    .X(_0197_));
 sky130_fd_sc_hd__o21ba_1 _3245_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(net988),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0198_));
 sky130_fd_sc_hd__a22o_4 _3246_ (.A1(net745),
    .A2(net725),
    .B1(_0197_),
    .B2(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__a221o_1 _3247_ (.A1(_0185_),
    .A2(_0174_),
    .B1(_0197_),
    .B2(_0198_),
    .C1(net617),
    .X(_0200_));
 sky130_fd_sc_hd__a21oi_1 _3248_ (.A1(_0036_),
    .A2(net617),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0201_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(net1),
    .A1(net5),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0202_));
 sky130_fd_sc_hd__a21o_1 _3250_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0202_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0203_));
 sky130_fd_sc_hd__a21o_1 _3251_ (.A1(_0201_),
    .A2(_0200_),
    .B1(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__mux4_1 _3252_ (.A0(net57),
    .A1(net61),
    .A2(net93),
    .A3(net1220),
    .S0(net617),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0205_));
 sky130_fd_sc_hd__o21ba_1 _3253_ (.A1(_0037_),
    .A2(_0205_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_0206_));
 sky130_fd_sc_hd__nand2b_1 _3254_ (.A_N(net1034),
    .B(net617),
    .Y(_0207_));
 sky130_fd_sc_hd__o21ba_1 _3255_ (.A1(net617),
    .A2(net1039),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(net1004),
    .A1(net1023),
    .S(net617),
    .X(_0209_));
 sky130_fd_sc_hd__a221o_1 _3257_ (.A1(_0207_),
    .A2(_0208_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .B2(_0209_),
    .C1(_0037_),
    .X(_0210_));
 sky130_fd_sc_hd__mux4_2 _3258_ (.A0(net1009),
    .A1(net1045),
    .A2(net1024),
    .A3(net1049),
    .S0(net617),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0211_));
 sky130_fd_sc_hd__o211a_1 _3259_ (.A1(_0211_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .B1(_0210_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_0212_));
 sky130_fd_sc_hd__a21o_4 _3260_ (.A1(_0206_),
    .A2(_0204_),
    .B1(_0212_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ));
 sky130_fd_sc_hd__a211o_1 _3261_ (.A1(_0204_),
    .A2(_0206_),
    .B1(_0212_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0213_));
 sky130_fd_sc_hd__a21oi_1 _3262_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .A2(_0038_),
    .B1(_0039_),
    .Y(_0214_));
 sky130_fd_sc_hd__mux2_1 _3263_ (.A0(net192),
    .A1(net138),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_4 _3264_ (.A1(_0213_),
    .A2(_0214_),
    .B1(_0215_),
    .B2(_0039_),
    .X(_0216_));
 sky130_fd_sc_hd__a221o_1 _3265_ (.A1(net711),
    .A2(_0214_),
    .B1(_0215_),
    .B2(_0039_),
    .C1(_0040_),
    .X(_0217_));
 sky130_fd_sc_hd__o21ba_1 _3266_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .A2(net993),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ),
    .X(_0218_));
 sky130_fd_sc_hd__mux4_2 _3267_ (.A0(net971),
    .A1(net691),
    .A2(net707),
    .A3(net743),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0219_));
 sky130_fd_sc_hd__and2b_1 _3268_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__mux4_2 _3269_ (.A0(net715),
    .A1(net995),
    .A2(net1016),
    .A3(net1013),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0221_));
 sky130_fd_sc_hd__a21bo_1 _3270_ (.A1(_0221_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0222_));
 sky130_fd_sc_hd__mux4_1 _3271_ (.A0(net181),
    .A1(net127),
    .A2(net1218),
    .A3(net1216),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0223_));
 sky130_fd_sc_hd__and2b_1 _3272_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(net73),
    .A1(net81),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0225_));
 sky130_fd_sc_hd__and2b_1 _3274_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .B(net217),
    .X(_0226_));
 sky130_fd_sc_hd__a21bo_1 _3275_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .A2(net233),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0227_));
 sky130_fd_sc_hd__o221a_1 _3276_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_0225_),
    .B1(_0226_),
    .B2(_0227_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0228_));
 sky130_fd_sc_hd__o32a_4 _3277_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0224_),
    .A3(_0228_),
    .B1(_0222_),
    .B2(_0220_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__inv_2 _3278_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .Y(_0229_));
 sky130_fd_sc_hd__mux4_2 _3279_ (.A0(net194),
    .A1(net90),
    .A2(net217),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0230_));
 sky130_fd_sc_hd__mux4_1 _3280_ (.A0(net983),
    .A1(net997),
    .A2(net1019),
    .A3(net1014),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0231_));
 sky130_fd_sc_hd__mux4_2 _3281_ (.A0(net969),
    .A1(net988),
    .A2(net993),
    .A3(net978),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_4 _3282_ (.A0(_0231_),
    .A1(_0232_),
    .S(_0041_),
    .X(_0233_));
 sky130_fd_sc_hd__and2b_1 _3283_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .B(net214),
    .X(_0234_));
 sky130_fd_sc_hd__a21bo_1 _3284_ (.A1(net230),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _3285_ (.A0(net70),
    .A1(net82),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0236_));
 sky130_fd_sc_hd__o221a_1 _3286_ (.A1(_0234_),
    .A2(_0235_),
    .B1(_0236_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0237_));
 sky130_fd_sc_hd__mux4_1 _3287_ (.A0(net176),
    .A1(net178),
    .A2(net124),
    .A3(net1215),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0238_));
 sky130_fd_sc_hd__a21o_1 _3288_ (.A1(_0041_),
    .A2(_0238_),
    .B1(_0237_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_2 _3289_ (.A0(_0239_),
    .A1(_0233_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0240_));
 sky130_fd_sc_hd__or2_4 _3290_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .B(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__o211a_4 _3291_ (.A1(_0040_),
    .A2(_0230_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ),
    .C1(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__a21o_4 _3292_ (.A1(net663),
    .A2(_0218_),
    .B1(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _3293_ (.A0(_0243_),
    .A1(net190),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _3294_ (.A0(net2),
    .A1(net10),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0245_));
 sky130_fd_sc_hd__or2_1 _3295_ (.A(_0084_),
    .B(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__o211a_1 _3296_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .A2(_0244_),
    .B1(_0246_),
    .C1(_0085_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _3297_ (.A0(net58),
    .A1(net66),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0248_));
 sky130_fd_sc_hd__or2_1 _3298_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .B(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _3299_ (.A0(net94),
    .A1(net1219),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0250_));
 sky130_fd_sc_hd__o211a_1 _3300_ (.A1(_0084_),
    .A2(_0250_),
    .B1(_0249_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0251_));
 sky130_fd_sc_hd__o32a_2 _3301_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0247_),
    .A3(_0251_),
    .B1(_0160_),
    .B2(_0162_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _3302_ (.A0(net200),
    .A1(net80),
    .A2(net23),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0252_));
 sky130_fd_sc_hd__mux4_2 _3303_ (.A0(net192),
    .A1(net68),
    .A2(net12),
    .A3(net115),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _3304_ (.A0(_0253_),
    .A1(_0252_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0254_));
 sky130_fd_sc_hd__mux4_1 _3305_ (.A0(net973),
    .A1(net968),
    .A2(net988),
    .A3(net992),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0255_));
 sky130_fd_sc_hd__or2_1 _3306_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .B(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__mux4_1 _3307_ (.A0(net979),
    .A1(net1019),
    .A2(net984),
    .A3(net1002),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0257_));
 sky130_fd_sc_hd__o211a_1 _3308_ (.A1(_0075_),
    .A2(_0257_),
    .B1(_0256_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0258_));
 sky130_fd_sc_hd__or2_1 _3309_ (.A(net205),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_0259_));
 sky130_fd_sc_hd__o21ai_1 _3310_ (.A1(net1256),
    .A2(_0052_),
    .B1(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__mux4_1 _3311_ (.A0(net1011),
    .A1(net1046),
    .A2(net1026),
    .A3(net1050),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3312_ (.A0(net1036),
    .A1(net1006),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0262_));
 sky130_fd_sc_hd__nand2b_1 _3313_ (.A_N(net1021),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .Y(_0263_));
 sky130_fd_sc_hd__o21a_1 _3314_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(net1031),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0264_));
 sky130_fd_sc_hd__a221o_1 _3315_ (.A1(_0053_),
    .A2(_0262_),
    .B1(_0263_),
    .B2(_0264_),
    .C1(_0054_),
    .X(_0265_));
 sky130_fd_sc_hd__o211a_1 _3316_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0261_),
    .B1(_0265_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0266_));
 sky130_fd_sc_hd__a211o_4 _3317_ (.A1(net664),
    .A2(_0218_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .C1(_0242_),
    .X(_0267_));
 sky130_fd_sc_hd__nand2b_1 _3318_ (.A_N(net190),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .Y(_0268_));
 sky130_fd_sc_hd__mux2_1 _3319_ (.A0(net2),
    .A1(net10),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0269_));
 sky130_fd_sc_hd__a21o_1 _3320_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0269_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0270_));
 sky130_fd_sc_hd__a31o_4 _3321_ (.A1(_0267_),
    .A2(_0053_),
    .A3(_0268_),
    .B1(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__mux4_1 _3322_ (.A0(net58),
    .A1(net66),
    .A2(net60),
    .A3(net94),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0272_));
 sky130_fd_sc_hd__o21ba_1 _3323_ (.A1(_0054_),
    .A2(_0272_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0273_));
 sky130_fd_sc_hd__a21o_1 _3324_ (.A1(_0271_),
    .A2(_0273_),
    .B1(_0266_),
    .X(_0274_));
 sky130_fd_sc_hd__a211oi_4 _3325_ (.A1(_0273_),
    .A2(_0271_),
    .B1(_0052_),
    .C1(_0266_),
    .Y(_0275_));
 sky130_fd_sc_hd__o21ai_1 _3326_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(net97),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_0276_));
 sky130_fd_sc_hd__o22a_1 _3327_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0260_),
    .B1(_0275_),
    .B2(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__clkinv_2 _3328_ (.A(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__o221a_4 _3329_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0260_),
    .B1(_0276_),
    .B2(_0275_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .X(_0279_));
 sky130_fd_sc_hd__mux4_2 _3330_ (.A0(net708),
    .A1(net750),
    .A2(net723),
    .A3(net1041),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0280_));
 sky130_fd_sc_hd__and2_4 _3331_ (.A(_0280_),
    .B(_0058_),
    .X(_0281_));
 sky130_fd_sc_hd__mux4_2 _3332_ (.A0(net737),
    .A1(net1005),
    .A2(net1030),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0282_));
 sky130_fd_sc_hd__a21bo_1 _3333_ (.A1(_0282_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_4 _3334_ (.A0(net744),
    .A1(net187),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _3335_ (.A0(net199),
    .A1(net7),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0285_));
 sky130_fd_sc_hd__or2_1 _3336_ (.A(_0057_),
    .B(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__o211a_1 _3337_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .A2(_0284_),
    .B1(_0286_),
    .C1(_0058_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _3338_ (.A0(net1256),
    .A1(net63),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0288_));
 sky130_fd_sc_hd__or2_1 _3339_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .B(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _3340_ (.A0(net99),
    .A1(net118),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0290_));
 sky130_fd_sc_hd__o211a_1 _3341_ (.A1(_0057_),
    .A2(_0290_),
    .B1(_0289_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_0291_));
 sky130_fd_sc_hd__o32a_4 _3342_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ),
    .A2(_0287_),
    .A3(_0291_),
    .B1(_0283_),
    .B2(_0281_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__o21ai_4 _3343_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ),
    .Y(_0292_));
 sky130_fd_sc_hd__mux4_1 _3344_ (.A0(net971),
    .A1(net728),
    .A2(net985),
    .A3(net975),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0293_));
 sky130_fd_sc_hd__mux4_1 _3345_ (.A0(net980),
    .A1(net995),
    .A2(net1016),
    .A3(net1013),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_4 _3346_ (.A0(_0293_),
    .A1(_0294_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0295_));
 sky130_fd_sc_hd__mux4_1 _3347_ (.A0(net181),
    .A1(net1218),
    .A2(net193),
    .A3(net127),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .X(_0296_));
 sky130_fd_sc_hd__mux4_1 _3348_ (.A0(net1216),
    .A1(net73),
    .A2(net217),
    .A3(net229),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _3349_ (.A0(_0296_),
    .A1(_0297_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_8 _3350_ (.A0(_0298_),
    .A1(_0295_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ));
 sky130_fd_sc_hd__mux4_1 _3351_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net16),
    .A2(net72),
    .A3(net108),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ),
    .X(_0299_));
 sky130_fd_sc_hd__o21ba_4 _3352_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .A2(net1004),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ),
    .X(_0300_));
 sky130_fd_sc_hd__o21ai_4 _3353_ (.A1(_0056_),
    .A2(net965),
    .B1(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__o21ai_4 _3354_ (.A1(_0292_),
    .A2(_0279_),
    .B1(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__o211ai_2 _3355_ (.A1(_0279_),
    .A2(_0292_),
    .B1(_0055_),
    .C1(_0301_),
    .Y(_0303_));
 sky130_fd_sc_hd__a21oi_1 _3356_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(_0059_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .Y(_0304_));
 sky130_fd_sc_hd__mux2_1 _3357_ (.A0(net209),
    .A1(net1068),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0305_));
 sky130_fd_sc_hd__a21bo_1 _3358_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .A2(_0305_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0306_));
 sky130_fd_sc_hd__a21o_1 _3359_ (.A1(_0304_),
    .A2(_0303_),
    .B1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__mux4_1 _3360_ (.A0(net175),
    .A1(net1218),
    .A2(net183),
    .A3(net129),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0308_));
 sky130_fd_sc_hd__o21ba_1 _3361_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_0308_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0309_));
 sky130_fd_sc_hd__o21ba_1 _3362_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(net978),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0310_));
 sky130_fd_sc_hd__o21a_1 _3363_ (.A1(_0055_),
    .A2(net997),
    .B1(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _3364_ (.A0(net1019),
    .A1(net1014),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0312_));
 sky130_fd_sc_hd__a21bo_1 _3365_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .A2(_0312_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0313_));
 sky130_fd_sc_hd__or2_1 _3366_ (.A(_0055_),
    .B(net968),
    .X(_0314_));
 sky130_fd_sc_hd__o21ba_1 _3367_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(net974),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(net988),
    .A1(net993),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0316_));
 sky130_fd_sc_hd__a221o_1 _3369_ (.A1(_0314_),
    .A2(_0315_),
    .B1(_0316_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0317_));
 sky130_fd_sc_hd__o211a_1 _3370_ (.A1(_0311_),
    .A2(_0313_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ),
    .C1(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__a21o_4 _3371_ (.A1(_0309_),
    .A2(net739),
    .B1(_0318_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ));
 sky130_fd_sc_hd__a211o_1 _3372_ (.A1(net712),
    .A2(_0309_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .C1(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__a21oi_1 _3373_ (.A1(_0060_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .Y(_0320_));
 sky130_fd_sc_hd__mux2_1 _3374_ (.A0(net74),
    .A1(net110),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .X(_0321_));
 sky130_fd_sc_hd__a22o_1 _3375_ (.A1(_0319_),
    .A2(_0320_),
    .B1(_0321_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0322_));
 sky130_fd_sc_hd__a221o_2 _3376_ (.A1(_0320_),
    .A2(_0319_),
    .B1(_0321_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .C1(_0074_),
    .X(_0323_));
 sky130_fd_sc_hd__o21ba_2 _3377_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .A2(net1030),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ),
    .X(_0324_));
 sky130_fd_sc_hd__a211oi_2 _3378_ (.A1(_0218_),
    .A2(_0217_),
    .B1(_0242_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .Y(_0325_));
 sky130_fd_sc_hd__and2_1 _3379_ (.A(_0042_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _3380_ (.A0(net200),
    .A1(net8),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0327_));
 sky130_fd_sc_hd__nand2_1 _3381_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__o311a_4 _3382_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0325_),
    .A3(_0326_),
    .B1(_0328_),
    .C1(_0043_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(net1255),
    .A1(net64),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0330_));
 sky130_fd_sc_hd__inv_1 _3384_ (.A(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__mux2_1 _3385_ (.A0(net100),
    .A1(net114),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_1 _3386_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .B(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__o211a_1 _3387_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0331_),
    .B1(_0333_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0334_));
 sky130_fd_sc_hd__mux4_1 _3388_ (.A0(net1034),
    .A1(net1004),
    .A2(net695),
    .A3(net676),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0335_));
 sky130_fd_sc_hd__mux4_2 _3389_ (.A0(net1009),
    .A1(net1045),
    .A2(net1049),
    .A3(net1039),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0336_));
 sky130_fd_sc_hd__o21a_1 _3390_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0336_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0337_));
 sky130_fd_sc_hd__o21ai_2 _3391_ (.A1(_0043_),
    .A2(_0335_),
    .B1(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__o31ai_2 _3392_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0329_),
    .A3(_0334_),
    .B1(_0338_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _3393_ (.A0(net708),
    .A1(net1024),
    .A2(net723),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0339_));
 sky130_fd_sc_hd__or2_4 _3394_ (.A(_0339_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0340_));
 sky130_fd_sc_hd__mux4_1 _3395_ (.A0(net1036),
    .A1(net1006),
    .A2(net1031),
    .A3(net1021),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0341_));
 sky130_fd_sc_hd__o21a_1 _3396_ (.A1(_0064_),
    .A2(_0341_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0342_));
 sky130_fd_sc_hd__mux4_1 _3397_ (.A0(net21),
    .A1(net99),
    .A2(net63),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0343_));
 sky130_fd_sc_hd__mux4_1 _3398_ (.A0(net187),
    .A1(net1),
    .A2(net199),
    .A3(net7),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _3399_ (.A0(_0343_),
    .A1(_0344_),
    .S(_0064_),
    .X(_0345_));
 sky130_fd_sc_hd__a22o_4 _3400_ (.A1(_0342_),
    .A2(_0340_),
    .B1(_0345_),
    .B2(_0065_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _3401_ (.A0(net208),
    .A1(net115),
    .A2(net80),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ),
    .X(_0346_));
 sky130_fd_sc_hd__or2_4 _3402_ (.A(_0346_),
    .B(_0074_),
    .X(_0347_));
 sky130_fd_sc_hd__o211a_4 _3403_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ),
    .B1(_0347_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ),
    .X(_0348_));
 sky130_fd_sc_hd__a21oi_4 _3404_ (.A1(_0324_),
    .A2(_0323_),
    .B1(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _3405_ (.A(net738),
    .Y(_0350_));
 sky130_fd_sc_hd__a211o_1 _3406_ (.A1(_0323_),
    .A2(_0324_),
    .B1(_0348_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0351_));
 sky130_fd_sc_hd__a21oi_1 _3407_ (.A1(_0045_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .Y(_0352_));
 sky130_fd_sc_hd__mux2_1 _3408_ (.A0(net210),
    .A1(net1067),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0353_));
 sky130_fd_sc_hd__a221o_1 _3409_ (.A1(_0351_),
    .A2(_0352_),
    .B1(_0353_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .C1(_0075_),
    .X(_0354_));
 sky130_fd_sc_hd__mux4_1 _3410_ (.A0(net176),
    .A1(net184),
    .A2(net1217),
    .A3(net130),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0355_));
 sky130_fd_sc_hd__o21ba_1 _3411_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_0355_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0356_));
 sky130_fd_sc_hd__a21o_2 _3412_ (.A1(_0354_),
    .A2(_0356_),
    .B1(_0258_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ));
 sky130_fd_sc_hd__or2_1 _3413_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .X(_0357_));
 sky130_fd_sc_hd__a21oi_1 _3414_ (.A1(_0083_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ),
    .Y(_0358_));
 sky130_fd_sc_hd__mux4_1 _3415_ (.A0(net1011),
    .A1(net1046),
    .A2(net1026),
    .A3(net1052),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _3416_ (.A(_0092_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__mux4_1 _3417_ (.A0(net1042),
    .A1(net1033),
    .A2(net1037),
    .A3(net1054),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0361_));
 sky130_fd_sc_hd__a21bo_1 _3418_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_0361_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0362_));
 sky130_fd_sc_hd__mux4_2 _3419_ (.A0(net981),
    .A1(net996),
    .A2(net1016),
    .A3(net1015),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0363_));
 sky130_fd_sc_hd__and2_4 _3420_ (.A(_0363_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0364_));
 sky130_fd_sc_hd__mux4_2 _3421_ (.A0(net972),
    .A1(net985),
    .A2(net991),
    .A3(net976),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0365_));
 sky130_fd_sc_hd__a21bo_1 _3422_ (.A1(_0022_),
    .A2(_0365_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0366_));
 sky130_fd_sc_hd__mux4_1 _3423_ (.A0(net179),
    .A1(net195),
    .A2(net119),
    .A3(net125),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _3424_ (.A(_0022_),
    .B(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _3425_ (.A0(net1216),
    .A1(net71),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(net215),
    .A1(net229),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0370_));
 sky130_fd_sc_hd__nand2b_1 _3427_ (.A_N(_0370_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .Y(_0371_));
 sky130_fd_sc_hd__o211a_1 _3428_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .A2(_0369_),
    .B1(_0371_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0372_));
 sky130_fd_sc_hd__o32a_4 _3429_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .A2(_0368_),
    .A3(_0372_),
    .B1(_0364_),
    .B2(_0366_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ));
 sky130_fd_sc_hd__mux4_2 _3430_ (.A0(net204),
    .A1(net231),
    .A2(net84),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .X(_0373_));
 sky130_fd_sc_hd__mux4_1 _3431_ (.A0(net971),
    .A1(net728),
    .A2(net991),
    .A3(net975),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0374_));
 sky130_fd_sc_hd__mux4_1 _3432_ (.A0(net980),
    .A1(net995),
    .A2(net1016),
    .A3(net1013),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_4 _3433_ (.A0(_0374_),
    .A1(_0375_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0376_));
 sky130_fd_sc_hd__mux4_1 _3434_ (.A0(net174),
    .A1(net180),
    .A2(net126),
    .A3(net1215),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0377_));
 sky130_fd_sc_hd__mux4_1 _3435_ (.A0(net72),
    .A1(net216),
    .A2(net84),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(_0377_),
    .A1(_0378_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0379_));
 sky130_fd_sc_hd__or2_1 _3437_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .B(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__o21ai_4 _3438_ (.A1(_0376_),
    .A2(_0046_),
    .B1(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_4 _3439_ (.A(_0381_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _3440_ (.A0(net190),
    .A1(net136),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A3(net226),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0382_));
 sky130_fd_sc_hd__mux4_2 _3441_ (.A0(net980),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .A2(_0382_),
    .A3(net688),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_4 _3442_ (.A0(net618),
    .A1(net192),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _3443_ (.A0(net1257),
    .A1(net12),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _3444_ (.A(_0091_),
    .B(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__o211a_1 _3445_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0384_),
    .B1(_0386_),
    .C1(_0092_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(net60),
    .A1(net68),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _3447_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .B(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(net94),
    .A1(net1219),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0390_));
 sky130_fd_sc_hd__o211a_1 _3449_ (.A1(_0091_),
    .A2(_0390_),
    .B1(_0389_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0391_));
 sky130_fd_sc_hd__o32a_4 _3450_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0391_),
    .A3(_0387_),
    .B1(_0360_),
    .B2(_0362_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(net75),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0392_));
 sky130_fd_sc_hd__a221o_1 _3452_ (.A1(_0357_),
    .A2(_0358_),
    .B1(_0392_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0393_));
 sky130_fd_sc_hd__o311a_4 _3453_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0329_),
    .A3(_0334_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .C1(_0338_),
    .X(_0394_));
 sky130_fd_sc_hd__o21ai_2 _3454_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .A2(net104),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2b_1 _3455_ (.A_N(net7),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .Y(_0396_));
 sky130_fd_sc_hd__o21ai_2 _3456_ (.A1(net199),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .B1(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__o22ai_4 _3457_ (.A1(_0395_),
    .A2(net627),
    .B1(_0397_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .Y(_0398_));
 sky130_fd_sc_hd__o221a_4 _3458_ (.A1(_0394_),
    .A2(_0395_),
    .B1(_0397_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .X(_0399_));
 sky130_fd_sc_hd__mux4_2 _3459_ (.A0(net1010),
    .A1(net724),
    .A2(net1024),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0400_));
 sky130_fd_sc_hd__mux4_1 _3460_ (.A0(net1034),
    .A1(net1005),
    .A2(net1029),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_4 _3461_ (.A0(_0400_),
    .A1(_0401_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_0402_));
 sky130_fd_sc_hd__mux4_2 _3462_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .A1(net197),
    .A2(net189),
    .A3(net9),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .X(_0403_));
 sky130_fd_sc_hd__mux4_1 _3463_ (.A0(net1256),
    .A1(net65),
    .A2(net101),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_4 _3464_ (.A0(_0403_),
    .A1(_0404_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_4 _3465_ (.A0(_0405_),
    .A1(_0402_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__o21ai_4 _3466_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .Y(_0406_));
 sky130_fd_sc_hd__mux4_2 _3467_ (.A0(net689),
    .A1(net70),
    .A2(net14),
    .A3(net106),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3468_ (.A0(net1039),
    .A1(_0407_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .X(_0408_));
 sky130_fd_sc_hd__nand2b_1 _3469_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__o21ai_4 _3470_ (.A1(_0399_),
    .A2(_0406_),
    .B1(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__o211a_1 _3471_ (.A1(_0399_),
    .A2(_0406_),
    .B1(_0409_),
    .C1(_0020_),
    .X(_0411_));
 sky130_fd_sc_hd__nor2_1 _3472_ (.A(_0020_),
    .B(net69),
    .Y(_0412_));
 sky130_fd_sc_hd__mux2_1 _3473_ (.A0(net209),
    .A1(net1068),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_0413_));
 sky130_fd_sc_hd__nand2_1 _3474_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__o311ai_4 _3475_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0412_),
    .A3(_0411_),
    .B1(_0414_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .Y(_0415_));
 sky130_fd_sc_hd__mux4_1 _3476_ (.A0(net173),
    .A1(net177),
    .A2(net119),
    .A3(net141),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0416_));
 sky130_fd_sc_hd__o21ba_1 _3477_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0416_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(net978),
    .A1(net983),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_0418_));
 sky130_fd_sc_hd__inv_2 _3479_ (.A(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(net997),
    .A1(net1014),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_0420_));
 sky130_fd_sc_hd__o21ai_1 _3481_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0419_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .Y(_0421_));
 sky130_fd_sc_hd__a21o_1 _3482_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0420_),
    .B1(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__mux4_1 _3483_ (.A0(net973),
    .A1(net968),
    .A2(net987),
    .A3(net992),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0423_));
 sky130_fd_sc_hd__o211a_1 _3484_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0423_),
    .B1(_0422_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0424_));
 sky130_fd_sc_hd__a21oi_2 _3485_ (.A1(_0415_),
    .A2(_0417_),
    .B1(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_1 _3486_ (.A(_0425_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ));
 sky130_fd_sc_hd__mux2_1 _3487_ (.A0(_0425_),
    .A1(_0044_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(net76),
    .A1(net112),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _3489_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__o211a_1 _3490_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ),
    .A2(_0426_),
    .B1(_0428_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0429_));
 sky130_fd_sc_hd__nor2_1 _3491_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__a22o_1 _3492_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ),
    .A2(_0254_),
    .B1(_0393_),
    .B2(_0430_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ),
    .S(net1064),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ),
    .A1(_0431_),
    .S(net1058),
    .X(_0432_));
 sky130_fd_sc_hd__mux4_1 _3495_ (.A0(net1011),
    .A1(net1046),
    .A2(net1050),
    .A3(net1042),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0433_));
 sky130_fd_sc_hd__or2_1 _3496_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .B(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__mux4_1 _3497_ (.A0(net1036),
    .A1(net1006),
    .A2(net1031),
    .A3(net1054),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0435_));
 sky130_fd_sc_hd__o21a_1 _3498_ (.A1(_0070_),
    .A2(_0435_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0436_));
 sky130_fd_sc_hd__mux4_1 _3499_ (.A0(net1255),
    .A1(net64),
    .A2(net100),
    .A3(net116),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0437_));
 sky130_fd_sc_hd__mux4_1 _3500_ (.A0(net188),
    .A1(net200),
    .A2(net2),
    .A3(net8),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _3501_ (.A0(_0437_),
    .A1(_0438_),
    .S(_0070_),
    .X(_0439_));
 sky130_fd_sc_hd__a22o_1 _3502_ (.A1(_0434_),
    .A2(_0436_),
    .B1(_0439_),
    .B2(_0071_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _3503_ (.A0(net8),
    .A1(net117),
    .A2(net88),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_0440_));
 sky130_fd_sc_hd__mux4_1 _3504_ (.A0(net208),
    .A1(net67),
    .A2(net11),
    .A3(net103),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _3505_ (.A0(_0441_),
    .A1(_0440_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _3506_ (.A0(_0425_),
    .A1(_0044_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(net76),
    .A1(net112),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0444_));
 sky130_fd_sc_hd__nand2_1 _3508_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__o211a_1 _3509_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ),
    .A2(_0443_),
    .B1(_0445_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0446_));
 sky130_fd_sc_hd__mux4_1 _3510_ (.A0(net19),
    .A1(net111),
    .A2(net75),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_0447_));
 sky130_fd_sc_hd__o21ba_1 _3511_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(_0447_),
    .B1_N(_0446_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_2 _3512_ (.A0(_0448_),
    .A1(_0442_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ));
 sky130_fd_sc_hd__nand2b_1 _3513_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ),
    .B(net1062),
    .Y(_0449_));
 sky130_fd_sc_hd__o21ai_4 _3514_ (.A1(net1062),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ),
    .B1(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__mux4_2 _3515_ (.A0(net691),
    .A1(net707),
    .A2(net991),
    .A3(net975),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0451_));
 sky130_fd_sc_hd__mux4_2 _3516_ (.A0(net715),
    .A1(net995),
    .A2(net1016),
    .A3(net714),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_4 _3517_ (.A0(_0451_),
    .A1(_0452_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .X(_0453_));
 sky130_fd_sc_hd__mux4_1 _3518_ (.A0(net178),
    .A1(net194),
    .A2(net1217),
    .A3(net124),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0454_));
 sky130_fd_sc_hd__mux4_1 _3519_ (.A0(net1215),
    .A1(net214),
    .A2(net90),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _3520_ (.A0(_0454_),
    .A1(_0455_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_4 _3521_ (.A0(_0456_),
    .A1(_0453_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ));
 sky130_fd_sc_hd__mux2_1 _3522_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .A1(net13),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_0457_));
 sky130_fd_sc_hd__and2b_1 _3523_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ),
    .B(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__mux4_1 _3524_ (.A0(net1010),
    .A1(net724),
    .A2(net1025),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0459_));
 sky130_fd_sc_hd__nor2_1 _3525_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__mux4_2 _3526_ (.A0(net737),
    .A1(net1005),
    .A2(net1029),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0461_));
 sky130_fd_sc_hd__o21ai_2 _3527_ (.A1(_0461_),
    .A2(_0082_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ),
    .Y(_0462_));
 sky130_fd_sc_hd__mux4_1 _3528_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .A1(net9),
    .A2(net189),
    .A3(net1256),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0463_));
 sky130_fd_sc_hd__nor2_1 _3529_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__mux4_1 _3530_ (.A0(net65),
    .A1(net101),
    .A2(net77),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0465_));
 sky130_fd_sc_hd__nor2_1 _3531_ (.A(_0082_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__o32a_4 _3532_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ),
    .A2(_0464_),
    .A3(_0466_),
    .B1(_0460_),
    .B2(_0462_),
    .X(_0467_));
 sky130_fd_sc_hd__inv_4 _3533_ (.A(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _3534_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ),
    .B(_0467_),
    .Y(_0469_));
 sky130_fd_sc_hd__o211a_1 _3535_ (.A1(net69),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ),
    .C1(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _3536_ (.A0(net689),
    .A1(net14),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0471_));
 sky130_fd_sc_hd__and2b_1 _3537_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ),
    .B(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(net70),
    .A1(net106),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0473_));
 sky130_fd_sc_hd__a21bo_1 _3539_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_0473_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0474_));
 sky130_fd_sc_hd__o32a_1 _3540_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0458_),
    .A3(_0470_),
    .B1(_0472_),
    .B2(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__mux4_2 _3541_ (.A0(net1009),
    .A1(net1024),
    .A2(net723),
    .A3(net1039),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0476_));
 sky130_fd_sc_hd__or2_4 _3542_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .B(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__mux4_2 _3543_ (.A0(net737),
    .A1(net736),
    .A2(net1029),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0478_));
 sky130_fd_sc_hd__o211a_1 _3544_ (.A1(_0478_),
    .A2(_0050_),
    .B1(_0477_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0479_));
 sky130_fd_sc_hd__or2_1 _3545_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .B(_0199_),
    .X(_0480_));
 sky130_fd_sc_hd__a21oi_1 _3546_ (.A1(_0049_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0481_));
 sky130_fd_sc_hd__mux2_1 _3547_ (.A0(net7),
    .A1(net1256),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0482_));
 sky130_fd_sc_hd__a221o_1 _3548_ (.A1(_0481_),
    .A2(_0480_),
    .B1(_0482_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(net63),
    .A1(net79),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0484_));
 sky130_fd_sc_hd__and2b_1 _3550_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .B(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3551_ (.A0(net99),
    .A1(net113),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0486_));
 sky130_fd_sc_hd__a211o_1 _3552_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0486_),
    .B1(_0485_),
    .C1(_0050_),
    .X(_0487_));
 sky130_fd_sc_hd__a31o_1 _3553_ (.A1(_0051_),
    .A2(_0483_),
    .A3(_0487_),
    .B1(_0479_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _3554_ (.A0(net197),
    .A1(net1256),
    .A2(net77),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ),
    .X(_0488_));
 sky130_fd_sc_hd__mux4_2 _3555_ (.A0(net185),
    .A1(net5),
    .A2(net61),
    .A3(net118),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_4 _3556_ (.A0(_0489_),
    .A1(_0488_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_4 _3557_ (.A0(_0475_),
    .A1(_0490_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ));
 sky130_fd_sc_hd__nand2b_1 _3558_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ),
    .B(net1060),
    .Y(_0491_));
 sky130_fd_sc_hd__o21ai_4 _3559_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ),
    .A2(net1060),
    .B1(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__or2_1 _3560_ (.A(_0450_),
    .B(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__mux4_2 _3561_ (.A0(net1036),
    .A1(net1006),
    .A2(net1031),
    .A3(net1021),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0494_));
 sky130_fd_sc_hd__mux4_2 _3562_ (.A0(net1009),
    .A1(net1045),
    .A2(net750),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0495_));
 sky130_fd_sc_hd__and2b_1 _3563_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__a21bo_1 _3564_ (.A1(_0494_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(net101),
    .A1(net117),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0498_));
 sky130_fd_sc_hd__nand2b_1 _3566_ (.A_N(_0498_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .Y(_0499_));
 sky130_fd_sc_hd__mux2_1 _3567_ (.A0(net65),
    .A1(net77),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0500_));
 sky130_fd_sc_hd__o211a_1 _3568_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_0500_),
    .B1(_0499_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0501_));
 sky130_fd_sc_hd__mux4_1 _3569_ (.A0(net189),
    .A1(net9),
    .A2(net1258),
    .A3(net1256),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0502_));
 sky130_fd_sc_hd__and2b_1 _3570_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__o32a_4 _3571_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0501_),
    .A3(_0503_),
    .B1(_0496_),
    .B2(_0497_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _3572_ (.A0(net974),
    .A1(net970),
    .A2(net989),
    .A3(net994),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0504_));
 sky130_fd_sc_hd__or2_1 _3573_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .B(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__mux4_1 _3574_ (.A0(net984),
    .A1(net998),
    .A2(net1020),
    .A3(net1001),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0506_));
 sky130_fd_sc_hd__o211a_1 _3575_ (.A1(_0079_),
    .A2(_0506_),
    .B1(_0505_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0507_));
 sky130_fd_sc_hd__mux4_2 _3576_ (.A0(net1045),
    .A1(net750),
    .A2(net713),
    .A3(net1039),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0508_));
 sky130_fd_sc_hd__or2_4 _3577_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ),
    .B(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__mux4_2 _3578_ (.A0(net1034),
    .A1(net736),
    .A2(net1029),
    .A3(net676),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0510_));
 sky130_fd_sc_hd__o211a_1 _3579_ (.A1(_0077_),
    .A2(_0510_),
    .B1(_0509_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0511_));
 sky130_fd_sc_hd__or2_4 _3580_ (.A(_0383_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0512_));
 sky130_fd_sc_hd__a21oi_1 _3581_ (.A1(_0024_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .Y(_0513_));
 sky130_fd_sc_hd__mux2_1 _3582_ (.A0(net198),
    .A1(net24),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0514_));
 sky130_fd_sc_hd__a221o_1 _3583_ (.A1(_0513_),
    .A2(_0512_),
    .B1(_0514_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(net1255),
    .A1(net62),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0516_));
 sky130_fd_sc_hd__and2b_1 _3585_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .B(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _3586_ (.A0(net98),
    .A1(net114),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0518_));
 sky130_fd_sc_hd__a211o_1 _3587_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_0518_),
    .B1(_0517_),
    .C1(_0077_),
    .X(_0519_));
 sky130_fd_sc_hd__a31o_4 _3588_ (.A1(_0515_),
    .A2(_0078_),
    .A3(_0519_),
    .B1(_0511_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__mux4_2 _3589_ (.A0(net198),
    .A1(net86),
    .A2(net101),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0520_));
 sky130_fd_sc_hd__or2_4 _3590_ (.A(_0076_),
    .B(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__o211a_4 _3591_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .B1(_0521_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ),
    .X(_0522_));
 sky130_fd_sc_hd__a211o_1 _3592_ (.A1(_0417_),
    .A2(_0415_),
    .B1(_0424_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0523_));
 sky130_fd_sc_hd__a21oi_1 _3593_ (.A1(_0044_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .Y(_0524_));
 sky130_fd_sc_hd__mux2_1 _3594_ (.A0(net76),
    .A1(net112),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0525_));
 sky130_fd_sc_hd__a22o_4 _3595_ (.A1(_0524_),
    .A2(_0523_),
    .B1(_0525_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_0526_));
 sky130_fd_sc_hd__a221o_1 _3596_ (.A1(_0524_),
    .A2(_0523_),
    .B1(_0525_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .C1(_0076_),
    .X(_0527_));
 sky130_fd_sc_hd__o21ba_1 _3597_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .A2(net1035),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ),
    .X(_0528_));
 sky130_fd_sc_hd__a21o_4 _3598_ (.A1(_0527_),
    .A2(_0528_),
    .B1(_0522_),
    .X(_0529_));
 sky130_fd_sc_hd__a211o_1 _3599_ (.A1(_0528_),
    .A2(_0527_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .C1(_0522_),
    .X(_0530_));
 sky130_fd_sc_hd__a21oi_1 _3600_ (.A1(_0061_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .Y(_0531_));
 sky130_fd_sc_hd__mux2_1 _3601_ (.A0(net210),
    .A1(net1067),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0532_));
 sky130_fd_sc_hd__a221o_1 _3602_ (.A1(_0531_),
    .A2(_0530_),
    .B1(_0532_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .C1(_0079_),
    .X(_0533_));
 sky130_fd_sc_hd__mux4_1 _3603_ (.A0(net174),
    .A1(net182),
    .A2(net120),
    .A3(net128),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0534_));
 sky130_fd_sc_hd__o21ba_1 _3604_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0534_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0535_));
 sky130_fd_sc_hd__a21o_4 _3605_ (.A1(_0535_),
    .A2(_0533_),
    .B1(_0507_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ));
 sky130_fd_sc_hd__inv_1 _3606_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .Y(_0536_));
 sky130_fd_sc_hd__mux4_2 _3607_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .A1(net109),
    .A2(net17),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_4 _3608_ (.A0(_0537_),
    .A1(_0322_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .X(_0538_));
 sky130_fd_sc_hd__mux4_1 _3609_ (.A0(net198),
    .A1(net114),
    .A2(net1255),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_0539_));
 sky130_fd_sc_hd__mux4_2 _3610_ (.A0(net189),
    .A1(net65),
    .A2(net23),
    .A3(net101),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _3611_ (.A0(_0540_),
    .A1(_0539_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_4 _3612_ (.A0(_0538_),
    .A1(_0541_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ));
 sky130_fd_sc_hd__nand2b_1 _3613_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ),
    .B(net1060),
    .Y(_0542_));
 sky130_fd_sc_hd__o21ai_4 _3614_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ),
    .A2(net1060),
    .B1(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__a211o_1 _3615_ (.A1(_0527_),
    .A2(_0528_),
    .B1(_0522_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0544_));
 sky130_fd_sc_hd__a211o_1 _3616_ (.A1(_0323_),
    .A2(_0324_),
    .B1(_0348_),
    .C1(_0107_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(net74),
    .A1(net210),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0546_));
 sky130_fd_sc_hd__a21bo_1 _3618_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0546_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0547_));
 sky130_fd_sc_hd__a31o_4 _3619_ (.A1(_0544_),
    .A2(_0108_),
    .A3(_0545_),
    .B1(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__mux4_1 _3620_ (.A0(net174),
    .A1(net182),
    .A2(net120),
    .A3(net128),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0549_));
 sky130_fd_sc_hd__o21ba_1 _3621_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0549_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0550_));
 sky130_fd_sc_hd__or2_1 _3622_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .B(net984),
    .X(_0551_));
 sky130_fd_sc_hd__o211a_1 _3623_ (.A1(_0107_),
    .A2(net998),
    .B1(_0551_),
    .C1(_0108_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_2 _3624_ (.A0(net734),
    .A1(net1015),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0553_));
 sky130_fd_sc_hd__a21bo_1 _3625_ (.A1(_0553_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0554_));
 sky130_fd_sc_hd__mux4_1 _3626_ (.A0(net974),
    .A1(net970),
    .A2(net989),
    .A3(net992),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0555_));
 sky130_fd_sc_hd__o221a_4 _3627_ (.A1(_0554_),
    .A2(_0552_),
    .B1(_0555_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0556_));
 sky130_fd_sc_hd__a21oi_4 _3628_ (.A1(_0548_),
    .A2(_0550_),
    .B1(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__a211o_1 _3629_ (.A1(_0548_),
    .A2(_0550_),
    .B1(_0106_),
    .C1(_0556_),
    .X(_0558_));
 sky130_fd_sc_hd__o21a_1 _3630_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .A2(net221),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .X(_0559_));
 sky130_fd_sc_hd__mux4_2 _3631_ (.A0(net724),
    .A1(net750),
    .A2(net1049),
    .A3(net1039),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0560_));
 sky130_fd_sc_hd__or2_4 _3632_ (.A(_0560_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0561_));
 sky130_fd_sc_hd__mux4_1 _3633_ (.A0(net1035),
    .A1(net736),
    .A2(net695),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0562_));
 sky130_fd_sc_hd__o21a_1 _3634_ (.A1(_0072_),
    .A2(_0562_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0563_));
 sky130_fd_sc_hd__mux4_1 _3635_ (.A0(net62),
    .A1(net78),
    .A2(net98),
    .A3(net114),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0564_));
 sky130_fd_sc_hd__mux4_1 _3636_ (.A0(net206),
    .A1(net1257),
    .A2(net6),
    .A3(net1255),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _3637_ (.A0(_0564_),
    .A1(_0565_),
    .S(_0072_),
    .X(_0566_));
 sky130_fd_sc_hd__a22o_4 _3638_ (.A1(_0561_),
    .A2(_0563_),
    .B1(_0566_),
    .B2(_0073_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ));
 sky130_fd_sc_hd__mux2_1 _3639_ (.A0(net185),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0567_));
 sky130_fd_sc_hd__a221o_1 _3640_ (.A1(_0559_),
    .A2(_0558_),
    .B1(_0567_),
    .B2(_0109_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0568_));
 sky130_fd_sc_hd__o21ba_1 _3641_ (.A1(_0110_),
    .A2(_0196_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0569_));
 sky130_fd_sc_hd__mux4_2 _3642_ (.A0(net193),
    .A1(net89),
    .A2(net229),
    .A3(net706),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .X(_0570_));
 sky130_fd_sc_hd__mux4_2 _3643_ (.A0(net177),
    .A1(net69),
    .A2(net142),
    .A3(net213),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0571_));
 sky130_fd_sc_hd__or2_1 _3644_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .B(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__o211a_1 _3645_ (.A1(_0110_),
    .A2(_0570_),
    .B1(_0572_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0573_));
 sky130_fd_sc_hd__a21o_1 _3646_ (.A1(_0568_),
    .A2(_0569_),
    .B1(_0573_),
    .X(\Tile_X0Y1_DSP_bot.B3 ));
 sky130_fd_sc_hd__a211o_4 _3647_ (.A1(_0569_),
    .A2(_0568_),
    .B1(_0573_),
    .C1(net1061),
    .X(_0574_));
 sky130_fd_sc_hd__nand2b_1 _3648_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ),
    .B(net1062),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _3649_ (.A(_0574_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__nor2_1 _3650_ (.A(_0543_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__nor2_1 _3651_ (.A(_0450_),
    .B(_0543_),
    .Y(_0578_));
 sky130_fd_sc_hd__nor2_1 _3652_ (.A(_0492_),
    .B(_0576_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2_1 _3653_ (.A(_0578_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2_1 _3654_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .B(_0183_),
    .Y(_0581_));
 sky130_fd_sc_hd__o211a_1 _3655_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .B1(_0581_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _3656_ (.A0(net185),
    .A1(net131),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_0583_));
 sky130_fd_sc_hd__and2b_1 _3657_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .B(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _3658_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A1(net222),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _3659_ (.A0(net186),
    .A1(net132),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0586_));
 sky130_fd_sc_hd__and2b_1 _3660_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .B(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__a21bo_1 _3661_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_0585_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0588_));
 sky130_fd_sc_hd__o32a_1 _3662_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0582_),
    .A3(_0584_),
    .B1(_0587_),
    .B2(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__mux4_2 _3663_ (.A0(net972),
    .A1(net986),
    .A2(net990),
    .A3(net976),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0590_));
 sky130_fd_sc_hd__mux4_2 _3664_ (.A0(net982),
    .A1(net996),
    .A2(net1018),
    .A3(net1001),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0591_));
 sky130_fd_sc_hd__or2_4 _3665_ (.A(_0591_),
    .B(_0100_),
    .X(_0592_));
 sky130_fd_sc_hd__o21a_1 _3666_ (.A1(_0590_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0593_));
 sky130_fd_sc_hd__mux4_1 _3667_ (.A0(net173),
    .A1(net179),
    .A2(net125),
    .A3(net1216),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0594_));
 sky130_fd_sc_hd__mux4_1 _3668_ (.A0(net71),
    .A1(net215),
    .A2(net83),
    .A3(net229),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _3669_ (.A0(_0594_),
    .A1(_0595_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0596_));
 sky130_fd_sc_hd__a22o_4 _3670_ (.A1(_0593_),
    .A2(_0592_),
    .B1(_0596_),
    .B2(_0101_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _3671_ (.A0(net193),
    .A1(net81),
    .A2(net1216),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0597_));
 sky130_fd_sc_hd__mux4_1 _3672_ (.A0(net177),
    .A1(net69),
    .A2(net123),
    .A3(net234),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _3673_ (.A0(_0598_),
    .A1(_0597_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_2 _3674_ (.A0(_0589_),
    .A1(_0599_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .X(\Tile_X0Y1_DSP_bot.A3 ));
 sky130_fd_sc_hd__nand2b_1 _3675_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ),
    .B(net1059),
    .Y(_0600_));
 sky130_fd_sc_hd__o21ai_4 _3676_ (.A1(net1059),
    .A2(\Tile_X0Y1_DSP_bot.A3 ),
    .B1(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__mux4_2 _3677_ (.A0(net708),
    .A1(net1045),
    .A2(net723),
    .A3(net1039),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0602_));
 sky130_fd_sc_hd__or2_4 _3678_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .B(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__mux4_1 _3679_ (.A0(net737),
    .A1(net736),
    .A2(net1030),
    .A3(net1023),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0604_));
 sky130_fd_sc_hd__o211a_1 _3680_ (.A1(_0062_),
    .A2(_0604_),
    .B1(_0603_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0605_));
 sky130_fd_sc_hd__or2_1 _3681_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .B(_0243_),
    .X(_0606_));
 sky130_fd_sc_hd__a21oi_1 _3682_ (.A1(_0042_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .Y(_0607_));
 sky130_fd_sc_hd__mux2_1 _3683_ (.A0(net8),
    .A1(net1255),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0608_));
 sky130_fd_sc_hd__a221o_1 _3684_ (.A1(_0606_),
    .A2(_0607_),
    .B1(_0608_),
    .B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _3685_ (.A0(net64),
    .A1(net80),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0610_));
 sky130_fd_sc_hd__and2b_1 _3686_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .B(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _3687_ (.A0(net100),
    .A1(net114),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0612_));
 sky130_fd_sc_hd__a211o_1 _3688_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0612_),
    .B1(_0611_),
    .C1(_0062_),
    .X(_0613_));
 sky130_fd_sc_hd__a31o_1 _3689_ (.A1(_0063_),
    .A2(_0609_),
    .A3(_0613_),
    .B1(_0605_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _3690_ (.A0(net197),
    .A1(net113),
    .A2(net85),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0614_));
 sky130_fd_sc_hd__mux4_1 _3691_ (.A0(net185),
    .A1(net61),
    .A2(net24),
    .A3(net97),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_4 _3692_ (.A0(_0615_),
    .A1(_0614_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0616_));
 sky130_fd_sc_hd__mux4_1 _3693_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .A1(net105),
    .A2(net69),
    .A3(_0274_),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _3694_ (.A0(_0617_),
    .A1(_0407_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_4 _3695_ (.A0(_0618_),
    .A1(_0616_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ));
 sky130_fd_sc_hd__nand2b_1 _3696_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ),
    .B(net1062),
    .Y(_0619_));
 sky130_fd_sc_hd__o21ai_4 _3697_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ),
    .A2(net1062),
    .B1(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__nor2_4 _3698_ (.A(_0601_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__mux4_1 _3699_ (.A0(net1010),
    .A1(net724),
    .A2(net1053),
    .A3(net1041),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0622_));
 sky130_fd_sc_hd__and2b_1 _3700_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .B(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__mux4_2 _3701_ (.A0(net1035),
    .A1(net1005),
    .A2(net1030),
    .A3(net1056),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0624_));
 sky130_fd_sc_hd__a21bo_1 _3702_ (.A1(_0624_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0625_));
 sky130_fd_sc_hd__mux4_1 _3703_ (.A0(net64),
    .A1(net100),
    .A2(net80),
    .A3(net114),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _3704_ (.A0(net8),
    .A1(net1255),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0627_));
 sky130_fd_sc_hd__nand2b_1 _3705_ (.A_N(_0627_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .Y(_0628_));
 sky130_fd_sc_hd__mux2_1 _3706_ (.A0(net208),
    .A1(net2),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0629_));
 sky130_fd_sc_hd__o21ba_1 _3707_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_0629_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .X(_0630_));
 sky130_fd_sc_hd__a221o_1 _3708_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .A2(_0626_),
    .B1(_0628_),
    .B2(_0630_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0631_));
 sky130_fd_sc_hd__o21ai_4 _3709_ (.A1(_0625_),
    .A2(_0623_),
    .B1(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__clkinv_2 _3710_ (.A(_0632_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _3711_ (.A0(net206),
    .A1(net24),
    .A2(net78),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ),
    .X(_0633_));
 sky130_fd_sc_hd__mux4_2 _3712_ (.A0(net189),
    .A1(net9),
    .A2(net87),
    .A3(net101),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _3713_ (.A0(_0634_),
    .A1(_0633_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0635_));
 sky130_fd_sc_hd__and2_1 _3714_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ),
    .B(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__mux4_1 _3715_ (.A0(net1011),
    .A1(net1046),
    .A2(net1027),
    .A3(net1051),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0637_));
 sky130_fd_sc_hd__and2_1 _3716_ (.A(_0088_),
    .B(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__mux4_1 _3717_ (.A0(net1036),
    .A1(net1008),
    .A2(net1032),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0639_));
 sky130_fd_sc_hd__a21bo_1 _3718_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0639_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_2 _3719_ (.A0(_0243_),
    .A1(net190),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _3720_ (.A0(net2),
    .A1(net10),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0642_));
 sky130_fd_sc_hd__or2_1 _3721_ (.A(_0087_),
    .B(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__o211a_1 _3722_ (.A1(_0641_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .B1(_0643_),
    .C1(_0088_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _3723_ (.A0(net58),
    .A1(net66),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0645_));
 sky130_fd_sc_hd__or2_1 _3724_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _3725_ (.A0(net94),
    .A1(net1219),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0647_));
 sky130_fd_sc_hd__o211a_1 _3726_ (.A1(_0087_),
    .A2(_0647_),
    .B1(_0646_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0648_));
 sky130_fd_sc_hd__o32a_4 _3727_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_0648_),
    .A3(_0644_),
    .B1(_0638_),
    .B2(_0640_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__mux2_1 _3728_ (.A0(net73),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0649_));
 sky130_fd_sc_hd__a211o_1 _3729_ (.A1(_0533_),
    .A2(_0535_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .C1(_0507_),
    .X(_0650_));
 sky130_fd_sc_hd__a21oi_1 _3730_ (.A1(_0080_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ),
    .Y(_0651_));
 sky130_fd_sc_hd__a22o_2 _3731_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ),
    .A2(_0649_),
    .B1(_0650_),
    .B2(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__a221o_1 _3732_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ),
    .A2(_0649_),
    .B1(_0650_),
    .B2(_0651_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0653_));
 sky130_fd_sc_hd__nor2_2 _3733_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ),
    .B(net710),
    .Y(_0654_));
 sky130_fd_sc_hd__a211o_1 _3734_ (.A1(_0060_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ),
    .C1(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _3735_ (.A0(net74),
    .A1(net110),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ),
    .X(_0656_));
 sky130_fd_sc_hd__nand2_1 _3736_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__a31oi_4 _3737_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_0657_),
    .A3(_0655_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_0658_));
 sky130_fd_sc_hd__a21o_1 _3738_ (.A1(_0653_),
    .A2(_0658_),
    .B1(_0636_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ));
 sky130_fd_sc_hd__a211o_4 _3739_ (.A1(_0653_),
    .A2(_0658_),
    .B1(net1061),
    .C1(_0636_),
    .X(_0659_));
 sky130_fd_sc_hd__nand2b_1 _3740_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ),
    .B(net1061),
    .Y(_0660_));
 sky130_fd_sc_hd__nand2_8 _3741_ (.A(_0659_),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__mux4_2 _3742_ (.A0(_0023_),
    .A1(_0102_),
    .A2(_0103_),
    .A3(_0229_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .X(_0662_));
 sky130_fd_sc_hd__nand2_1 _3743_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .B(_0382_),
    .Y(_0663_));
 sky130_fd_sc_hd__mux4_1 _3744_ (.A0(net692),
    .A1(net747),
    .A2(net733),
    .A3(net1013),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0664_));
 sky130_fd_sc_hd__mux4_2 _3745_ (.A0(net971),
    .A1(net985),
    .A2(net716),
    .A3(net976),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0665_));
 sky130_fd_sc_hd__or2_4 _3746_ (.A(_0665_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0666_));
 sky130_fd_sc_hd__o21a_1 _3747_ (.A1(_0104_),
    .A2(_0664_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0667_));
 sky130_fd_sc_hd__mux4_1 _3748_ (.A0(net203),
    .A1(net143),
    .A2(net119),
    .A3(net1216),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0668_));
 sky130_fd_sc_hd__mux4_1 _3749_ (.A0(net83),
    .A1(net91),
    .A2(net215),
    .A3(net229),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _3750_ (.A0(_0668_),
    .A1(_0669_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0670_));
 sky130_fd_sc_hd__a22o_4 _3751_ (.A1(_0667_),
    .A2(_0666_),
    .B1(_0670_),
    .B2(_0105_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _3752_ (.A0(net194),
    .A1(net230),
    .A2(net1215),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_0671_));
 sky130_fd_sc_hd__mux4_2 _3753_ (.A0(net181),
    .A1(net73),
    .A2(net141),
    .A3(net217),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_4 _3754_ (.A0(_0672_),
    .A1(_0671_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0673_));
 sky130_fd_sc_hd__o21ai_2 _3755_ (.A1(_0662_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .B1(_0663_),
    .Y(_0674_));
 sky130_fd_sc_hd__mux2_4 _3756_ (.A0(_0674_),
    .A1(_0673_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Tile_X0Y1_DSP_bot.A2 ));
 sky130_fd_sc_hd__nand2b_1 _3757_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ),
    .B(net1059),
    .Y(_0675_));
 sky130_fd_sc_hd__o21ai_4 _3758_ (.A1(\Tile_X0Y1_DSP_bot.A2 ),
    .A2(net1059),
    .B1(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__inv_2 _3759_ (.A(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__and3_1 _3760_ (.A(_0659_),
    .B(_0660_),
    .C(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__nor2_1 _3761_ (.A(_0601_),
    .B(_0661_),
    .Y(_0679_));
 sky130_fd_sc_hd__nor2_1 _3762_ (.A(_0620_),
    .B(_0676_),
    .Y(_0680_));
 sky130_fd_sc_hd__and2_4 _3763_ (.A(_0621_),
    .B(_0678_),
    .X(_0681_));
 sky130_fd_sc_hd__mux4_1 _3764_ (.A0(net1012),
    .A1(net1047),
    .A2(net1027),
    .A3(net1051),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0682_));
 sky130_fd_sc_hd__nand2b_1 _3765_ (.A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__mux4_2 _3766_ (.A0(net1038),
    .A1(net740),
    .A2(net1032),
    .A3(net1021),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0684_));
 sky130_fd_sc_hd__nand2_2 _3767_ (.A(_0684_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .Y(_0685_));
 sky130_fd_sc_hd__mux2_1 _3768_ (.A0(_0243_),
    .A1(net190),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0686_));
 sky130_fd_sc_hd__nor2_1 _3769_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__mux2_1 _3770_ (.A0(net2),
    .A1(net10),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0688_));
 sky130_fd_sc_hd__inv_1 _3771_ (.A(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__a211o_1 _3772_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .A2(_0689_),
    .B1(_0687_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _3773_ (.A0(net58),
    .A1(net60),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0691_));
 sky130_fd_sc_hd__or2_1 _3774_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .B(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _3775_ (.A0(net66),
    .A1(net94),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0693_));
 sky130_fd_sc_hd__o211a_1 _3776_ (.A1(_0086_),
    .A2(_0693_),
    .B1(_0692_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0694_));
 sky130_fd_sc_hd__nor2_1 _3777_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__a32o_2 _3778_ (.A1(_0685_),
    .A2(_0683_),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ),
    .B1(_0690_),
    .B2(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__inv_4 _3779_ (.A(_0696_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__mux4_2 _3780_ (.A0(net982),
    .A1(net747),
    .A2(net1018),
    .A3(net714),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0697_));
 sky130_fd_sc_hd__mux4_1 _3781_ (.A0(net972),
    .A1(net967),
    .A2(net990),
    .A3(net976),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_4 _3782_ (.A0(_0698_),
    .A1(_0697_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .X(_0699_));
 sky130_fd_sc_hd__mux4_1 _3783_ (.A0(net1215),
    .A1(net72),
    .A2(net216),
    .A3(net232),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0700_));
 sky130_fd_sc_hd__mux4_1 _3784_ (.A0(net180),
    .A1(net196),
    .A2(net120),
    .A3(net126),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _3785_ (.A0(_0701_),
    .A1(_0700_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_4 _3786_ (.A0(_0702_),
    .A1(_0699_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ));
 sky130_fd_sc_hd__mux4_2 _3787_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A1(net107),
    .A2(net15),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0703_));
 sky130_fd_sc_hd__mux4_2 _3788_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net16),
    .A2(net72),
    .A3(net108),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_4 _3789_ (.A0(_0703_),
    .A1(_0704_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0705_));
 sky130_fd_sc_hd__mux4_2 _3790_ (.A0(net187),
    .A1(net63),
    .A2(net7),
    .A3(net117),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_4 _3791_ (.A0(_0706_),
    .A1(_0398_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_4 _3792_ (.A0(_0705_),
    .A1(_0707_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ));
 sky130_fd_sc_hd__nand2b_1 _3793_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ),
    .B(net1061),
    .Y(_0708_));
 sky130_fd_sc_hd__o21ai_4 _3794_ (.A1(net1061),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .B1(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__mux4_2 _3795_ (.A0(net191),
    .A1(net11),
    .A2(net88),
    .A3(net103),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _3796_ (.A0(_0710_),
    .A1(_0346_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0711_));
 sky130_fd_sc_hd__a211o_1 _3797_ (.A1(_0354_),
    .A2(_0356_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .C1(_0258_),
    .X(_0712_));
 sky130_fd_sc_hd__a21oi_1 _3798_ (.A1(_0059_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ),
    .Y(_0713_));
 sky130_fd_sc_hd__mux4_2 _3799_ (.A0(net708),
    .A1(net724),
    .A2(net750),
    .A3(net1040),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0714_));
 sky130_fd_sc_hd__or2_4 _3800_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ),
    .B(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__mux4_2 _3801_ (.A0(net1035),
    .A1(net736),
    .A2(net695),
    .A3(net1023),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0716_));
 sky130_fd_sc_hd__o21a_1 _3802_ (.A1(_0716_),
    .A2(_0066_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0717_));
 sky130_fd_sc_hd__mux4_1 _3803_ (.A0(net189),
    .A1(net197),
    .A2(net1258),
    .A3(net9),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0718_));
 sky130_fd_sc_hd__mux4_1 _3804_ (.A0(net1256),
    .A1(net65),
    .A2(net101),
    .A3(net113),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _3805_ (.A0(_0718_),
    .A1(_0719_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0720_));
 sky130_fd_sc_hd__a22o_4 _3806_ (.A1(_0717_),
    .A2(_0715_),
    .B1(_0720_),
    .B2(_0067_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ));
 sky130_fd_sc_hd__mux2_1 _3807_ (.A0(net111),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .X(_0721_));
 sky130_fd_sc_hd__a221o_1 _3808_ (.A1(_0712_),
    .A2(_0713_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ),
    .B2(_0721_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _3809_ (.A0(_0425_),
    .A1(_0044_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _3810_ (.A0(net76),
    .A1(net112),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0724_));
 sky130_fd_sc_hd__nand2_1 _3811_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__o211a_1 _3812_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ),
    .A2(_0723_),
    .B1(_0725_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0726_));
 sky130_fd_sc_hd__nor2_1 _3813_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__a22o_4 _3814_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ),
    .A2(_0711_),
    .B1(_0727_),
    .B2(_0722_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ));
 sky130_fd_sc_hd__nand2b_1 _3815_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ),
    .B(net1059),
    .Y(_0728_));
 sky130_fd_sc_hd__o21ai_4 _3816_ (.A1(net1059),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ),
    .B1(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__or2_1 _3817_ (.A(net665),
    .B(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__xnor2_1 _3818_ (.A(_0679_),
    .B(_0680_),
    .Y(_0731_));
 sky130_fd_sc_hd__nor2_1 _3819_ (.A(_0730_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__mux4_2 _3820_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net16),
    .A2(net72),
    .A3(net108),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0733_));
 sky130_fd_sc_hd__mux4_1 _3821_ (.A0(net15),
    .A1(net107),
    .A2(net71),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _3822_ (.A0(_0734_),
    .A1(_0733_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0735_));
 sky130_fd_sc_hd__mux4_1 _3823_ (.A0(net25),
    .A1(net79),
    .A2(net104),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ),
    .X(_0736_));
 sky130_fd_sc_hd__mux4_2 _3824_ (.A0(net205),
    .A1(net63),
    .A2(net7),
    .A3(net99),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_1 _3825_ (.A0(_0737_),
    .A1(_0736_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_2 _3826_ (.A0(_0735_),
    .A1(_0738_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ));
 sky130_fd_sc_hd__nand2b_1 _3827_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ),
    .B(net1059),
    .Y(_0739_));
 sky130_fd_sc_hd__o21ai_4 _3828_ (.A1(net1059),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ),
    .B1(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__or2_1 _3829_ (.A(net665),
    .B(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__nor2_4 _3830_ (.A(net662),
    .B(_0661_),
    .Y(_0742_));
 sky130_fd_sc_hd__nor2_1 _3831_ (.A(_0620_),
    .B(_0729_),
    .Y(_0743_));
 sky130_fd_sc_hd__nand2_1 _3832_ (.A(_0679_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__xnor2_2 _3833_ (.A(_0621_),
    .B(_0742_),
    .Y(_0745_));
 sky130_fd_sc_hd__or2_4 _3834_ (.A(_0741_),
    .B(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__xnor2_1 _3835_ (.A(_0741_),
    .B(_0745_),
    .Y(_0747_));
 sky130_fd_sc_hd__o21ba_4 _3836_ (.A1(_0681_),
    .A2(_0732_),
    .B1_N(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__or3b_1 _3837_ (.A(_0681_),
    .B(_0732_),
    .C_N(_0747_),
    .X(_0749_));
 sky130_fd_sc_hd__nand2b_4 _3838_ (.A_N(_0748_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__or2_1 _3839_ (.A(_0578_),
    .B(_0579_),
    .X(_0751_));
 sky130_fd_sc_hd__nand2_1 _3840_ (.A(_0580_),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__nor2_4 _3841_ (.A(_0752_),
    .B(_0750_),
    .Y(_0753_));
 sky130_fd_sc_hd__or2_4 _3842_ (.A(_0543_),
    .B(net665),
    .X(_0754_));
 sky130_fd_sc_hd__nor2_1 _3843_ (.A(_0661_),
    .B(_0740_),
    .Y(_0755_));
 sky130_fd_sc_hd__nor2_1 _3844_ (.A(_0620_),
    .B(_0740_),
    .Y(_0756_));
 sky130_fd_sc_hd__xnor2_1 _3845_ (.A(_0743_),
    .B(_0755_),
    .Y(_0757_));
 sky130_fd_sc_hd__xnor2_4 _3846_ (.A(_0757_),
    .B(_0754_),
    .Y(_0758_));
 sky130_fd_sc_hd__nand3_4 _3847_ (.A(_0744_),
    .B(_0746_),
    .C(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__a21o_1 _3848_ (.A1(_0744_),
    .A2(_0746_),
    .B1(_0758_),
    .X(_0760_));
 sky130_fd_sc_hd__nand2_4 _3849_ (.A(_0760_),
    .B(_0759_),
    .Y(_0761_));
 sky130_fd_sc_hd__xnor2_2 _3850_ (.A(_0761_),
    .B(_0493_),
    .Y(_0762_));
 sky130_fd_sc_hd__nor3b_2 _3851_ (.A(_0748_),
    .B(_0753_),
    .C_N(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__o21ba_1 _3852_ (.A1(_0748_),
    .A2(_0753_),
    .B1_N(_0762_),
    .X(_0764_));
 sky130_fd_sc_hd__nor2_2 _3853_ (.A(_0764_),
    .B(_0763_),
    .Y(_0765_));
 sky130_fd_sc_hd__xnor2_2 _3854_ (.A(_0765_),
    .B(_0580_),
    .Y(_0766_));
 sky130_fd_sc_hd__mux4_2 _3855_ (.A0(net188),
    .A1(net134),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(net224),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0767_));
 sky130_fd_sc_hd__mux4_1 _3856_ (.A0(net972),
    .A1(net986),
    .A2(net990),
    .A3(net976),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0768_));
 sky130_fd_sc_hd__mux4_1 _3857_ (.A0(net982),
    .A1(net996),
    .A2(net1018),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0769_));
 sky130_fd_sc_hd__or2_1 _3858_ (.A(_0113_),
    .B(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__o21a_1 _3859_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .A2(_0768_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0771_));
 sky130_fd_sc_hd__mux4_1 _3860_ (.A0(net173),
    .A1(net179),
    .A2(net195),
    .A3(net125),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0772_));
 sky130_fd_sc_hd__mux4_1 _3861_ (.A0(net1216),
    .A1(net71),
    .A2(net215),
    .A3(net234),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _3862_ (.A0(_0772_),
    .A1(_0773_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _3863_ (.A1(_0770_),
    .A2(_0771_),
    .B1(_0774_),
    .B2(_0114_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _3864_ (.A0(net715),
    .A1(net995),
    .A2(net1016),
    .A3(net714),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0775_));
 sky130_fd_sc_hd__mux4_2 _3865_ (.A0(net971),
    .A1(net691),
    .A2(net707),
    .A3(net975),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_4 _3866_ (.A0(_0776_),
    .A1(_0775_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_0777_));
 sky130_fd_sc_hd__mux4_1 _3867_ (.A0(net175),
    .A1(net181),
    .A2(net193),
    .A3(net127),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0778_));
 sky130_fd_sc_hd__mux4_1 _3868_ (.A0(net1216),
    .A1(net73),
    .A2(net217),
    .A3(net229),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_1 _3869_ (.A0(_0778_),
    .A1(_0779_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_4 _3870_ (.A0(_0780_),
    .A1(_0777_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__mux4_2 _3871_ (.A0(net201),
    .A1(net71),
    .A2(net125),
    .A3(net215),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0781_));
 sky130_fd_sc_hd__mux4_2 _3872_ (.A0(net143),
    .A1(net83),
    .A2(net220),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .X(_0782_));
 sky130_fd_sc_hd__mux4_2 _3873_ (.A0(net133),
    .A1(net223),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0783_));
 sky130_fd_sc_hd__mux4_2 _3874_ (.A0(_0783_),
    .A1(_0781_),
    .A2(_0767_),
    .A3(_0782_),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ),
    .X(\Tile_X0Y1_DSP_bot.A1 ));
 sky130_fd_sc_hd__mux2_4 _3875_ (.A0(\Tile_X0Y1_DSP_bot.A1 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ),
    .S(net1060),
    .X(_0784_));
 sky130_fd_sc_hd__clkinv_2 _3876_ (.A(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__and3_1 _3877_ (.A(_0659_),
    .B(_0660_),
    .C(_0784_),
    .X(_0786_));
 sky130_fd_sc_hd__nor2_1 _3878_ (.A(_0620_),
    .B(_0785_),
    .Y(_0787_));
 sky130_fd_sc_hd__or2_1 _3879_ (.A(_0601_),
    .B(_0709_),
    .X(_0788_));
 sky130_fd_sc_hd__xnor2_1 _3880_ (.A(_0678_),
    .B(_0787_),
    .Y(_0789_));
 sky130_fd_sc_hd__o2bb2ai_1 _3881_ (.A1_N(_0680_),
    .A2_N(_0786_),
    .B1(_0788_),
    .B2(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__xnor2_1 _3882_ (.A(_0730_),
    .B(_0731_),
    .Y(_0791_));
 sky130_fd_sc_hd__and2b_1 _3883_ (.A_N(_0791_),
    .B(_0790_),
    .X(_0792_));
 sky130_fd_sc_hd__xor2_1 _3884_ (.A(_0790_),
    .B(_0791_),
    .X(_0793_));
 sky130_fd_sc_hd__mux4_1 _3885_ (.A0(net971),
    .A1(net967),
    .A2(net990),
    .A3(net976),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0794_));
 sky130_fd_sc_hd__or2_1 _3886_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .B(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__mux4_2 _3887_ (.A0(net982),
    .A1(net996),
    .A2(net1018),
    .A3(net1000),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0796_));
 sky130_fd_sc_hd__o21a_1 _3888_ (.A1(_0796_),
    .A2(_0118_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0797_));
 sky130_fd_sc_hd__mux4_1 _3889_ (.A0(net204),
    .A1(net120),
    .A2(net126),
    .A3(net1215),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0798_));
 sky130_fd_sc_hd__mux4_1 _3890_ (.A0(net72),
    .A1(net216),
    .A2(net84),
    .A3(net230),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0799_));
 sky130_fd_sc_hd__mux2_1 _3891_ (.A0(_0798_),
    .A1(_0799_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .X(_0800_));
 sky130_fd_sc_hd__a22o_4 _3892_ (.A1(_0797_),
    .A2(_0795_),
    .B1(_0800_),
    .B2(_0119_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _3893_ (.A0(net202),
    .A1(net142),
    .A2(net82),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .X(_0801_));
 sky130_fd_sc_hd__mux4_2 _3894_ (.A0(net181),
    .A1(net127),
    .A2(net91),
    .A3(net217),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_4 _3895_ (.A0(_0802_),
    .A1(_0801_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0803_));
 sky130_fd_sc_hd__and2_4 _3896_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .B(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _3897_ (.A0(net189),
    .A1(net135),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0805_));
 sky130_fd_sc_hd__mux4_2 _3898_ (.A0(net974),
    .A1(net970),
    .A2(net989),
    .A3(net994),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0806_));
 sky130_fd_sc_hd__or2_4 _3899_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .B(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__mux4_1 _3900_ (.A0(net984),
    .A1(net998),
    .A2(net1020),
    .A3(net1001),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0808_));
 sky130_fd_sc_hd__o211a_1 _3901_ (.A1(_0116_),
    .A2(_0808_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .C1(_0807_),
    .X(_0809_));
 sky130_fd_sc_hd__a211o_1 _3902_ (.A1(_0527_),
    .A2(_0528_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .C1(_0522_),
    .X(_0810_));
 sky130_fd_sc_hd__a21oi_1 _3903_ (.A1(_0061_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0811_));
 sky130_fd_sc_hd__mux2_1 _3904_ (.A0(net210),
    .A1(net1067),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0812_));
 sky130_fd_sc_hd__a221o_1 _3905_ (.A1(_0811_),
    .A2(_0810_),
    .B1(_0812_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .C1(_0116_),
    .X(_0813_));
 sky130_fd_sc_hd__mux4_1 _3906_ (.A0(net174),
    .A1(net182),
    .A2(net120),
    .A3(net128),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0814_));
 sky130_fd_sc_hd__o21ba_1 _3907_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0814_),
    .B1_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0815_));
 sky130_fd_sc_hd__a21o_1 _3908_ (.A1(_0813_),
    .A2(_0815_),
    .B1(_0809_),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__a211o_1 _3909_ (.A1(_0815_),
    .A2(_0813_),
    .B1(_0115_),
    .C1(_0809_),
    .X(_0816_));
 sky130_fd_sc_hd__o21a_1 _3910_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .X(_0817_));
 sky130_fd_sc_hd__a22o_4 _3911_ (.A1(_0117_),
    .A2(_0805_),
    .B1(_0817_),
    .B2(_0816_),
    .X(_0818_));
 sky130_fd_sc_hd__inv_2 _3912_ (.A(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__a221o_1 _3913_ (.A1(_0117_),
    .A2(_0805_),
    .B1(_0817_),
    .B2(_0816_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _3914_ (.A0(net190),
    .A1(net136),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .X(_0821_));
 sky130_fd_sc_hd__inv_1 _3915_ (.A(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__mux2_1 _3916_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A1(net226),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_1 _3917_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__o211a_1 _3918_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .A2(_0822_),
    .B1(_0824_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0825_));
 sky130_fd_sc_hd__nor2_1 _3919_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .B(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__a21o_1 _3920_ (.A1(_0820_),
    .A2(_0826_),
    .B1(_0804_),
    .X(\Tile_X0Y1_DSP_bot.B2 ));
 sky130_fd_sc_hd__a211o_4 _3921_ (.A1(_0820_),
    .A2(_0826_),
    .B1(_0804_),
    .C1(net1061),
    .X(_0827_));
 sky130_fd_sc_hd__nand2b_1 _3922_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ),
    .B(net1062),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2_8 _3923_ (.A(_0827_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__or2_4 _3924_ (.A(_0492_),
    .B(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__nor2_1 _3925_ (.A(_0450_),
    .B(_0740_),
    .Y(_0831_));
 sky130_fd_sc_hd__nor2_1 _3926_ (.A(_0576_),
    .B(_0740_),
    .Y(_0832_));
 sky130_fd_sc_hd__xnor2_1 _3927_ (.A(_0577_),
    .B(_0831_),
    .Y(_0833_));
 sky130_fd_sc_hd__xnor2_4 _3928_ (.A(_0830_),
    .B(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__o21ba_4 _3929_ (.A1(_0793_),
    .A2(_0834_),
    .B1_N(_0792_),
    .X(_0835_));
 sky130_fd_sc_hd__xor2_1 _3930_ (.A(_0750_),
    .B(_0752_),
    .X(_0836_));
 sky130_fd_sc_hd__nand2b_1 _3931_ (.A_N(_0835_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__o2bb2ai_1 _3932_ (.A1_N(_0577_),
    .A2_N(_0831_),
    .B1(_0833_),
    .B2(_0830_),
    .Y(_0838_));
 sky130_fd_sc_hd__xnor2_1 _3933_ (.A(_0835_),
    .B(_0836_),
    .Y(_0839_));
 sky130_fd_sc_hd__a21bo_4 _3934_ (.A1(_0838_),
    .A2(_0839_),
    .B1_N(_0837_),
    .X(_0840_));
 sky130_fd_sc_hd__nand2_4 _3935_ (.A(_0840_),
    .B(_0766_),
    .Y(_0841_));
 sky130_fd_sc_hd__or2_4 _3936_ (.A(_0492_),
    .B(_0709_),
    .X(_0842_));
 sky130_fd_sc_hd__nor2_1 _3937_ (.A(_0543_),
    .B(_0661_),
    .Y(_0843_));
 sky130_fd_sc_hd__nor2_1 _3938_ (.A(_0756_),
    .B(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__and2_1 _3939_ (.A(_0756_),
    .B(_0843_),
    .X(_0845_));
 sky130_fd_sc_hd__or2_1 _3940_ (.A(_0844_),
    .B(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__and2_1 _3941_ (.A(_0842_),
    .B(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__nor2_1 _3942_ (.A(_0842_),
    .B(_0846_),
    .Y(_0848_));
 sky130_fd_sc_hd__or2_4 _3943_ (.A(_0847_),
    .B(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__o2bb2ai_1 _3944_ (.A1_N(_0743_),
    .A2_N(_0755_),
    .B1(_0757_),
    .B2(_0754_),
    .Y(_0850_));
 sky130_fd_sc_hd__and2b_1 _3945_ (.A_N(_0849_),
    .B(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__xor2_1 _3946_ (.A(_0849_),
    .B(_0850_),
    .X(_0852_));
 sky130_fd_sc_hd__o21a_1 _3947_ (.A1(_0493_),
    .A2(_0761_),
    .B1(_0760_),
    .X(_0853_));
 sky130_fd_sc_hd__nor2_2 _3948_ (.A(_0852_),
    .B(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__xnor2_1 _3949_ (.A(_0852_),
    .B(_0853_),
    .Y(_0855_));
 sky130_fd_sc_hd__o21ba_1 _3950_ (.A1(_0580_),
    .A2(_0763_),
    .B1_N(_0764_),
    .X(_0856_));
 sky130_fd_sc_hd__nor2_1 _3951_ (.A(_0855_),
    .B(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__xnor2_1 _3952_ (.A(_0855_),
    .B(_0856_),
    .Y(_0858_));
 sky130_fd_sc_hd__nor2_1 _3953_ (.A(_0841_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__mux4_1 _3954_ (.A0(net183),
    .A1(net129),
    .A2(net92),
    .A3(net219),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(_0860_),
    .A1(net672),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_0861_));
 sky130_fd_sc_hd__mux4_2 _3956_ (.A0(net192),
    .A1(net138),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .A3(net228),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .X(_0862_));
 sky130_fd_sc_hd__mux4_1 _3957_ (.A0(net1012),
    .A1(net1047),
    .A2(net1028),
    .A3(net1052),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0863_));
 sky130_fd_sc_hd__mux4_1 _3958_ (.A0(net1043),
    .A1(net1032),
    .A2(net1038),
    .A3(net1055),
    .S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0864_));
 sky130_fd_sc_hd__and2_1 _3959_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .B(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__a21bo_1 _3960_ (.A1(_0096_),
    .A2(_0863_),
    .B1_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ),
    .X(_0866_));
 sky130_fd_sc_hd__mux2_1 _3961_ (.A0(net673),
    .A1(net192),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _3962_ (.A0(net1257),
    .A1(net12),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0868_));
 sky130_fd_sc_hd__or2_1 _3963_ (.A(_0095_),
    .B(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__o211a_1 _3964_ (.A1(_0867_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .B1(_0869_),
    .C1(_0096_),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _3965_ (.A0(net60),
    .A1(net68),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0871_));
 sky130_fd_sc_hd__or2_1 _3966_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .B(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _3967_ (.A0(net94),
    .A1(net1219),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0873_));
 sky130_fd_sc_hd__o211a_1 _3968_ (.A1(_0095_),
    .A2(_0873_),
    .B1(_0872_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0874_));
 sky130_fd_sc_hd__o32a_4 _3969_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0870_),
    .A3(_0874_),
    .B1(_0865_),
    .B2(_0866_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _3970_ (.A0(net191),
    .A1(net227),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .A3(net658),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_4 _3971_ (.A0(_0875_),
    .A1(_0862_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_4 _3972_ (.A0(_0876_),
    .A1(_0861_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ),
    .X(\Tile_X0Y1_DSP_bot.A0 ));
 sky130_fd_sc_hd__nand2b_1 _3973_ (.A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ),
    .B(net1059),
    .Y(_0877_));
 sky130_fd_sc_hd__o21ai_4 _3974_ (.A1(\Tile_X0Y1_DSP_bot.A0 ),
    .A2(net1059),
    .B1(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__nor2_1 _3975_ (.A(_0620_),
    .B(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__nor2_1 _3976_ (.A(_0676_),
    .B(_0709_),
    .Y(_0880_));
 sky130_fd_sc_hd__inv_2 _3977_ (.A(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__xnor2_1 _3978_ (.A(_0786_),
    .B(_0879_),
    .Y(_0882_));
 sky130_fd_sc_hd__o2bb2a_1 _3979_ (.A1_N(_0786_),
    .A2_N(_0879_),
    .B1(_0881_),
    .B2(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__xnor2_1 _3980_ (.A(_0788_),
    .B(_0789_),
    .Y(_0884_));
 sky130_fd_sc_hd__or2_1 _3981_ (.A(_0883_),
    .B(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__xnor2_1 _3982_ (.A(_0883_),
    .B(_0884_),
    .Y(_0886_));
 sky130_fd_sc_hd__or2_1 _3983_ (.A(_0543_),
    .B(_0829_),
    .X(_0887_));
 sky130_fd_sc_hd__nor2_1 _3984_ (.A(_0450_),
    .B(_0729_),
    .Y(_0888_));
 sky130_fd_sc_hd__nor2_1 _3985_ (.A(_0576_),
    .B(_0729_),
    .Y(_0889_));
 sky130_fd_sc_hd__xnor2_1 _3986_ (.A(_0832_),
    .B(_0888_),
    .Y(_0890_));
 sky130_fd_sc_hd__xnor2_1 _3987_ (.A(_0887_),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__o21a_1 _3988_ (.A1(_0886_),
    .A2(_0891_),
    .B1(_0885_),
    .X(_0892_));
 sky130_fd_sc_hd__xor2_1 _3989_ (.A(_0793_),
    .B(_0834_),
    .X(_0893_));
 sky130_fd_sc_hd__nand2b_1 _3990_ (.A_N(_0892_),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__o2bb2ai_1 _3991_ (.A1_N(_0832_),
    .A2_N(_0888_),
    .B1(_0890_),
    .B2(_0887_),
    .Y(_0895_));
 sky130_fd_sc_hd__xnor2_1 _3992_ (.A(_0892_),
    .B(_0893_),
    .Y(_0896_));
 sky130_fd_sc_hd__a21bo_1 _3993_ (.A1(_0895_),
    .A2(_0896_),
    .B1_N(_0894_),
    .X(_0897_));
 sky130_fd_sc_hd__xnor2_1 _3994_ (.A(_0838_),
    .B(_0839_),
    .Y(_0898_));
 sky130_fd_sc_hd__and2b_1 _3995_ (.A_N(_0898_),
    .B(_0897_),
    .X(_0899_));
 sky130_fd_sc_hd__xor2_1 _3996_ (.A(_0766_),
    .B(_0840_),
    .X(_0900_));
 sky130_fd_sc_hd__and2_4 _3997_ (.A(_0899_),
    .B(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__nor2_1 _3998_ (.A(_0899_),
    .B(_0900_),
    .Y(_0902_));
 sky130_fd_sc_hd__nor2_1 _3999_ (.A(_0901_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__xnor2_1 _4000_ (.A(_0897_),
    .B(_0898_),
    .Y(_0904_));
 sky130_fd_sc_hd__nor2_1 _4001_ (.A(_0709_),
    .B(_0878_),
    .Y(_0905_));
 sky130_fd_sc_hd__nand2_1 _4002_ (.A(_0786_),
    .B(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__xnor2_1 _4003_ (.A(_0881_),
    .B(_0882_),
    .Y(_0907_));
 sky130_fd_sc_hd__nor2_1 _4004_ (.A(_0906_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__xor2_1 _4005_ (.A(_0906_),
    .B(_0907_),
    .X(_0909_));
 sky130_fd_sc_hd__dlxtp_1 _4006_ (.D(net1228),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4007_ (.D(net1229),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4008_ (.D(net46),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4009_ (.D(net1232),
    .GATE(net1178),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4010_ (.D(net1234),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4011_ (.D(net1236),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4012_ (.D(net44),
    .GATE(net1178),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4013_ (.D(net1238),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4014_ (.D(net1239),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4015_ (.D(net1240),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4016_ (.D(net1241),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4017_ (.D(net1242),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4018_ (.D(net1244),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4019_ (.D(net1245),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4020_ (.D(net1246),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4021_ (.D(net1247),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4022_ (.D(net1248),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4023_ (.D(net1249),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4024_ (.D(net1250),
    .GATE(net1178),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4025_ (.D(net1251),
    .GATE(net1178),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4026_ (.D(net1252),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4027_ (.D(net1253),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4028_ (.D(net1221),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4029_ (.D(net55),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4030_ (.D(net1223),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4031_ (.D(net1224),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4032_ (.D(net1225),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4033_ (.D(net1226),
    .GATE(net1175),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4034_ (.D(net1227),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4035_ (.D(net1230),
    .GATE(net1177),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4036_ (.D(net38),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4037_ (.D(net27),
    .GATE(net1176),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4038_ (.D(net49),
    .GATE(net1143),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4039_ (.D(net1229),
    .GATE(net1144),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4040_ (.D(net1231),
    .GATE(net1143),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4041_ (.D(net1232),
    .GATE(net1143),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4042_ (.D(net1233),
    .GATE(net1143),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4043_ (.D(net1235),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4044_ (.D(net44),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4045_ (.D(net43),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4046_ (.D(net1239),
    .GATE(net1143),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4047_ (.D(net1240),
    .GATE(net1143),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4048_ (.D(net1241),
    .GATE(net1143),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4049_ (.D(net1242),
    .GATE(net1143),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4050_ (.D(net1244),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4051_ (.D(net1245),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4052_ (.D(net35),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4053_ (.D(net1247),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4054_ (.D(net1248),
    .GATE(net1144),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4055_ (.D(net1249),
    .GATE(net1144),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4056_ (.D(net1250),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4057_ (.D(net1251),
    .GATE(net1144),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4058_ (.D(net1252),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4059_ (.D(net1253),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4060_ (.D(net1221),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4061_ (.D(net1222),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4062_ (.D(net1223),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4063_ (.D(net1224),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4064_ (.D(net1225),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4065_ (.D(net1226),
    .GATE(net1141),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4066_ (.D(net1227),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4067_ (.D(net1230),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4068_ (.D(net1243),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4069_ (.D(net1254),
    .GATE(net1142),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4070_ (.D(net1228),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4071_ (.D(net1229),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4072_ (.D(net1231),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4073_ (.D(net1232),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4074_ (.D(net1233),
    .GATE(net1135),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4075_ (.D(net1235),
    .GATE(net1135),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4076_ (.D(net44),
    .GATE(net1135),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4077_ (.D(net43),
    .GATE(net1135),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4078_ (.D(net1239),
    .GATE(net1135),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4079_ (.D(net1240),
    .GATE(net1135),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4080_ (.D(net1241),
    .GATE(net1135),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4081_ (.D(net1242),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4082_ (.D(net1244),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4083_ (.D(net1245),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4084_ (.D(net1246),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4085_ (.D(net1247),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4086_ (.D(net1248),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4087_ (.D(net1249),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4088_ (.D(net31),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4089_ (.D(net30),
    .GATE(net1134),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4090_ (.D(net29),
    .GATE(net1133),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4091_ (.D(net28),
    .GATE(net1133),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4092_ (.D(net1221),
    .GATE(net1133),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4093_ (.D(net1222),
    .GATE(net1133),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4094_ (.D(net1223),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4095_ (.D(net1224),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4096_ (.D(net1225),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4097_ (.D(net1226),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4098_ (.D(net1227),
    .GATE(net1133),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4099_ (.D(net1230),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4100_ (.D(net1243),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4101_ (.D(net1254),
    .GATE(net1132),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4102_ (.D(net1228),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4103_ (.D(net48),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4104_ (.D(net1231),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4105_ (.D(net1232),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4106_ (.D(net1234),
    .GATE(net1126),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4107_ (.D(net1235),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4108_ (.D(net1237),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4109_ (.D(net1238),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4110_ (.D(net1239),
    .GATE(net1126),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4111_ (.D(net1240),
    .GATE(net1126),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4112_ (.D(net40),
    .GATE(net1126),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4113_ (.D(net1242),
    .GATE(net1126),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4114_ (.D(net37),
    .GATE(net1127),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4115_ (.D(net36),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4116_ (.D(net1246),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4117_ (.D(net34),
    .GATE(net1125),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4118_ (.D(net1248),
    .GATE(net1124),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4119_ (.D(net1249),
    .GATE(net1124),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4120_ (.D(net1250),
    .GATE(net1124),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4121_ (.D(net1251),
    .GATE(net1124),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4122_ (.D(net1252),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4123_ (.D(net1253),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4124_ (.D(net1221),
    .GATE(net1124),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4125_ (.D(net1222),
    .GATE(net1124),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4126_ (.D(net1223),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4127_ (.D(net1224),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4128_ (.D(net1225),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4129_ (.D(net1226),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4130_ (.D(net1227),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4131_ (.D(net1230),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4132_ (.D(net1243),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4133_ (.D(net1254),
    .GATE(net1123),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4134_ (.D(net49),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4135_ (.D(net48),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4136_ (.D(net1231),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4137_ (.D(net1232),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4138_ (.D(net1233),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4139_ (.D(net1235),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4140_ (.D(net44),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4141_ (.D(net43),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4142_ (.D(net42),
    .GATE(net1117),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4143_ (.D(net41),
    .GATE(net1117),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4144_ (.D(net1241),
    .GATE(net1117),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4145_ (.D(net1242),
    .GATE(net1117),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4146_ (.D(net1244),
    .GATE(net1117),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4147_ (.D(net1245),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4148_ (.D(net35),
    .GATE(net1117),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4149_ (.D(net34),
    .GATE(net1115),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4150_ (.D(net1248),
    .GATE(net1118),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4151_ (.D(net1249),
    .GATE(net1118),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4152_ (.D(net31),
    .GATE(net1118),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4153_ (.D(net30),
    .GATE(net1118),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4154_ (.D(net1252),
    .GATE(net1116),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4155_ (.D(net1253),
    .GATE(net1116),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4156_ (.D(net56),
    .GATE(net1116),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4157_ (.D(net1222),
    .GATE(net1116),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4158_ (.D(net54),
    .GATE(net1116),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4159_ (.D(net53),
    .GATE(net1118),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4160_ (.D(net1225),
    .GATE(net1118),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4161_ (.D(net1226),
    .GATE(net1118),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4162_ (.D(net1227),
    .GATE(net1116),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4163_ (.D(net1230),
    .GATE(net1116),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4164_ (.D(net1243),
    .GATE(net1116),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4165_ (.D(net1254),
    .GATE(net1116),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4166_ (.D(net1228),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4167_ (.D(net1229),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4168_ (.D(net46),
    .GATE(net1108),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4169_ (.D(net1232),
    .GATE(net1108),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4170_ (.D(net1233),
    .GATE(net1108),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4171_ (.D(net1235),
    .GATE(net1108),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4172_ (.D(net1237),
    .GATE(net1109),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4173_ (.D(net1238),
    .GATE(net1109),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4174_ (.D(net1239),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4175_ (.D(net1240),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4176_ (.D(net1241),
    .GATE(net1109),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4177_ (.D(net1242),
    .GATE(net1108),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4178_ (.D(net1244),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4179_ (.D(net1245),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4180_ (.D(net1246),
    .GATE(net1108),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4181_ (.D(net1247),
    .GATE(net1108),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4182_ (.D(net33),
    .GATE(net1110),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4183_ (.D(net32),
    .GATE(net1110),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4184_ (.D(net1250),
    .GATE(net1110),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4185_ (.D(net1251),
    .GATE(net1110),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4186_ (.D(net1252),
    .GATE(net1108),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4187_ (.D(net1253),
    .GATE(net1108),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4188_ (.D(net56),
    .GATE(net1109),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4189_ (.D(net55),
    .GATE(net1109),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4190_ (.D(net54),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4191_ (.D(net53),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4192_ (.D(net1225),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4193_ (.D(net51),
    .GATE(net1107),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4194_ (.D(net1227),
    .GATE(net1110),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4195_ (.D(net1230),
    .GATE(net1110),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4196_ (.D(net38),
    .GATE(net1109),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4197_ (.D(net27),
    .GATE(net1109),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4198_ (.D(net1228),
    .GATE(net1101),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4199_ (.D(net1229),
    .GATE(net1101),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4200_ (.D(net1231),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4201_ (.D(net1232),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4202_ (.D(net1233),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4203_ (.D(net1235),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4204_ (.D(net1237),
    .GATE(net1100),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4205_ (.D(net1238),
    .GATE(net1100),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4206_ (.D(net42),
    .GATE(net1100),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4207_ (.D(net41),
    .GATE(net1101),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4208_ (.D(net1241),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4209_ (.D(net1242),
    .GATE(net1102),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4210_ (.D(net1244),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4211_ (.D(net1245),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4212_ (.D(net1246),
    .GATE(net1101),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4213_ (.D(net1247),
    .GATE(net1101),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4214_ (.D(net1248),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4215_ (.D(net1249),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4216_ (.D(net1250),
    .GATE(net1101),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4217_ (.D(net1251),
    .GATE(net1101),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4218_ (.D(net29),
    .GATE(net1100),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4219_ (.D(net28),
    .GATE(net1100),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4220_ (.D(net56),
    .GATE(net1100),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4221_ (.D(net55),
    .GATE(net1100),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4222_ (.D(net1223),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4223_ (.D(net1224),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4224_ (.D(net1225),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4225_ (.D(net1226),
    .GATE(net1099),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4226_ (.D(net50),
    .GATE(net1100),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4227_ (.D(net47),
    .GATE(net1100),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4228_ (.D(net38),
    .GATE(net1101),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4229_ (.D(net27),
    .GATE(net1101),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4230_ (.D(net1228),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4231_ (.D(net1229),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4232_ (.D(net1231),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4233_ (.D(net45),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4234_ (.D(net1233),
    .GATE(net1091),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4235_ (.D(net1236),
    .GATE(net1091),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4236_ (.D(net1237),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4237_ (.D(net1238),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4238_ (.D(net42),
    .GATE(net1091),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4239_ (.D(net41),
    .GATE(net1091),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4240_ (.D(net1241),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4241_ (.D(net1242),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4242_ (.D(net37),
    .GATE(net1091),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4243_ (.D(net36),
    .GATE(net1091),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4244_ (.D(net35),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4245_ (.D(net34),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4246_ (.D(net33),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4247_ (.D(net32),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4248_ (.D(net1250),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4249_ (.D(net1251),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4250_ (.D(net1252),
    .GATE(net1091),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4251_ (.D(net1253),
    .GATE(net1091),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4252_ (.D(net1221),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4253_ (.D(net1222),
    .GATE(net1090),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4254_ (.D(net1223),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4255_ (.D(net1224),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4256_ (.D(net52),
    .GATE(net1092),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4257_ (.D(net51),
    .GATE(net1092),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4258_ (.D(net1227),
    .GATE(net1092),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4259_ (.D(net1230),
    .GATE(net1092),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4260_ (.D(net1243),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4261_ (.D(net1254),
    .GATE(net1093),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4262_ (.D(net1228),
    .GATE(net1085),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4263_ (.D(net1229),
    .GATE(net1084),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4264_ (.D(net46),
    .GATE(net1084),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4265_ (.D(net45),
    .GATE(net1084),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4266_ (.D(net1234),
    .GATE(net1084),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4267_ (.D(net1235),
    .GATE(net1084),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4268_ (.D(net1237),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4269_ (.D(net1238),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4270_ (.D(net1239),
    .GATE(net1084),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4271_ (.D(net1240),
    .GATE(net1084),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4272_ (.D(net40),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4273_ (.D(net39),
    .GATE(net1083),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4274_ (.D(net1244),
    .GATE(net1083),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4275_ (.D(net1245),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4276_ (.D(net1246),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4277_ (.D(net1247),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4278_ (.D(net1248),
    .GATE(net1084),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4279_ (.D(net1249),
    .GATE(net1084),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4280_ (.D(net1250),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4281_ (.D(net1251),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4282_ (.D(net29),
    .GATE(net1083),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4283_ (.D(net28),
    .GATE(net1083),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4284_ (.D(net1221),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4285_ (.D(net1222),
    .GATE(net1082),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4286_ (.D(net1223),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4287_ (.D(net1224),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4288_ (.D(net52),
    .GATE(net1083),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4289_ (.D(net1226),
    .GATE(net1083),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4290_ (.D(net50),
    .GATE(net1083),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4291_ (.D(net47),
    .GATE(net1083),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4292_ (.D(net1243),
    .GATE(net1081),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4293_ (.D(net1254),
    .GATE(net1085),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4294_ (.D(net1228),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4295_ (.D(net1229),
    .GATE(net1074),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4296_ (.D(net1231),
    .GATE(net1074),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4297_ (.D(net1232),
    .GATE(net1077),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4298_ (.D(net1234),
    .GATE(net1074),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4299_ (.D(net1236),
    .GATE(net1074),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4300_ (.D(net1237),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4301_ (.D(net43),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4302_ (.D(net1239),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4303_ (.D(net1240),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4304_ (.D(net1241),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4305_ (.D(net1242),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4306_ (.D(net1244),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4307_ (.D(net1245),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4308_ (.D(net35),
    .GATE(net1076),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4309_ (.D(net34),
    .GATE(net1076),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4310_ (.D(net1248),
    .GATE(net1076),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4311_ (.D(net1249),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4312_ (.D(net1250),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4313_ (.D(net1251),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4314_ (.D(net1252),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4315_ (.D(net1253),
    .GATE(net1076),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4316_ (.D(net1221),
    .GATE(net1075),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4317_ (.D(net1222),
    .GATE(net1076),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4318_ (.D(net1223),
    .GATE(net1076),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4319_ (.D(net1224),
    .GATE(net1076),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4320_ (.D(net1225),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4321_ (.D(net1226),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4322_ (.D(net1227),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4323_ (.D(net1230),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4324_ (.D(net1243),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4325_ (.D(net1254),
    .GATE(net1073),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4326_ (.D(net1228),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4327_ (.D(net1229),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4328_ (.D(net1231),
    .GATE(net1169),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4329_ (.D(net1232),
    .GATE(net1169),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4330_ (.D(net1233),
    .GATE(net1169),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4331_ (.D(net1236),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4332_ (.D(net1237),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4333_ (.D(net1238),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4334_ (.D(net1239),
    .GATE(net1170),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4335_ (.D(net1240),
    .GATE(net1169),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4336_ (.D(net1241),
    .GATE(net1169),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4337_ (.D(net39),
    .GATE(net1170),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4338_ (.D(net37),
    .GATE(net1169),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4339_ (.D(net1245),
    .GATE(net1169),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4340_ (.D(net1246),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4341_ (.D(net1247),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4342_ (.D(net33),
    .GATE(net1170),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4343_ (.D(net32),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4344_ (.D(net1250),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4345_ (.D(net1251),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4346_ (.D(net1252),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4347_ (.D(net1253),
    .GATE(net1167),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4348_ (.D(net1221),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4349_ (.D(net1222),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4350_ (.D(net1223),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4351_ (.D(net1224),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4352_ (.D(net1225),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4353_ (.D(net1226),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4354_ (.D(net1227),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4355_ (.D(net1230),
    .GATE(net1168),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4356_ (.D(net1243),
    .GATE(net1169),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4357_ (.D(net1254),
    .GATE(net1169),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4358_ (.D(net49),
    .GATE(net1160),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4359_ (.D(net48),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4360_ (.D(net46),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4361_ (.D(net45),
    .GATE(net1160),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4362_ (.D(net1233),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4363_ (.D(net1235),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4364_ (.D(net1237),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4365_ (.D(net1238),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4366_ (.D(net1239),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4367_ (.D(net41),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4368_ (.D(net40),
    .GATE(net1161),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4369_ (.D(net39),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4370_ (.D(net37),
    .GATE(net1160),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4371_ (.D(net36),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4372_ (.D(net1246),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4373_ (.D(net1247),
    .GATE(net1160),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4374_ (.D(net1248),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4375_ (.D(net1249),
    .GATE(net1159),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4376_ (.D(net1250),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4377_ (.D(net30),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4378_ (.D(net29),
    .GATE(net1162),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4379_ (.D(net28),
    .GATE(net1162),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4380_ (.D(net1221),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4381_ (.D(net1222),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4382_ (.D(net1223),
    .GATE(net1162),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4383_ (.D(net1224),
    .GATE(net1162),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4384_ (.D(net52),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4385_ (.D(net1226),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4386_ (.D(net1227),
    .GATE(net1158),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4387_ (.D(net1230),
    .GATE(net1161),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4388_ (.D(net1243),
    .GATE(net1161),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4389_ (.D(net1254),
    .GATE(net1161),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4390_ (.D(net49),
    .GATE(net1151),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4391_ (.D(net48),
    .GATE(net1151),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4392_ (.D(net1231),
    .GATE(net1151),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4393_ (.D(net1232),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4394_ (.D(net1233),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4395_ (.D(net1235),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4396_ (.D(net1237),
    .GATE(net1152),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4397_ (.D(net1238),
    .GATE(net1152),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4398_ (.D(net1239),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4399_ (.D(net1240),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4400_ (.D(net1241),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4401_ (.D(net1242),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4402_ (.D(net1244),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4403_ (.D(net1245),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4404_ (.D(net1246),
    .GATE(net1152),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4405_ (.D(net1247),
    .GATE(net1152),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4406_ (.D(net1248),
    .GATE(net1152),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4407_ (.D(net1249),
    .GATE(net1152),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4408_ (.D(net31),
    .GATE(net1151),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4409_ (.D(net1251),
    .GATE(net1150),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4410_ (.D(net1252),
    .GATE(net1152),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4411_ (.D(net1253),
    .GATE(net1152),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ));
 sky130_fd_sc_hd__dfxtp_1 _4412_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0000_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4413_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0001_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4414_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0002_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4415_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0003_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4416_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0004_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4417_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0005_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4418_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0006_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4419_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0007_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4420_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0008_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4421_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0009_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4422_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0010_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4423_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0011_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4424_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0012_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4425_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0013_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4426_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0014_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4427_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0015_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4428_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0016_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4429_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0017_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4430_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0018_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4431_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(_0019_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4432_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(net735),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4433_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.A1 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4434_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.A2 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4435_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.A3 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4436_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4437_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4438_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4439_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4440_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.B0 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4441_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.B1 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4442_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.B2 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4443_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.B3 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4444_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4445_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4446_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4447_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4448_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C0 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4449_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C1 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4450_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C2 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4451_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C3 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4452_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C4 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4453_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C5 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4454_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C6 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4455_ (.CLK(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C7 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4456_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C8 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4457_ (.CLK(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y1_DSP_bot.C9 ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4458_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4459_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4460_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4461_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4462_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4463_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4464_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4465_ (.CLK(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4466_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4467_ (.CLK(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ));
 sky130_fd_sc_hd__dlxtp_1 _4468_ (.D(net1186),
    .GATE(net1173),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4469_ (.D(net1188),
    .GATE(net1173),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4470_ (.D(net164),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4471_ (.D(net163),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4472_ (.D(net1193),
    .GATE(net1174),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4473_ (.D(net1195),
    .GATE(net1174),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4474_ (.D(net1196),
    .GATE(net1174),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4475_ (.D(net1197),
    .GATE(net1174),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4476_ (.D(net1198),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4477_ (.D(net1199),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4478_ (.D(net1200),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4479_ (.D(net1201),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4480_ (.D(net1203),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4481_ (.D(net1204),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4482_ (.D(net1205),
    .GATE(net1174),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4483_ (.D(net1206),
    .GATE(net1174),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4484_ (.D(net1208),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4485_ (.D(net1209),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4486_ (.D(net1210),
    .GATE(net1173),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4487_ (.D(net1211),
    .GATE(net1173),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4488_ (.D(net1212),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4489_ (.D(net1213),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4490_ (.D(net172),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4491_ (.D(net1180),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4492_ (.D(net1181),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4493_ (.D(net1182),
    .GATE(net1171),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4494_ (.D(net1183),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4495_ (.D(net1184),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4496_ (.D(net1185),
    .GATE(net1173),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4497_ (.D(net1190),
    .GATE(net1173),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4498_ (.D(net155),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4499_ (.D(net145),
    .GATE(net1172),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4500_ (.D(net1186),
    .GATE(net1139),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4501_ (.D(net1188),
    .GATE(net1139),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4502_ (.D(net1191),
    .GATE(net1139),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4503_ (.D(net1192),
    .GATE(net1139),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4504_ (.D(net1194),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4505_ (.D(net1195),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4506_ (.D(net1196),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4507_ (.D(net1197),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4508_ (.D(net1198),
    .GATE(net1139),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4509_ (.D(net1199),
    .GATE(net1139),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4510_ (.D(net1200),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4511_ (.D(net1201),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4512_ (.D(net1203),
    .GATE(net1140),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4513_ (.D(net1204),
    .GATE(net1140),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4514_ (.D(net1205),
    .GATE(net1140),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4515_ (.D(net1206),
    .GATE(net1140),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4516_ (.D(net1208),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4517_ (.D(net1209),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4518_ (.D(net1210),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4519_ (.D(net1211),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4520_ (.D(net1212),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4521_ (.D(net1213),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4522_ (.D(net1179),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4523_ (.D(net1180),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4524_ (.D(net170),
    .GATE(net1145),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4525_ (.D(net169),
    .GATE(net1145),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4526_ (.D(net1183),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4527_ (.D(net167),
    .GATE(net1137),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4528_ (.D(net1185),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4529_ (.D(net1190),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4530_ (.D(net1202),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4531_ (.D(net1214),
    .GATE(net1138),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4532_ (.D(net1187),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4533_ (.D(net1189),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4534_ (.D(net1191),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4535_ (.D(net1192),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4536_ (.D(net1193),
    .GATE(net1131),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4537_ (.D(net1195),
    .GATE(net1131),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4538_ (.D(net1196),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4539_ (.D(net1197),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4540_ (.D(net1198),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4541_ (.D(net1199),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4542_ (.D(net1200),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4543_ (.D(net1201),
    .GATE(net1130),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4544_ (.D(net154),
    .GATE(net1131),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4545_ (.D(net153),
    .GATE(net1131),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4546_ (.D(net152),
    .GATE(net1131),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4547_ (.D(net1207),
    .GATE(net1131),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4548_ (.D(net1208),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4549_ (.D(net1209),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4550_ (.D(net1210),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4551_ (.D(net1211),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4552_ (.D(net147),
    .GATE(net1129),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4553_ (.D(net146),
    .GATE(net1129),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4554_ (.D(net172),
    .GATE(net1129),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4555_ (.D(net171),
    .GATE(net1129),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4556_ (.D(net1181),
    .GATE(net1129),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4557_ (.D(net1182),
    .GATE(net1129),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4558_ (.D(net1183),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4559_ (.D(net1184),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4560_ (.D(net1185),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4561_ (.D(net1190),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4562_ (.D(net1202),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4563_ (.D(net1214),
    .GATE(net1128),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4564_ (.D(net1186),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4565_ (.D(net1188),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4566_ (.D(net1191),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4567_ (.D(net1192),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4568_ (.D(net1193),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4569_ (.D(net1195),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4570_ (.D(net1196),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4571_ (.D(net1197),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4572_ (.D(net159),
    .GATE(net1122),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4573_ (.D(net158),
    .GATE(net1122),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4574_ (.D(net157),
    .GATE(net1122),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4575_ (.D(net156),
    .GATE(net1122),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4576_ (.D(net1203),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4577_ (.D(net1204),
    .GATE(net1122),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4578_ (.D(net1205),
    .GATE(net1121),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4579_ (.D(net1206),
    .GATE(net1122),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4580_ (.D(net1208),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4581_ (.D(net1209),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4582_ (.D(net1210),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4583_ (.D(net1211),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4584_ (.D(net1212),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4585_ (.D(net1213),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4586_ (.D(net1179),
    .GATE(net1120),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4587_ (.D(net1180),
    .GATE(net1120),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4588_ (.D(net170),
    .GATE(net1120),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4589_ (.D(net169),
    .GATE(net1120),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4590_ (.D(net1183),
    .GATE(net1120),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4591_ (.D(net1184),
    .GATE(net1120),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4592_ (.D(net1185),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4593_ (.D(net1190),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4594_ (.D(net1202),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4595_ (.D(net1214),
    .GATE(net1119),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4596_ (.D(net1186),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4597_ (.D(net1188),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4598_ (.D(net1191),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4599_ (.D(net1192),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4600_ (.D(net1193),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4601_ (.D(net1195),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4602_ (.D(net1196),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4603_ (.D(net1197),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4604_ (.D(net1198),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4605_ (.D(net1199),
    .GATE(net1114),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4606_ (.D(net1200),
    .GATE(net1114),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4607_ (.D(net1201),
    .GATE(net1113),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4608_ (.D(net154),
    .GATE(net1114),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4609_ (.D(net153),
    .GATE(net1114),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4610_ (.D(net152),
    .GATE(net1114),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4611_ (.D(net1207),
    .GATE(net1114),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4612_ (.D(net1208),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4613_ (.D(net1209),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4614_ (.D(net1210),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4615_ (.D(net1211),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4616_ (.D(net147),
    .GATE(net1112),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4617_ (.D(net146),
    .GATE(net1112),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4618_ (.D(net172),
    .GATE(net1112),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4619_ (.D(net171),
    .GATE(net1112),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4620_ (.D(net1181),
    .GATE(net1112),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4621_ (.D(net1182),
    .GATE(net1112),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4622_ (.D(net1183),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4623_ (.D(net1184),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4624_ (.D(net1185),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4625_ (.D(net1190),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4626_ (.D(net1202),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4627_ (.D(net1214),
    .GATE(net1111),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4628_ (.D(net1186),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4629_ (.D(net1188),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4630_ (.D(net1191),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4631_ (.D(net1192),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4632_ (.D(net1193),
    .GATE(net1106),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4633_ (.D(net1195),
    .GATE(net1106),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4634_ (.D(net1196),
    .GATE(net1106),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4635_ (.D(net1197),
    .GATE(net1106),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4636_ (.D(net1198),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4637_ (.D(net1199),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4638_ (.D(net157),
    .GATE(net1105),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4639_ (.D(net156),
    .GATE(net1105),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4640_ (.D(net1203),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4641_ (.D(net1204),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4642_ (.D(net1205),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4643_ (.D(net1207),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4644_ (.D(net1208),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4645_ (.D(net1209),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4646_ (.D(net1210),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4647_ (.D(net1211),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4648_ (.D(net1212),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4649_ (.D(net1213),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4650_ (.D(net1179),
    .GATE(net1105),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4651_ (.D(net171),
    .GATE(net1105),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4652_ (.D(net1181),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4653_ (.D(net1182),
    .GATE(net1103),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4654_ (.D(net1183),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4655_ (.D(net1184),
    .GATE(net1104),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4656_ (.D(net1185),
    .GATE(net1105),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4657_ (.D(net1190),
    .GATE(net1105),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4658_ (.D(net155),
    .GATE(net1105),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4659_ (.D(net1214),
    .GATE(net1105),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4660_ (.D(net1186),
    .GATE(net1095),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4661_ (.D(net1188),
    .GATE(net1095),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4662_ (.D(net164),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4663_ (.D(net163),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4664_ (.D(net1193),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4665_ (.D(net1195),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4666_ (.D(net161),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4667_ (.D(net160),
    .GATE(net1098),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4668_ (.D(net1198),
    .GATE(net1095),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4669_ (.D(net1199),
    .GATE(net1095),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4670_ (.D(net157),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4671_ (.D(net156),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4672_ (.D(net1203),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4673_ (.D(net1204),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4674_ (.D(net1205),
    .GATE(net1096),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4675_ (.D(net1206),
    .GATE(net1096),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4676_ (.D(net1208),
    .GATE(net1096),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4677_ (.D(net1209),
    .GATE(net1096),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4678_ (.D(net149),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4679_ (.D(net148),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4680_ (.D(net1212),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4681_ (.D(net1213),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4682_ (.D(net1179),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4683_ (.D(net1180),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4684_ (.D(net1181),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4685_ (.D(net1182),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4686_ (.D(net168),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4687_ (.D(net167),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4688_ (.D(net1185),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4689_ (.D(net1190),
    .GATE(net1094),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4690_ (.D(net1202),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4691_ (.D(net1214),
    .GATE(net1097),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4692_ (.D(net1186),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4693_ (.D(net1188),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4694_ (.D(net1191),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4695_ (.D(net1192),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4696_ (.D(net1193),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4697_ (.D(net1195),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4698_ (.D(net161),
    .GATE(net1089),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4699_ (.D(net160),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4700_ (.D(net1198),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4701_ (.D(net1199),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4702_ (.D(net1200),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4703_ (.D(net1201),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4704_ (.D(net1203),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4705_ (.D(net1204),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4706_ (.D(net1205),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4707_ (.D(net1206),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4708_ (.D(net151),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4709_ (.D(net150),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4710_ (.D(net1210),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4711_ (.D(net148),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4712_ (.D(net1212),
    .GATE(net1089),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4713_ (.D(net1213),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4714_ (.D(net1179),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4715_ (.D(net1180),
    .GATE(net1088),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4716_ (.D(net1181),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4717_ (.D(net1182),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4718_ (.D(net1183),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4719_ (.D(net1184),
    .GATE(net1086),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4720_ (.D(net166),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4721_ (.D(net165),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4722_ (.D(net1202),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4723_ (.D(net145),
    .GATE(net1087),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4724_ (.D(net1186),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4725_ (.D(net1188),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4726_ (.D(net1191),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4727_ (.D(net1192),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4728_ (.D(net1193),
    .GATE(net1081),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4729_ (.D(net162),
    .GATE(net1081),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4730_ (.D(net1196),
    .GATE(net1081),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4731_ (.D(net1197),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4732_ (.D(net1198),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4733_ (.D(net1199),
    .GATE(net1079),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4734_ (.D(net1200),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4735_ (.D(net1201),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4736_ (.D(net154),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4737_ (.D(net153),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4738_ (.D(net1205),
    .GATE(net1079),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4739_ (.D(net1206),
    .GATE(net1079),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4740_ (.D(net151),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4741_ (.D(net150),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4742_ (.D(net1210),
    .GATE(net1079),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4743_ (.D(net1211),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4744_ (.D(net1212),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4745_ (.D(net146),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4746_ (.D(net1179),
    .GATE(net1079),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4747_ (.D(net1180),
    .GATE(net1079),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4748_ (.D(net1181),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4749_ (.D(net1182),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4750_ (.D(net168),
    .GATE(net1081),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4751_ (.D(net167),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4752_ (.D(net166),
    .GATE(net1080),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4753_ (.D(net165),
    .GATE(net1078),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4754_ (.D(net1202),
    .GATE(net1079),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4755_ (.D(net1214),
    .GATE(net1079),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4756_ (.D(net1187),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4757_ (.D(net1189),
    .GATE(net1072),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4758_ (.D(net1191),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4759_ (.D(net1192),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4760_ (.D(net1194),
    .GATE(net1070),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4761_ (.D(net162),
    .GATE(net1070),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4762_ (.D(net1196),
    .GATE(net1070),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4763_ (.D(net160),
    .GATE(net1070),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4764_ (.D(net159),
    .GATE(net1070),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4765_ (.D(net1199),
    .GATE(net1070),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4766_ (.D(net1200),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4767_ (.D(net1201),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4768_ (.D(net1203),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4769_ (.D(net1204),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4770_ (.D(net1205),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4771_ (.D(net1206),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4772_ (.D(net1208),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4773_ (.D(net1209),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4774_ (.D(net1210),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4775_ (.D(net1211),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4776_ (.D(net1212),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4777_ (.D(net1213),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4778_ (.D(net1179),
    .GATE(net1070),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4779_ (.D(net1180),
    .GATE(net1070),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4780_ (.D(net170),
    .GATE(net1070),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4781_ (.D(net169),
    .GATE(net1072),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4782_ (.D(net168),
    .GATE(net1072),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4783_ (.D(net1184),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4784_ (.D(net1185),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4785_ (.D(net1190),
    .GATE(net1071),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4786_ (.D(net1202),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4787_ (.D(net1214),
    .GATE(net1069),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4788_ (.D(net1186),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4789_ (.D(net1188),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4790_ (.D(net1191),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4791_ (.D(net1192),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4792_ (.D(net1193),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4793_ (.D(net1195),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4794_ (.D(net1196),
    .GATE(net1164),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4795_ (.D(net1197),
    .GATE(net1164),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4796_ (.D(net1198),
    .GATE(net1164),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4797_ (.D(net158),
    .GATE(net1166),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4798_ (.D(net157),
    .GATE(net1164),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4799_ (.D(net156),
    .GATE(net1166),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4800_ (.D(net1203),
    .GATE(net1166),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4801_ (.D(net1204),
    .GATE(net1164),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4802_ (.D(net152),
    .GATE(net1164),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4803_ (.D(net1207),
    .GATE(net1164),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4804_ (.D(net151),
    .GATE(net1164),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4805_ (.D(net150),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4806_ (.D(net149),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4807_ (.D(net148),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4808_ (.D(net147),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4809_ (.D(net146),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4810_ (.D(net1179),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4811_ (.D(net1180),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4812_ (.D(net1181),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4813_ (.D(net1182),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4814_ (.D(net1183),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4815_ (.D(net1184),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4816_ (.D(net166),
    .GATE(net1164),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4817_ (.D(net1190),
    .GATE(net1163),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4818_ (.D(net1202),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4819_ (.D(net1214),
    .GATE(net1165),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4820_ (.D(net1186),
    .GATE(net1156),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4821_ (.D(net1188),
    .GATE(net1156),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4822_ (.D(net164),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4823_ (.D(net163),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4824_ (.D(net1194),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4825_ (.D(net162),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4826_ (.D(net161),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4827_ (.D(net1197),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4828_ (.D(net159),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4829_ (.D(net158),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4830_ (.D(net1200),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4831_ (.D(net1201),
    .GATE(net1156),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4832_ (.D(net1203),
    .GATE(net1156),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4833_ (.D(net153),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4834_ (.D(net152),
    .GATE(net1156),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4835_ (.D(net1206),
    .GATE(net1156),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4836_ (.D(net1208),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4837_ (.D(net1209),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4838_ (.D(net149),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4839_ (.D(net148),
    .GATE(net1157),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4840_ (.D(net147),
    .GATE(net1157),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4841_ (.D(net1213),
    .GATE(net1157),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4842_ (.D(net172),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4843_ (.D(net171),
    .GATE(net1155),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4844_ (.D(net170),
    .GATE(net1156),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4845_ (.D(net169),
    .GATE(net1156),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4846_ (.D(net168),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4847_ (.D(net167),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4848_ (.D(net166),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4849_ (.D(net1190),
    .GATE(net1154),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4850_ (.D(net1202),
    .GATE(net1157),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4851_ (.D(net1214),
    .GATE(net1156),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4852_ (.D(net1187),
    .GATE(net1148),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4853_ (.D(net1189),
    .GATE(net1148),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4854_ (.D(net1191),
    .GATE(net1148),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4855_ (.D(net1192),
    .GATE(net1148),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4856_ (.D(net1193),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4857_ (.D(net1195),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4858_ (.D(net1196),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4859_ (.D(net1197),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4860_ (.D(net1198),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4861_ (.D(net1199),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4862_ (.D(net1200),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4863_ (.D(net1201),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4864_ (.D(net1203),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4865_ (.D(net1204),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4866_ (.D(net1205),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4867_ (.D(net1206),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4868_ (.D(net1208),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4869_ (.D(net1209),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4870_ (.D(net1210),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4871_ (.D(net1211),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4872_ (.D(net1212),
    .GATE(net1153),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4873_ (.D(net1213),
    .GATE(net1153),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4874_ (.D(net1179),
    .GATE(net1148),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4875_ (.D(net1180),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4876_ (.D(net1181),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4877_ (.D(net1182),
    .GATE(net1147),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4878_ (.D(net1183),
    .GATE(net1149),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4879_ (.D(net1184),
    .GATE(net1149),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4880_ (.D(net1185),
    .GATE(net1149),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4881_ (.D(net165),
    .GATE(net1149),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4882_ (.D(net155),
    .GATE(net1146),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _4883_ (.D(net145),
    .GATE(net1149),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ));
 sky130_fd_sc_hd__buf_1 _4884_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ),
    .X(net235));
 sky130_fd_sc_hd__buf_6 _4885_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ),
    .X(net236));
 sky130_fd_sc_hd__buf_1 _4886_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ),
    .X(net237));
 sky130_fd_sc_hd__buf_1 _4887_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ),
    .X(net238));
 sky130_fd_sc_hd__buf_2 _4888_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 _4889_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 _4890_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ),
    .X(net241));
 sky130_fd_sc_hd__buf_4 _4891_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .X(net242));
 sky130_fd_sc_hd__buf_1 _4892_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .X(net243));
 sky130_fd_sc_hd__buf_4 _4893_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .X(net244));
 sky130_fd_sc_hd__buf_1 _4894_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .X(net245));
 sky130_fd_sc_hd__buf_1 _4895_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 _4896_ (.A(net13),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 _4897_ (.A(net14),
    .X(net248));
 sky130_fd_sc_hd__buf_1 _4898_ (.A(net15),
    .X(net249));
 sky130_fd_sc_hd__buf_1 _4899_ (.A(net16),
    .X(net250));
 sky130_fd_sc_hd__buf_1 _4900_ (.A(net17),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 _4901_ (.A(net18),
    .X(net252));
 sky130_fd_sc_hd__buf_1 _4902_ (.A(net19),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 _4903_ (.A(net20),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 _4904_ (.A(Tile_X0Y0_E6END[2]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 _4905_ (.A(Tile_X0Y0_E6END[3]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 _4906_ (.A(Tile_X0Y0_E6END[4]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 _4907_ (.A(Tile_X0Y0_E6END[5]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 _4908_ (.A(Tile_X0Y0_E6END[6]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 _4909_ (.A(Tile_X0Y0_E6END[7]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 _4910_ (.A(Tile_X0Y0_E6END[8]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 _4911_ (.A(Tile_X0Y0_E6END[9]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 _4912_ (.A(Tile_X0Y0_E6END[10]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 _4913_ (.A(Tile_X0Y0_E6END[11]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 _4914_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 _4915_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ),
    .X(net257));
 sky130_fd_sc_hd__buf_1 _4916_ (.A(Tile_X0Y0_EE4END[4]),
    .X(net267));
 sky130_fd_sc_hd__buf_1 _4917_ (.A(Tile_X0Y0_EE4END[5]),
    .X(net274));
 sky130_fd_sc_hd__buf_1 _4918_ (.A(Tile_X0Y0_EE4END[6]),
    .X(net275));
 sky130_fd_sc_hd__buf_1 _4919_ (.A(Tile_X0Y0_EE4END[7]),
    .X(net276));
 sky130_fd_sc_hd__buf_1 _4920_ (.A(Tile_X0Y0_EE4END[8]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 _4921_ (.A(Tile_X0Y0_EE4END[9]),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 _4922_ (.A(Tile_X0Y0_EE4END[10]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 _4923_ (.A(Tile_X0Y0_EE4END[11]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 _4924_ (.A(Tile_X0Y0_EE4END[12]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 _4925_ (.A(Tile_X0Y0_EE4END[13]),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 _4926_ (.A(Tile_X0Y0_EE4END[14]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 _4927_ (.A(Tile_X0Y0_EE4END[15]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 _4928_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 _4929_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ),
    .X(net271));
 sky130_fd_sc_hd__buf_1 _4930_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 _4931_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ),
    .X(net273));
 sky130_fd_sc_hd__buf_4 _4932_ (.A(net1254),
    .X(net283));
 sky130_fd_sc_hd__buf_4 _4933_ (.A(net1243),
    .X(net294));
 sky130_fd_sc_hd__buf_1 _4934_ (.A(net47),
    .X(net305));
 sky130_fd_sc_hd__buf_1 _4935_ (.A(net50),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 _4936_ (.A(net51),
    .X(net309));
 sky130_fd_sc_hd__buf_2 _4937_ (.A(net1225),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_2 _4938_ (.A(net53),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_2 _4939_ (.A(net54),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 _4940_ (.A(net1222),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 _4941_ (.A(net1221),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_2 _4942_ (.A(net1253),
    .X(net284));
 sky130_fd_sc_hd__buf_2 _4943_ (.A(net1252),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 _4944_ (.A(net30),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 _4945_ (.A(net31),
    .X(net287));
 sky130_fd_sc_hd__buf_2 _4946_ (.A(net32),
    .X(net288));
 sky130_fd_sc_hd__buf_2 _4947_ (.A(net33),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 _4948_ (.A(net1247),
    .X(net290));
 sky130_fd_sc_hd__buf_1 _4949_ (.A(net1246),
    .X(net291));
 sky130_fd_sc_hd__buf_1 _4950_ (.A(net36),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_1 _4951_ (.A(net1244),
    .X(net293));
 sky130_fd_sc_hd__buf_1 _4952_ (.A(net39),
    .X(net295));
 sky130_fd_sc_hd__buf_1 _4953_ (.A(net40),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 _4954_ (.A(net1240),
    .X(net297));
 sky130_fd_sc_hd__buf_1 _4955_ (.A(net42),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 _4956_ (.A(net1238),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_2 _4957_ (.A(net1237),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 _4958_ (.A(net1235),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_2 _4959_ (.A(net1233),
    .X(net302));
 sky130_fd_sc_hd__buf_1 _4960_ (.A(net45),
    .X(net303));
 sky130_fd_sc_hd__buf_1 _4961_ (.A(net1231),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 _4962_ (.A(net1229),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 _4963_ (.A(net1228),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 _4964_ (.A(net1176),
    .X(net315));
 sky130_fd_sc_hd__buf_1 _4965_ (.A(net1143),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 _4966_ (.A(net1135),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 _4967_ (.A(net1126),
    .X(net328));
 sky130_fd_sc_hd__buf_1 _4968_ (.A(net1117),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 _4969_ (.A(net1109),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 _4970_ (.A(net1100),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_2 _4971_ (.A(net1091),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 _4972_ (.A(net1084),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_2 _4973_ (.A(net1077),
    .X(net334));
 sky130_fd_sc_hd__buf_1 _4974_ (.A(net1169),
    .X(net316));
 sky130_fd_sc_hd__buf_1 _4975_ (.A(net1160),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 _4976_ (.A(net1151),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 _4977_ (.A(Tile_X0Y1_FrameStrobe[13]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 _4978_ (.A(Tile_X0Y1_FrameStrobe[14]),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 _4979_ (.A(Tile_X0Y1_FrameStrobe[15]),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 _4980_ (.A(Tile_X0Y1_FrameStrobe[16]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 _4981_ (.A(Tile_X0Y1_FrameStrobe[17]),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 _4982_ (.A(Tile_X0Y1_FrameStrobe[18]),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 _4983_ (.A(Tile_X0Y1_FrameStrobe[19]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 _4984_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ),
    .X(net335));
 sky130_fd_sc_hd__buf_6 clone133 (.A(net1025),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_2 _4986_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 _4987_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ),
    .X(net338));
 sky130_fd_sc_hd__buf_1 _4988_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_2 _4989_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 _4990_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .X(net341));
 sky130_fd_sc_hd__buf_4 _4991_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 _4992_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 _4993_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ),
    .X(net344));
 sky130_fd_sc_hd__buf_1 _4994_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_2 _4995_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ),
    .X(net346));
 sky130_fd_sc_hd__buf_6 _4996_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .X(net347));
 sky130_fd_sc_hd__buf_6 _4997_ (.A(net666),
    .X(net348));
 sky130_fd_sc_hd__buf_6 _4998_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .X(net349));
 sky130_fd_sc_hd__buf_6 _4999_ (.A(net694),
    .X(net350));
 sky130_fd_sc_hd__buf_4 _5000_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .X(net351));
 sky130_fd_sc_hd__buf_4 _5001_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .X(net352));
 sky130_fd_sc_hd__buf_2 _5002_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .X(net353));
 sky130_fd_sc_hd__buf_4 _5003_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_1 _5004_ (.A(Tile_X0Y1_N4END[8]),
    .X(net355));
 sky130_fd_sc_hd__buf_1 _5005_ (.A(Tile_X0Y1_N4END[9]),
    .X(net362));
 sky130_fd_sc_hd__buf_1 _5006_ (.A(Tile_X0Y1_N4END[10]),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 _5007_ (.A(Tile_X0Y1_N4END[11]),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 _5008_ (.A(Tile_X0Y1_N4END[12]),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 _5009_ (.A(Tile_X0Y1_N4END[13]),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_1 _5010_ (.A(Tile_X0Y1_N4END[14]),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 _5011_ (.A(Tile_X0Y1_N4END[15]),
    .X(net368));
 sky130_fd_sc_hd__buf_6 _5012_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ),
    .X(net369));
 sky130_fd_sc_hd__buf_4 _5013_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ),
    .X(net370));
 sky130_fd_sc_hd__buf_4 _5014_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ),
    .X(net356));
 sky130_fd_sc_hd__buf_6 _5015_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ),
    .X(net357));
 sky130_fd_sc_hd__buf_1 _5016_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ),
    .X(net358));
 sky130_fd_sc_hd__buf_1 _5017_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ),
    .X(net359));
 sky130_fd_sc_hd__buf_1 _5018_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 _5019_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ),
    .X(net361));
 sky130_fd_sc_hd__buf_1 _5020_ (.A(Tile_X0Y1_NN4END[8]),
    .X(net371));
 sky130_fd_sc_hd__buf_1 _5021_ (.A(Tile_X0Y1_NN4END[9]),
    .X(net378));
 sky130_fd_sc_hd__buf_1 _5022_ (.A(Tile_X0Y1_NN4END[10]),
    .X(net379));
 sky130_fd_sc_hd__buf_1 _5023_ (.A(Tile_X0Y1_NN4END[11]),
    .X(net380));
 sky130_fd_sc_hd__buf_1 _5024_ (.A(Tile_X0Y1_NN4END[12]),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 _5025_ (.A(Tile_X0Y1_NN4END[13]),
    .X(net382));
 sky130_fd_sc_hd__buf_1 _5026_ (.A(Tile_X0Y1_NN4END[14]),
    .X(net383));
 sky130_fd_sc_hd__buf_1 _5027_ (.A(Tile_X0Y1_NN4END[15]),
    .X(net384));
 sky130_fd_sc_hd__buf_6 _5028_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ),
    .X(net385));
 sky130_fd_sc_hd__buf_6 _5029_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ),
    .X(net386));
 sky130_fd_sc_hd__buf_4 _5030_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ),
    .X(net372));
 sky130_fd_sc_hd__buf_4 _5031_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ),
    .X(net373));
 sky130_fd_sc_hd__buf_1 _5032_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 _5033_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ),
    .X(net375));
 sky130_fd_sc_hd__buf_1 _5034_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ),
    .X(net376));
 sky130_fd_sc_hd__buf_4 _5035_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ),
    .X(net377));
 sky130_fd_sc_hd__buf_2 _5036_ (.A(clknet_1_0__leaf_Tile_X0Y1_UserCLK),
    .X(net387));
 sky130_fd_sc_hd__buf_1 _5037_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 _5038_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 _5039_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ),
    .X(net390));
 sky130_fd_sc_hd__buf_1 _5040_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ),
    .X(net391));
 sky130_fd_sc_hd__buf_1 _5041_ (.A(net97),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 _5042_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .X(net393));
 sky130_fd_sc_hd__buf_1 _5043_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .X(net394));
 sky130_fd_sc_hd__buf_1 _5044_ (.A(net100),
    .X(net395));
 sky130_fd_sc_hd__buf_1 _5045_ (.A(net101),
    .X(net396));
 sky130_fd_sc_hd__buf_4 _5046_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ),
    .X(net397));
 sky130_fd_sc_hd__buf_4 _5047_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .X(net398));
 sky130_fd_sc_hd__buf_1 _5048_ (.A(net104),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_2 _5049_ (.A(net105),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 _5050_ (.A(net106),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_2 _5051_ (.A(net107),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 _5052_ (.A(net108),
    .X(net403));
 sky130_fd_sc_hd__buf_1 _5053_ (.A(net109),
    .X(net404));
 sky130_fd_sc_hd__buf_1 _5054_ (.A(net110),
    .X(net405));
 sky130_fd_sc_hd__buf_1 _5055_ (.A(net111),
    .X(net406));
 sky130_fd_sc_hd__buf_1 _5056_ (.A(net112),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 _5057_ (.A(Tile_X0Y0_W6END[2]),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_2 _5058_ (.A(Tile_X0Y0_W6END[3]),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 _5059_ (.A(Tile_X0Y0_W6END[4]),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_2 _5060_ (.A(Tile_X0Y0_W6END[5]),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_2 _5061_ (.A(Tile_X0Y0_W6END[6]),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_2 _5062_ (.A(Tile_X0Y0_W6END[7]),
    .X(net415));
 sky130_fd_sc_hd__buf_4 _5063_ (.A(Tile_X0Y0_W6END[8]),
    .X(net416));
 sky130_fd_sc_hd__buf_4 _5064_ (.A(Tile_X0Y0_W6END[9]),
    .X(net417));
 sky130_fd_sc_hd__buf_2 _5065_ (.A(Tile_X0Y0_W6END[10]),
    .X(net418));
 sky130_fd_sc_hd__buf_4 _5066_ (.A(Tile_X0Y0_W6END[11]),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_2 _5067_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ),
    .X(net409));
 sky130_fd_sc_hd__buf_4 _5068_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_2 _5069_ (.A(Tile_X0Y0_WW4END[4]),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 _5070_ (.A(Tile_X0Y0_WW4END[5]),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 _5071_ (.A(Tile_X0Y0_WW4END[6]),
    .X(net428));
 sky130_fd_sc_hd__buf_2 _5072_ (.A(Tile_X0Y0_WW4END[7]),
    .X(net429));
 sky130_fd_sc_hd__buf_2 _5073_ (.A(Tile_X0Y0_WW4END[8]),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 _5074_ (.A(Tile_X0Y0_WW4END[9]),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_2 _5075_ (.A(Tile_X0Y0_WW4END[10]),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_2 _5076_ (.A(Tile_X0Y0_WW4END[11]),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_2 _5077_ (.A(Tile_X0Y0_WW4END[12]),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_2 _5078_ (.A(Tile_X0Y0_WW4END[13]),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 _5079_ (.A(Tile_X0Y0_WW4END[14]),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_2 _5080_ (.A(Tile_X0Y0_WW4END[15]),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_2 _5081_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ),
    .X(net423));
 sky130_fd_sc_hd__buf_4 _5082_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_1 _5083_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ),
    .X(net425));
 sky130_fd_sc_hd__buf_2 _5084_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ),
    .X(net426));
 sky130_fd_sc_hd__buf_1 _5085_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ),
    .X(net436));
 sky130_fd_sc_hd__buf_1 _5086_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_1 _5087_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ),
    .X(net438));
 sky130_fd_sc_hd__buf_1 _5088_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_2 _5089_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ),
    .X(net440));
 sky130_fd_sc_hd__buf_1 _5090_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_2 _5091_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 _5092_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .X(net443));
 sky130_fd_sc_hd__buf_1 _5093_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_2 _5094_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .X(net445));
 sky130_fd_sc_hd__buf_6 _5095_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .X(net446));
 sky130_fd_sc_hd__buf_6 _5096_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_2 _5097_ (.A(net131),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_2 _5098_ (.A(net132),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 _5099_ (.A(net133),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 _5100_ (.A(net134),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 _5101_ (.A(net135),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 _5102_ (.A(net136),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_2 _5103_ (.A(net137),
    .X(net454));
 sky130_fd_sc_hd__buf_1 _5104_ (.A(net138),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 _5105_ (.A(Tile_X0Y1_E6END[2]),
    .X(net456));
 sky130_fd_sc_hd__buf_1 _5106_ (.A(Tile_X0Y1_E6END[3]),
    .X(net459));
 sky130_fd_sc_hd__buf_1 _5107_ (.A(Tile_X0Y1_E6END[4]),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_2 _5108_ (.A(Tile_X0Y1_E6END[5]),
    .X(net461));
 sky130_fd_sc_hd__buf_1 _5109_ (.A(Tile_X0Y1_E6END[6]),
    .X(net462));
 sky130_fd_sc_hd__buf_1 _5110_ (.A(Tile_X0Y1_E6END[7]),
    .X(net463));
 sky130_fd_sc_hd__buf_1 _5111_ (.A(Tile_X0Y1_E6END[8]),
    .X(net464));
 sky130_fd_sc_hd__buf_1 _5112_ (.A(Tile_X0Y1_E6END[9]),
    .X(net465));
 sky130_fd_sc_hd__buf_1 _5113_ (.A(Tile_X0Y1_E6END[10]),
    .X(net466));
 sky130_fd_sc_hd__buf_1 _5114_ (.A(Tile_X0Y1_E6END[11]),
    .X(net467));
 sky130_fd_sc_hd__buf_1 _5115_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ),
    .X(net457));
 sky130_fd_sc_hd__buf_6 _5116_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 _5117_ (.A(Tile_X0Y1_EE4END[4]),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_1 _5118_ (.A(Tile_X0Y1_EE4END[5]),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_1 _5119_ (.A(Tile_X0Y1_EE4END[6]),
    .X(net476));
 sky130_fd_sc_hd__buf_1 _5120_ (.A(Tile_X0Y1_EE4END[7]),
    .X(net477));
 sky130_fd_sc_hd__buf_1 _5121_ (.A(Tile_X0Y1_EE4END[8]),
    .X(net478));
 sky130_fd_sc_hd__buf_1 _5122_ (.A(Tile_X0Y1_EE4END[9]),
    .X(net479));
 sky130_fd_sc_hd__buf_1 _5123_ (.A(Tile_X0Y1_EE4END[10]),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 _5124_ (.A(Tile_X0Y1_EE4END[11]),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 _5125_ (.A(Tile_X0Y1_EE4END[12]),
    .X(net482));
 sky130_fd_sc_hd__buf_1 _5126_ (.A(Tile_X0Y1_EE4END[13]),
    .X(net483));
 sky130_fd_sc_hd__buf_1 _5127_ (.A(Tile_X0Y1_EE4END[14]),
    .X(net469));
 sky130_fd_sc_hd__buf_1 _5128_ (.A(Tile_X0Y1_EE4END[15]),
    .X(net470));
 sky130_fd_sc_hd__buf_1 _5129_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ),
    .X(net471));
 sky130_fd_sc_hd__buf_2 _5130_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ),
    .X(net472));
 sky130_fd_sc_hd__buf_6 _5131_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ),
    .X(net473));
 sky130_fd_sc_hd__buf_6 clone90 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .X(net707));
 sky130_fd_sc_hd__buf_1 _5133_ (.A(net145),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_1 _5134_ (.A(net155),
    .X(net495));
 sky130_fd_sc_hd__buf_1 _5135_ (.A(net165),
    .X(net506));
 sky130_fd_sc_hd__buf_2 _5136_ (.A(net1185),
    .X(net509));
 sky130_fd_sc_hd__buf_4 _5137_ (.A(net1184),
    .X(net510));
 sky130_fd_sc_hd__buf_2 _5138_ (.A(net1183),
    .X(net511));
 sky130_fd_sc_hd__buf_4 _5139_ (.A(net1182),
    .X(net512));
 sky130_fd_sc_hd__buf_4 _5140_ (.A(net1181),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_2 _5141_ (.A(net1180),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_2 _5142_ (.A(net1179),
    .X(net515));
 sky130_fd_sc_hd__buf_2 _5143_ (.A(net1213),
    .X(net485));
 sky130_fd_sc_hd__buf_4 _5144_ (.A(net1212),
    .X(net486));
 sky130_fd_sc_hd__buf_4 _5145_ (.A(net1211),
    .X(net487));
 sky130_fd_sc_hd__buf_1 _5146_ (.A(net149),
    .X(net488));
 sky130_fd_sc_hd__buf_1 _5147_ (.A(net150),
    .X(net489));
 sky130_fd_sc_hd__buf_1 _5148_ (.A(net151),
    .X(net490));
 sky130_fd_sc_hd__buf_1 _5149_ (.A(net1206),
    .X(net491));
 sky130_fd_sc_hd__buf_1 _5150_ (.A(net1205),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_2 _5151_ (.A(net1204),
    .X(net493));
 sky130_fd_sc_hd__buf_1 _5152_ (.A(net154),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_2 _5153_ (.A(net1201),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_2 _5154_ (.A(net1200),
    .X(net497));
 sky130_fd_sc_hd__buf_1 _5155_ (.A(net158),
    .X(net498));
 sky130_fd_sc_hd__buf_1 _5156_ (.A(net159),
    .X(net499));
 sky130_fd_sc_hd__buf_1 _5157_ (.A(net160),
    .X(net500));
 sky130_fd_sc_hd__buf_1 _5158_ (.A(net161),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_2 _5159_ (.A(net162),
    .X(net502));
 sky130_fd_sc_hd__buf_2 _5160_ (.A(net1194),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_2 _5161_ (.A(net163),
    .X(net504));
 sky130_fd_sc_hd__buf_1 _5162_ (.A(net164),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_2 _5163_ (.A(net1189),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_2 _5164_ (.A(net1187),
    .X(net508));
 sky130_fd_sc_hd__buf_1 _5165_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_1 _5166_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ),
    .X(net517));
 sky130_fd_sc_hd__buf_1 _5167_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ),
    .X(net518));
 sky130_fd_sc_hd__buf_1 _5168_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_1 _5169_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_1 _5170_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .X(net521));
 sky130_fd_sc_hd__buf_1 _5171_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .X(net522));
 sky130_fd_sc_hd__buf_1 _5172_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .X(net523));
 sky130_fd_sc_hd__buf_6 _5173_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .X(net524));
 sky130_fd_sc_hd__buf_4 _5174_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_2 _5175_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .X(net526));
 sky130_fd_sc_hd__buf_6 _5176_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ),
    .X(net527));
 sky130_fd_sc_hd__buf_4 _5177_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .X(net528));
 sky130_fd_sc_hd__buf_4 _5178_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .X(net529));
 sky130_fd_sc_hd__buf_2 _5179_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .X(net530));
 sky130_fd_sc_hd__buf_4 _5180_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .X(net531));
 sky130_fd_sc_hd__buf_2 _5181_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .X(net532));
 sky130_fd_sc_hd__buf_4 _5182_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .X(net533));
 sky130_fd_sc_hd__buf_4 _5183_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_2 _5184_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .X(net535));
 sky130_fd_sc_hd__buf_6 _5185_ (.A(Tile_X0Y0_S4END[8]),
    .X(net536));
 sky130_fd_sc_hd__buf_6 _5186_ (.A(Tile_X0Y0_S4END[9]),
    .X(net543));
 sky130_fd_sc_hd__buf_6 _5187_ (.A(Tile_X0Y0_S4END[10]),
    .X(net544));
 sky130_fd_sc_hd__buf_6 _5188_ (.A(Tile_X0Y0_S4END[11]),
    .X(net545));
 sky130_fd_sc_hd__buf_6 _5189_ (.A(Tile_X0Y0_S4END[12]),
    .X(net546));
 sky130_fd_sc_hd__buf_6 _5190_ (.A(Tile_X0Y0_S4END[13]),
    .X(net547));
 sky130_fd_sc_hd__buf_6 _5191_ (.A(Tile_X0Y0_S4END[14]),
    .X(net548));
 sky130_fd_sc_hd__buf_6 _5192_ (.A(Tile_X0Y0_S4END[15]),
    .X(net549));
 sky130_fd_sc_hd__buf_4 _5193_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ),
    .X(net550));
 sky130_fd_sc_hd__buf_4 _5194_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ),
    .X(net551));
 sky130_fd_sc_hd__buf_4 _5195_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ),
    .X(net537));
 sky130_fd_sc_hd__buf_6 _5196_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_1 _5197_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_1 _5198_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ),
    .X(net540));
 sky130_fd_sc_hd__buf_1 _5199_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ),
    .X(net541));
 sky130_fd_sc_hd__buf_1 _5200_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ),
    .X(net542));
 sky130_fd_sc_hd__buf_6 _5201_ (.A(Tile_X0Y0_SS4END[8]),
    .X(net552));
 sky130_fd_sc_hd__buf_6 _5202_ (.A(Tile_X0Y0_SS4END[9]),
    .X(net559));
 sky130_fd_sc_hd__buf_6 _5203_ (.A(Tile_X0Y0_SS4END[10]),
    .X(net560));
 sky130_fd_sc_hd__buf_6 _5204_ (.A(Tile_X0Y0_SS4END[11]),
    .X(net561));
 sky130_fd_sc_hd__buf_6 _5205_ (.A(Tile_X0Y0_SS4END[12]),
    .X(net562));
 sky130_fd_sc_hd__buf_6 _5206_ (.A(Tile_X0Y0_SS4END[13]),
    .X(net563));
 sky130_fd_sc_hd__buf_6 _5207_ (.A(Tile_X0Y0_SS4END[14]),
    .X(net564));
 sky130_fd_sc_hd__buf_6 _5208_ (.A(Tile_X0Y0_SS4END[15]),
    .X(net565));
 sky130_fd_sc_hd__buf_6 _5209_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ),
    .X(net566));
 sky130_fd_sc_hd__buf_6 _5210_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ),
    .X(net567));
 sky130_fd_sc_hd__buf_4 _5211_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ),
    .X(net553));
 sky130_fd_sc_hd__buf_6 _5212_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_1 _5213_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ),
    .X(net555));
 sky130_fd_sc_hd__buf_4 _5214_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ),
    .X(net556));
 sky130_fd_sc_hd__buf_1 _5215_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_2 _5216_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ),
    .X(net558));
 sky130_fd_sc_hd__buf_1 _5217_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ),
    .X(net568));
 sky130_fd_sc_hd__buf_1 _5218_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ),
    .X(net569));
 sky130_fd_sc_hd__buf_1 _5219_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ),
    .X(net570));
 sky130_fd_sc_hd__buf_1 _5220_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ),
    .X(net571));
 sky130_fd_sc_hd__buf_1 _5221_ (.A(net213),
    .X(net572));
 sky130_fd_sc_hd__buf_1 _5222_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .X(net573));
 sky130_fd_sc_hd__buf_1 _5223_ (.A(net705),
    .X(net574));
 sky130_fd_sc_hd__buf_1 _5224_ (.A(net216),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_1 _5225_ (.A(net217),
    .X(net576));
 sky130_fd_sc_hd__buf_4 _5226_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .X(net577));
 sky130_fd_sc_hd__buf_6 clone106 (.A(net1053),
    .X(net723));
 sky130_fd_sc_hd__buf_1 _5228_ (.A(net220),
    .X(net579));
 sky130_fd_sc_hd__buf_1 _5229_ (.A(net221),
    .X(net580));
 sky130_fd_sc_hd__buf_1 _5230_ (.A(net222),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 _5231_ (.A(net223),
    .X(net582));
 sky130_fd_sc_hd__buf_1 _5232_ (.A(net224),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_2 _5233_ (.A(net225),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_2 _5234_ (.A(net226),
    .X(net585));
 sky130_fd_sc_hd__buf_4 _5235_ (.A(net227),
    .X(net586));
 sky130_fd_sc_hd__buf_4 _5236_ (.A(net228),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_2 _5237_ (.A(Tile_X0Y1_W6END[2]),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_2 _5238_ (.A(Tile_X0Y1_W6END[3]),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_2 _5239_ (.A(Tile_X0Y1_W6END[4]),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_2 _5240_ (.A(Tile_X0Y1_W6END[5]),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_2 _5241_ (.A(Tile_X0Y1_W6END[6]),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_2 _5242_ (.A(Tile_X0Y1_W6END[7]),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_2 _5243_ (.A(Tile_X0Y1_W6END[8]),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_2 _5244_ (.A(Tile_X0Y1_W6END[9]),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_2 _5245_ (.A(Tile_X0Y1_W6END[10]),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_2 _5246_ (.A(Tile_X0Y1_W6END[11]),
    .X(net599));
 sky130_fd_sc_hd__buf_1 _5247_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_1 clone74 (.A(net704),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_2 _5249_ (.A(Tile_X0Y1_WW4END[4]),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_2 _5250_ (.A(Tile_X0Y1_WW4END[5]),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_2 _5251_ (.A(Tile_X0Y1_WW4END[6]),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_2 _5252_ (.A(Tile_X0Y1_WW4END[7]),
    .X(net609));
 sky130_fd_sc_hd__buf_2 _5253_ (.A(Tile_X0Y1_WW4END[8]),
    .X(net610));
 sky130_fd_sc_hd__buf_2 _5254_ (.A(Tile_X0Y1_WW4END[9]),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_2 _5255_ (.A(Tile_X0Y1_WW4END[10]),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_2 _5256_ (.A(Tile_X0Y1_WW4END[11]),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_2 _5257_ (.A(Tile_X0Y1_WW4END[12]),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_2 _5258_ (.A(Tile_X0Y1_WW4END[13]),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_2 _5259_ (.A(Tile_X0Y1_WW4END[14]),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_2 _5260_ (.A(Tile_X0Y1_WW4END[15]),
    .X(net602));
 sky130_fd_sc_hd__buf_1 _5261_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ),
    .X(net603));
 sky130_fd_sc_hd__o21ai_4 clone48 (.A1(net1061),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .B1(_0708_),
    .Y(net665));
 sky130_fd_sc_hd__clkbuf_1 _5263_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_2 rebuffer96 (.A(net1049),
    .X(net713));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1660 ();
 sky130_fd_sc_hd__buf_2 fanout963 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_4 fanout964 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .X(net964));
 sky130_fd_sc_hd__buf_6 fanout965 (.A(_0299_),
    .X(net965));
 sky130_fd_sc_hd__buf_8 fanout966 (.A(net731),
    .X(net966));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout967 (.A(net732),
    .X(net967));
 sky130_fd_sc_hd__buf_8 fanout968 (.A(net969),
    .X(net968));
 sky130_fd_sc_hd__buf_6 fanout969 (.A(net970),
    .X(net969));
 sky130_fd_sc_hd__buf_6 fanout970 (.A(net726),
    .X(net970));
 sky130_fd_sc_hd__buf_4 fanout971 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .X(net971));
 sky130_fd_sc_hd__clkbuf_2 fanout972 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .X(net972));
 sky130_fd_sc_hd__buf_2 fanout973 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__buf_2 fanout974 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .X(net974));
 sky130_fd_sc_hd__buf_8 fanout975 (.A(net977),
    .X(net975));
 sky130_fd_sc_hd__buf_2 fanout976 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__buf_8 fanout977 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .X(net977));
 sky130_fd_sc_hd__buf_2 fanout978 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_4 fanout979 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .X(net979));
 sky130_fd_sc_hd__buf_12 fanout980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__buf_8 fanout981 (.A(net982),
    .X(net981));
 sky130_fd_sc_hd__buf_8 fanout982 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .X(net982));
 sky130_fd_sc_hd__buf_2 fanout983 (.A(net984),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_4 fanout984 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .X(net984));
 sky130_fd_sc_hd__buf_8 fanout985 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .X(net985));
 sky130_fd_sc_hd__buf_6 fanout986 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .X(net986));
 sky130_fd_sc_hd__buf_2 fanout987 (.A(net988),
    .X(net987));
 sky130_fd_sc_hd__buf_2 fanout988 (.A(net989),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_2 fanout989 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .X(net989));
 sky130_fd_sc_hd__buf_2 fanout990 (.A(net991),
    .X(net990));
 sky130_fd_sc_hd__buf_8 fanout991 (.A(net994),
    .X(net991));
 sky130_fd_sc_hd__buf_2 fanout992 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_2 fanout993 (.A(net994),
    .X(net993));
 sky130_fd_sc_hd__buf_12 fanout994 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .X(net994));
 sky130_fd_sc_hd__buf_2 fanout995 (.A(net999),
    .X(net995));
 sky130_fd_sc_hd__buf_8 fanout996 (.A(net999),
    .X(net996));
 sky130_fd_sc_hd__buf_2 fanout997 (.A(net998),
    .X(net997));
 sky130_fd_sc_hd__buf_2 fanout998 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__buf_8 fanout999 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .X(net999));
 sky130_fd_sc_hd__buf_8 fanout1000 (.A(net1001),
    .X(net1000));
 sky130_fd_sc_hd__buf_12 fanout1001 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_2 fanout1002 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_4 fanout1003 (.A(_1361_),
    .X(net1003));
 sky130_fd_sc_hd__buf_8 fanout1004 (.A(net1005),
    .X(net1004));
 sky130_fd_sc_hd__buf_8 fanout1005 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .X(net1005));
 sky130_fd_sc_hd__buf_6 fanout1006 (.A(net1007),
    .X(net1006));
 sky130_fd_sc_hd__buf_8 fanout1007 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_2 fanout1008 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .X(net1008));
 sky130_fd_sc_hd__buf_8 fanout1009 (.A(net1010),
    .X(net1009));
 sky130_fd_sc_hd__buf_8 fanout1010 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_4 fanout1011 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .X(net1011));
 sky130_fd_sc_hd__buf_2 fanout1012 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .X(net1012));
 sky130_fd_sc_hd__buf_8 fanout1013 (.A(net1015),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout1014 (.A(net1015),
    .X(net1014));
 sky130_fd_sc_hd__buf_12 fanout1015 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .X(net1015));
 sky130_fd_sc_hd__buf_6 fanout1016 (.A(net1017),
    .X(net1016));
 sky130_fd_sc_hd__buf_4 fanout1017 (.A(net1020),
    .X(net1017));
 sky130_fd_sc_hd__buf_8 fanout1018 (.A(net1020),
    .X(net1018));
 sky130_fd_sc_hd__buf_2 fanout1019 (.A(net1020),
    .X(net1019));
 sky130_fd_sc_hd__buf_12 fanout1020 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_4 fanout1021 (.A(net1023),
    .X(net1021));
 sky130_fd_sc_hd__buf_8 fanout1022 (.A(net676),
    .X(net1022));
 sky130_fd_sc_hd__buf_8 fanout1023 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .X(net1023));
 sky130_fd_sc_hd__buf_8 fanout1024 (.A(net1025),
    .X(net1024));
 sky130_fd_sc_hd__buf_8 fanout1025 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .X(net1025));
 sky130_fd_sc_hd__buf_2 fanout1026 (.A(net1028),
    .X(net1026));
 sky130_fd_sc_hd__buf_2 fanout1027 (.A(net1028),
    .X(net1027));
 sky130_fd_sc_hd__buf_2 fanout1028 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .X(net1028));
 sky130_fd_sc_hd__buf_8 fanout1029 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .X(net1029));
 sky130_fd_sc_hd__buf_2 fanout1030 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .X(net1030));
 sky130_fd_sc_hd__buf_2 fanout1031 (.A(net1033),
    .X(net1031));
 sky130_fd_sc_hd__buf_2 fanout1032 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__buf_2 fanout1033 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .X(net1033));
 sky130_fd_sc_hd__buf_8 fanout1034 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__buf_8 fanout1035 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .X(net1035));
 sky130_fd_sc_hd__clkbuf_4 fanout1036 (.A(net1038),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_2 fanout1037 (.A(net1038),
    .X(net1037));
 sky130_fd_sc_hd__buf_2 fanout1038 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .X(net1038));
 sky130_fd_sc_hd__buf_2 fanout1039 (.A(net1041),
    .X(net1039));
 sky130_fd_sc_hd__buf_6 fanout1040 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__buf_8 fanout1041 (.A(net1044),
    .X(net1041));
 sky130_fd_sc_hd__buf_2 fanout1042 (.A(net1044),
    .X(net1042));
 sky130_fd_sc_hd__buf_2 fanout1043 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__buf_8 fanout1044 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .X(net1044));
 sky130_fd_sc_hd__buf_8 fanout1045 (.A(net1048),
    .X(net1045));
 sky130_fd_sc_hd__clkbuf_4 fanout1046 (.A(net1047),
    .X(net1046));
 sky130_fd_sc_hd__buf_2 fanout1047 (.A(net1048),
    .X(net1047));
 sky130_fd_sc_hd__buf_12 fanout1048 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .X(net1048));
 sky130_fd_sc_hd__buf_8 fanout1049 (.A(net1053),
    .X(net1049));
 sky130_fd_sc_hd__buf_2 fanout1050 (.A(net1052),
    .X(net1050));
 sky130_fd_sc_hd__buf_2 fanout1051 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__buf_2 fanout1052 (.A(net1053),
    .X(net1052));
 sky130_fd_sc_hd__buf_8 fanout1053 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_4 fanout1054 (.A(net1056),
    .X(net1054));
 sky130_fd_sc_hd__buf_2 fanout1055 (.A(net1056),
    .X(net1055));
 sky130_fd_sc_hd__buf_8 fanout1056 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .X(net1056));
 sky130_fd_sc_hd__clkbuf_4 fanout1057 (.A(_0099_),
    .X(net1057));
 sky130_fd_sc_hd__buf_4 fanout1058 (.A(_0099_),
    .X(net1058));
 sky130_fd_sc_hd__clkbuf_8 fanout1059 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .X(net1059));
 sky130_fd_sc_hd__buf_2 fanout1060 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .X(net1060));
 sky130_fd_sc_hd__buf_4 fanout1061 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .X(net1061));
 sky130_fd_sc_hd__clkbuf_4 fanout1062 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_4 fanout1063 (.A(net1064),
    .X(net1063));
 sky130_fd_sc_hd__buf_4 fanout1064 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .X(net1064));
 sky130_fd_sc_hd__clkbuf_4 fanout1065 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .X(net1065));
 sky130_fd_sc_hd__clkbuf_4 fanout1066 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_4 fanout1067 (.A(net212),
    .X(net1067));
 sky130_fd_sc_hd__buf_4 fanout1068 (.A(net211),
    .X(net1068));
 sky130_fd_sc_hd__buf_2 fanout1069 (.A(net1070),
    .X(net1069));
 sky130_fd_sc_hd__clkbuf_4 fanout1070 (.A(net1072),
    .X(net1070));
 sky130_fd_sc_hd__buf_2 fanout1071 (.A(net1072),
    .X(net1071));
 sky130_fd_sc_hd__buf_2 fanout1072 (.A(net1077),
    .X(net1072));
 sky130_fd_sc_hd__buf_2 fanout1073 (.A(net1074),
    .X(net1073));
 sky130_fd_sc_hd__buf_1 fanout1074 (.A(net1077),
    .X(net1074));
 sky130_fd_sc_hd__clkbuf_2 fanout1075 (.A(net1076),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sky130_fd_sc_hd__clkbuf_2 fanout1077 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net1077));
 sky130_fd_sc_hd__buf_2 fanout1078 (.A(net1081),
    .X(net1078));
 sky130_fd_sc_hd__buf_2 fanout1079 (.A(net1081),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_2 fanout1080 (.A(net1081),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_4 fanout1081 (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(net1081));
 sky130_fd_sc_hd__buf_2 fanout1082 (.A(net1085),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_2 fanout1083 (.A(net1085),
    .X(net1083));
 sky130_fd_sc_hd__buf_2 fanout1084 (.A(net1085),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_2 fanout1085 (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(net1085));
 sky130_fd_sc_hd__buf_2 fanout1086 (.A(net1089),
    .X(net1086));
 sky130_fd_sc_hd__buf_2 fanout1087 (.A(net1089),
    .X(net1087));
 sky130_fd_sc_hd__clkbuf_2 fanout1088 (.A(net1089),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_2 fanout1089 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_2 fanout1090 (.A(net1091),
    .X(net1090));
 sky130_fd_sc_hd__buf_2 fanout1091 (.A(net1092),
    .X(net1091));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1092 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net1092));
 sky130_fd_sc_hd__clkbuf_2 fanout1093 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net1093));
 sky130_fd_sc_hd__clkbuf_2 fanout1094 (.A(net1095),
    .X(net1094));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1095 (.A(net1096),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_2 fanout1096 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net1096));
 sky130_fd_sc_hd__clkbuf_2 fanout1097 (.A(net1098),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_2 fanout1098 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net1098));
 sky130_fd_sc_hd__buf_2 fanout1099 (.A(net1102),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_2 fanout1100 (.A(net1101),
    .X(net1100));
 sky130_fd_sc_hd__buf_2 fanout1101 (.A(net1102),
    .X(net1101));
 sky130_fd_sc_hd__clkbuf_2 fanout1102 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net1102));
 sky130_fd_sc_hd__buf_2 fanout1103 (.A(net1105),
    .X(net1103));
 sky130_fd_sc_hd__buf_2 fanout1104 (.A(net1105),
    .X(net1104));
 sky130_fd_sc_hd__buf_2 fanout1105 (.A(net1106),
    .X(net1105));
 sky130_fd_sc_hd__clkbuf_2 fanout1106 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net1106));
 sky130_fd_sc_hd__clkbuf_2 fanout1107 (.A(net1108),
    .X(net1107));
 sky130_fd_sc_hd__clkbuf_2 fanout1108 (.A(net1109),
    .X(net1108));
 sky130_fd_sc_hd__clkbuf_2 fanout1109 (.A(net1110),
    .X(net1109));
 sky130_fd_sc_hd__clkbuf_4 fanout1110 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net1110));
 sky130_fd_sc_hd__clkbuf_2 fanout1111 (.A(net1112),
    .X(net1111));
 sky130_fd_sc_hd__clkbuf_2 fanout1112 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net1112));
 sky130_fd_sc_hd__clkbuf_2 fanout1113 (.A(net1114),
    .X(net1113));
 sky130_fd_sc_hd__clkbuf_2 fanout1114 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net1114));
 sky130_fd_sc_hd__clkbuf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sky130_fd_sc_hd__buf_2 fanout1116 (.A(net1117),
    .X(net1116));
 sky130_fd_sc_hd__clkbuf_2 fanout1117 (.A(net1118),
    .X(net1117));
 sky130_fd_sc_hd__clkbuf_4 fanout1118 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net1118));
 sky130_fd_sc_hd__clkbuf_2 fanout1119 (.A(net1120),
    .X(net1119));
 sky130_fd_sc_hd__buf_2 fanout1120 (.A(net1127),
    .X(net1120));
 sky130_fd_sc_hd__buf_2 fanout1121 (.A(net1122),
    .X(net1121));
 sky130_fd_sc_hd__clkbuf_2 fanout1122 (.A(net1127),
    .X(net1122));
 sky130_fd_sc_hd__buf_2 fanout1123 (.A(net1124),
    .X(net1123));
 sky130_fd_sc_hd__clkbuf_2 fanout1124 (.A(net1127),
    .X(net1124));
 sky130_fd_sc_hd__buf_2 fanout1125 (.A(net1127),
    .X(net1125));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1126 (.A(net1127),
    .X(net1126));
 sky130_fd_sc_hd__buf_4 fanout1127 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net1127));
 sky130_fd_sc_hd__clkbuf_2 fanout1128 (.A(net1136),
    .X(net1128));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1129 (.A(net1136),
    .X(net1129));
 sky130_fd_sc_hd__clkbuf_2 fanout1130 (.A(net1131),
    .X(net1130));
 sky130_fd_sc_hd__clkbuf_2 fanout1131 (.A(net1136),
    .X(net1131));
 sky130_fd_sc_hd__clkbuf_2 fanout1132 (.A(net1133),
    .X(net1132));
 sky130_fd_sc_hd__clkbuf_2 fanout1133 (.A(net1136),
    .X(net1133));
 sky130_fd_sc_hd__buf_2 fanout1134 (.A(net1136),
    .X(net1134));
 sky130_fd_sc_hd__clkbuf_2 fanout1135 (.A(net1136),
    .X(net1135));
 sky130_fd_sc_hd__buf_4 fanout1136 (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(net1136));
 sky130_fd_sc_hd__buf_2 fanout1137 (.A(net1145),
    .X(net1137));
 sky130_fd_sc_hd__buf_2 fanout1138 (.A(net1140),
    .X(net1138));
 sky130_fd_sc_hd__buf_1 fanout1139 (.A(net1140),
    .X(net1139));
 sky130_fd_sc_hd__clkbuf_2 fanout1140 (.A(net1145),
    .X(net1140));
 sky130_fd_sc_hd__clkbuf_2 fanout1141 (.A(net1144),
    .X(net1141));
 sky130_fd_sc_hd__buf_2 fanout1142 (.A(net1143),
    .X(net1142));
 sky130_fd_sc_hd__clkbuf_2 fanout1143 (.A(net1144),
    .X(net1143));
 sky130_fd_sc_hd__buf_2 fanout1144 (.A(net1145),
    .X(net1144));
 sky130_fd_sc_hd__buf_2 fanout1145 (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(net1145));
 sky130_fd_sc_hd__clkbuf_4 fanout1146 (.A(net1153),
    .X(net1146));
 sky130_fd_sc_hd__buf_2 fanout1147 (.A(net1149),
    .X(net1147));
 sky130_fd_sc_hd__buf_1 fanout1148 (.A(net1149),
    .X(net1148));
 sky130_fd_sc_hd__clkbuf_2 fanout1149 (.A(net1153),
    .X(net1149));
 sky130_fd_sc_hd__clkbuf_2 fanout1150 (.A(net1151),
    .X(net1150));
 sky130_fd_sc_hd__clkbuf_2 fanout1151 (.A(net1152),
    .X(net1151));
 sky130_fd_sc_hd__buf_4 fanout1152 (.A(net1153),
    .X(net1152));
 sky130_fd_sc_hd__clkbuf_2 fanout1153 (.A(Tile_X0Y1_FrameStrobe[12]),
    .X(net1153));
 sky130_fd_sc_hd__clkbuf_2 fanout1154 (.A(net1155),
    .X(net1154));
 sky130_fd_sc_hd__buf_2 fanout1155 (.A(net1156),
    .X(net1155));
 sky130_fd_sc_hd__clkbuf_4 fanout1156 (.A(net1157),
    .X(net1156));
 sky130_fd_sc_hd__clkbuf_2 fanout1157 (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(net1157));
 sky130_fd_sc_hd__buf_2 fanout1158 (.A(net1161),
    .X(net1158));
 sky130_fd_sc_hd__buf_2 fanout1159 (.A(net1161),
    .X(net1159));
 sky130_fd_sc_hd__clkbuf_2 fanout1160 (.A(net1161),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_2 fanout1161 (.A(net1162),
    .X(net1161));
 sky130_fd_sc_hd__clkbuf_2 fanout1162 (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(net1162));
 sky130_fd_sc_hd__buf_2 fanout1163 (.A(net1164),
    .X(net1163));
 sky130_fd_sc_hd__buf_2 fanout1164 (.A(net1166),
    .X(net1164));
 sky130_fd_sc_hd__clkbuf_2 fanout1165 (.A(net1166),
    .X(net1165));
 sky130_fd_sc_hd__buf_2 fanout1166 (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net1166));
 sky130_fd_sc_hd__clkbuf_2 fanout1167 (.A(net1170),
    .X(net1167));
 sky130_fd_sc_hd__clkbuf_2 fanout1168 (.A(net1170),
    .X(net1168));
 sky130_fd_sc_hd__buf_2 fanout1169 (.A(net1170),
    .X(net1169));
 sky130_fd_sc_hd__buf_2 fanout1170 (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net1170));
 sky130_fd_sc_hd__clkbuf_2 fanout1171 (.A(net1173),
    .X(net1171));
 sky130_fd_sc_hd__buf_2 fanout1172 (.A(net1173),
    .X(net1172));
 sky130_fd_sc_hd__clkbuf_2 fanout1173 (.A(net1174),
    .X(net1173));
 sky130_fd_sc_hd__clkbuf_2 fanout1174 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net1174));
 sky130_fd_sc_hd__clkbuf_2 fanout1175 (.A(net1178),
    .X(net1175));
 sky130_fd_sc_hd__clkbuf_2 fanout1176 (.A(net1177),
    .X(net1176));
 sky130_fd_sc_hd__buf_2 fanout1177 (.A(net1178),
    .X(net1177));
 sky130_fd_sc_hd__buf_2 fanout1178 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net1178));
 sky130_fd_sc_hd__buf_4 fanout1179 (.A(net172),
    .X(net1179));
 sky130_fd_sc_hd__buf_4 fanout1180 (.A(net171),
    .X(net1180));
 sky130_fd_sc_hd__buf_4 fanout1181 (.A(net170),
    .X(net1181));
 sky130_fd_sc_hd__buf_4 fanout1182 (.A(net169),
    .X(net1182));
 sky130_fd_sc_hd__buf_4 fanout1183 (.A(net168),
    .X(net1183));
 sky130_fd_sc_hd__buf_4 fanout1184 (.A(net167),
    .X(net1184));
 sky130_fd_sc_hd__buf_4 fanout1185 (.A(net166),
    .X(net1185));
 sky130_fd_sc_hd__buf_4 fanout1186 (.A(net1187),
    .X(net1186));
 sky130_fd_sc_hd__clkbuf_2 fanout1187 (.A(Tile_X0Y1_FrameData[31]),
    .X(net1187));
 sky130_fd_sc_hd__buf_4 fanout1188 (.A(net1189),
    .X(net1188));
 sky130_fd_sc_hd__clkbuf_2 fanout1189 (.A(Tile_X0Y1_FrameData[30]),
    .X(net1189));
 sky130_fd_sc_hd__clkbuf_4 fanout1190 (.A(net165),
    .X(net1190));
 sky130_fd_sc_hd__clkbuf_4 fanout1191 (.A(net164),
    .X(net1191));
 sky130_fd_sc_hd__clkbuf_4 fanout1192 (.A(net163),
    .X(net1192));
 sky130_fd_sc_hd__clkbuf_4 fanout1193 (.A(net1194),
    .X(net1193));
 sky130_fd_sc_hd__clkbuf_2 fanout1194 (.A(Tile_X0Y1_FrameData[27]),
    .X(net1194));
 sky130_fd_sc_hd__clkbuf_4 fanout1195 (.A(net162),
    .X(net1195));
 sky130_fd_sc_hd__clkbuf_4 fanout1196 (.A(net161),
    .X(net1196));
 sky130_fd_sc_hd__clkbuf_4 fanout1197 (.A(net160),
    .X(net1197));
 sky130_fd_sc_hd__buf_4 fanout1198 (.A(net159),
    .X(net1198));
 sky130_fd_sc_hd__buf_4 fanout1199 (.A(net158),
    .X(net1199));
 sky130_fd_sc_hd__buf_4 fanout1200 (.A(net157),
    .X(net1200));
 sky130_fd_sc_hd__buf_4 fanout1201 (.A(net156),
    .X(net1201));
 sky130_fd_sc_hd__clkbuf_4 fanout1202 (.A(net155),
    .X(net1202));
 sky130_fd_sc_hd__buf_4 fanout1203 (.A(net154),
    .X(net1203));
 sky130_fd_sc_hd__buf_4 fanout1204 (.A(net153),
    .X(net1204));
 sky130_fd_sc_hd__clkbuf_4 fanout1205 (.A(net152),
    .X(net1205));
 sky130_fd_sc_hd__buf_4 fanout1206 (.A(net1207),
    .X(net1206));
 sky130_fd_sc_hd__clkbuf_2 fanout1207 (.A(Tile_X0Y1_FrameData[16]),
    .X(net1207));
 sky130_fd_sc_hd__buf_4 fanout1208 (.A(net151),
    .X(net1208));
 sky130_fd_sc_hd__buf_4 fanout1209 (.A(net150),
    .X(net1209));
 sky130_fd_sc_hd__clkbuf_4 fanout1210 (.A(net149),
    .X(net1210));
 sky130_fd_sc_hd__buf_4 fanout1211 (.A(net148),
    .X(net1211));
 sky130_fd_sc_hd__buf_4 fanout1212 (.A(net147),
    .X(net1212));
 sky130_fd_sc_hd__buf_4 fanout1213 (.A(net146),
    .X(net1213));
 sky130_fd_sc_hd__clkbuf_4 fanout1214 (.A(net145),
    .X(net1214));
 sky130_fd_sc_hd__buf_2 fanout1215 (.A(net140),
    .X(net1215));
 sky130_fd_sc_hd__clkbuf_4 fanout1216 (.A(net139),
    .X(net1216));
 sky130_fd_sc_hd__clkbuf_4 fanout1217 (.A(net122),
    .X(net1217));
 sky130_fd_sc_hd__buf_4 fanout1218 (.A(net121),
    .X(net1218));
 sky130_fd_sc_hd__clkbuf_4 fanout1219 (.A(net96),
    .X(net1219));
 sky130_fd_sc_hd__buf_4 fanout1220 (.A(net95),
    .X(net1220));
 sky130_fd_sc_hd__buf_4 fanout1221 (.A(net56),
    .X(net1221));
 sky130_fd_sc_hd__clkbuf_4 fanout1222 (.A(net55),
    .X(net1222));
 sky130_fd_sc_hd__buf_4 fanout1223 (.A(net54),
    .X(net1223));
 sky130_fd_sc_hd__buf_4 fanout1224 (.A(net53),
    .X(net1224));
 sky130_fd_sc_hd__buf_4 fanout1225 (.A(net52),
    .X(net1225));
 sky130_fd_sc_hd__buf_4 fanout1226 (.A(net51),
    .X(net1226));
 sky130_fd_sc_hd__buf_4 fanout1227 (.A(net50),
    .X(net1227));
 sky130_fd_sc_hd__buf_4 fanout1228 (.A(net49),
    .X(net1228));
 sky130_fd_sc_hd__buf_4 fanout1229 (.A(net48),
    .X(net1229));
 sky130_fd_sc_hd__buf_4 fanout1230 (.A(net47),
    .X(net1230));
 sky130_fd_sc_hd__buf_4 fanout1231 (.A(net46),
    .X(net1231));
 sky130_fd_sc_hd__clkbuf_4 fanout1232 (.A(net45),
    .X(net1232));
 sky130_fd_sc_hd__buf_4 fanout1233 (.A(net1234),
    .X(net1233));
 sky130_fd_sc_hd__clkbuf_2 fanout1234 (.A(Tile_X0Y0_FrameData[27]),
    .X(net1234));
 sky130_fd_sc_hd__buf_4 fanout1235 (.A(net1236),
    .X(net1235));
 sky130_fd_sc_hd__clkbuf_2 fanout1236 (.A(Tile_X0Y0_FrameData[26]),
    .X(net1236));
 sky130_fd_sc_hd__buf_4 fanout1237 (.A(net44),
    .X(net1237));
 sky130_fd_sc_hd__buf_4 fanout1238 (.A(net43),
    .X(net1238));
 sky130_fd_sc_hd__buf_4 fanout1239 (.A(net42),
    .X(net1239));
 sky130_fd_sc_hd__buf_4 fanout1240 (.A(net41),
    .X(net1240));
 sky130_fd_sc_hd__buf_4 fanout1241 (.A(net40),
    .X(net1241));
 sky130_fd_sc_hd__buf_4 fanout1242 (.A(net39),
    .X(net1242));
 sky130_fd_sc_hd__buf_4 fanout1243 (.A(net38),
    .X(net1243));
 sky130_fd_sc_hd__buf_4 fanout1244 (.A(net37),
    .X(net1244));
 sky130_fd_sc_hd__clkbuf_4 fanout1245 (.A(net36),
    .X(net1245));
 sky130_fd_sc_hd__buf_4 fanout1246 (.A(net35),
    .X(net1246));
 sky130_fd_sc_hd__buf_4 fanout1247 (.A(net34),
    .X(net1247));
 sky130_fd_sc_hd__buf_4 fanout1248 (.A(net33),
    .X(net1248));
 sky130_fd_sc_hd__buf_4 fanout1249 (.A(net32),
    .X(net1249));
 sky130_fd_sc_hd__buf_4 fanout1250 (.A(net31),
    .X(net1250));
 sky130_fd_sc_hd__buf_4 fanout1251 (.A(net30),
    .X(net1251));
 sky130_fd_sc_hd__buf_4 fanout1252 (.A(net29),
    .X(net1252));
 sky130_fd_sc_hd__buf_4 fanout1253 (.A(net28),
    .X(net1253));
 sky130_fd_sc_hd__buf_4 fanout1254 (.A(net27),
    .X(net1254));
 sky130_fd_sc_hd__clkbuf_4 fanout1255 (.A(net22),
    .X(net1255));
 sky130_fd_sc_hd__buf_2 fanout1256 (.A(net21),
    .X(net1256));
 sky130_fd_sc_hd__buf_4 fanout1257 (.A(net4),
    .X(net1257));
 sky130_fd_sc_hd__clkbuf_4 fanout1258 (.A(net3),
    .X(net1258));
 sky130_fd_sc_hd__buf_6 input1 (.A(Tile_X0Y0_E1END[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(Tile_X0Y0_E1END[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(Tile_X0Y0_E1END[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(Tile_X0Y0_E1END[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(Tile_X0Y0_E2END[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(Tile_X0Y0_E2END[1]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(Tile_X0Y0_E2END[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(Tile_X0Y0_E2END[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(Tile_X0Y0_E2END[4]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(Tile_X0Y0_E2END[5]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(Tile_X0Y0_E2END[6]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(Tile_X0Y0_E2END[7]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(Tile_X0Y0_E2MID[0]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(Tile_X0Y0_E2MID[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(Tile_X0Y0_E2MID[2]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(Tile_X0Y0_E2MID[3]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(Tile_X0Y0_E2MID[4]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(Tile_X0Y0_E2MID[5]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(Tile_X0Y0_E2MID[6]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(Tile_X0Y0_E2MID[7]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(Tile_X0Y0_E6END[0]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(Tile_X0Y0_E6END[1]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(Tile_X0Y0_EE4END[0]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(Tile_X0Y0_EE4END[1]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(Tile_X0Y0_EE4END[2]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(Tile_X0Y0_EE4END[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(Tile_X0Y0_FrameData[0]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(Tile_X0Y0_FrameData[10]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(Tile_X0Y0_FrameData[11]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(Tile_X0Y0_FrameData[12]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(Tile_X0Y0_FrameData[13]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(Tile_X0Y0_FrameData[14]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(Tile_X0Y0_FrameData[15]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(Tile_X0Y0_FrameData[16]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(Tile_X0Y0_FrameData[17]),
    .X(net35));
 sky130_fd_sc_hd__buf_2 input36 (.A(Tile_X0Y0_FrameData[18]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(Tile_X0Y0_FrameData[19]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(Tile_X0Y0_FrameData[1]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(Tile_X0Y0_FrameData[20]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input40 (.A(Tile_X0Y0_FrameData[21]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(Tile_X0Y0_FrameData[22]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(Tile_X0Y0_FrameData[23]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(Tile_X0Y0_FrameData[24]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(Tile_X0Y0_FrameData[25]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(Tile_X0Y0_FrameData[28]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(Tile_X0Y0_FrameData[29]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(Tile_X0Y0_FrameData[2]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(Tile_X0Y0_FrameData[30]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(Tile_X0Y0_FrameData[31]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input50 (.A(Tile_X0Y0_FrameData[3]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(Tile_X0Y0_FrameData[4]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(Tile_X0Y0_FrameData[5]),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s2s_1 input53 (.A(Tile_X0Y0_FrameData[6]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(Tile_X0Y0_FrameData[7]),
    .X(net54));
 sky130_fd_sc_hd__buf_2 input55 (.A(Tile_X0Y0_FrameData[8]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(Tile_X0Y0_FrameData[9]),
    .X(net56));
 sky130_fd_sc_hd__buf_8 input57 (.A(Tile_X0Y0_S1END[0]),
    .X(net57));
 sky130_fd_sc_hd__buf_2 input58 (.A(Tile_X0Y0_S1END[1]),
    .X(net58));
 sky130_fd_sc_hd__buf_6 input59 (.A(Tile_X0Y0_S1END[2]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input60 (.A(Tile_X0Y0_S1END[3]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input61 (.A(Tile_X0Y0_S2END[0]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(Tile_X0Y0_S2END[1]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(Tile_X0Y0_S2END[2]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(Tile_X0Y0_S2END[3]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(Tile_X0Y0_S2END[4]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(Tile_X0Y0_S2END[5]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(Tile_X0Y0_S2END[6]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(Tile_X0Y0_S2END[7]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_8 input69 (.A(Tile_X0Y0_S2MID[0]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_8 input70 (.A(Tile_X0Y0_S2MID[1]),
    .X(net70));
 sky130_fd_sc_hd__buf_4 input71 (.A(Tile_X0Y0_S2MID[2]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 input72 (.A(Tile_X0Y0_S2MID[3]),
    .X(net72));
 sky130_fd_sc_hd__buf_4 input73 (.A(Tile_X0Y0_S2MID[4]),
    .X(net73));
 sky130_fd_sc_hd__buf_4 input74 (.A(Tile_X0Y0_S2MID[5]),
    .X(net74));
 sky130_fd_sc_hd__buf_4 input75 (.A(Tile_X0Y0_S2MID[6]),
    .X(net75));
 sky130_fd_sc_hd__buf_4 input76 (.A(Tile_X0Y0_S2MID[7]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(Tile_X0Y0_S4END[0]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 input78 (.A(Tile_X0Y0_S4END[1]),
    .X(net78));
 sky130_fd_sc_hd__buf_2 input79 (.A(Tile_X0Y0_S4END[2]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input80 (.A(Tile_X0Y0_S4END[3]),
    .X(net80));
 sky130_fd_sc_hd__buf_4 input81 (.A(Tile_X0Y0_S4END[4]),
    .X(net81));
 sky130_fd_sc_hd__buf_4 input82 (.A(Tile_X0Y0_S4END[5]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(Tile_X0Y0_S4END[6]),
    .X(net83));
 sky130_fd_sc_hd__buf_4 input84 (.A(Tile_X0Y0_S4END[7]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(Tile_X0Y0_SS4END[0]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(Tile_X0Y0_SS4END[1]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(Tile_X0Y0_SS4END[2]),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 input88 (.A(Tile_X0Y0_SS4END[3]),
    .X(net88));
 sky130_fd_sc_hd__buf_4 input89 (.A(Tile_X0Y0_SS4END[4]),
    .X(net89));
 sky130_fd_sc_hd__buf_4 input90 (.A(Tile_X0Y0_SS4END[5]),
    .X(net90));
 sky130_fd_sc_hd__buf_4 input91 (.A(Tile_X0Y0_SS4END[6]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(Tile_X0Y0_SS4END[7]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(Tile_X0Y0_W1END[0]),
    .X(net93));
 sky130_fd_sc_hd__buf_4 input94 (.A(Tile_X0Y0_W1END[1]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(Tile_X0Y0_W1END[2]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(Tile_X0Y0_W1END[3]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(Tile_X0Y0_W2END[0]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 input98 (.A(Tile_X0Y0_W2END[1]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input99 (.A(Tile_X0Y0_W2END[2]),
    .X(net99));
 sky130_fd_sc_hd__buf_2 input100 (.A(Tile_X0Y0_W2END[3]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 input101 (.A(Tile_X0Y0_W2END[4]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(Tile_X0Y0_W2END[5]),
    .X(net102));
 sky130_fd_sc_hd__dlymetal6s2s_1 input103 (.A(Tile_X0Y0_W2END[6]),
    .X(net103));
 sky130_fd_sc_hd__buf_2 input104 (.A(Tile_X0Y0_W2END[7]),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 input105 (.A(Tile_X0Y0_W2MID[0]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(Tile_X0Y0_W2MID[1]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(Tile_X0Y0_W2MID[2]),
    .X(net107));
 sky130_fd_sc_hd__dlymetal6s2s_1 input108 (.A(Tile_X0Y0_W2MID[3]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(Tile_X0Y0_W2MID[4]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(Tile_X0Y0_W2MID[5]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(Tile_X0Y0_W2MID[6]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(Tile_X0Y0_W2MID[7]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 input113 (.A(Tile_X0Y0_W6END[0]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 input114 (.A(Tile_X0Y0_W6END[1]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(Tile_X0Y0_WW4END[0]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(Tile_X0Y0_WW4END[1]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(Tile_X0Y0_WW4END[2]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(Tile_X0Y0_WW4END[3]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(Tile_X0Y1_E1END[0]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 input120 (.A(Tile_X0Y1_E1END[1]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(Tile_X0Y1_E1END[2]),
    .X(net121));
 sky130_fd_sc_hd__buf_1 input122 (.A(Tile_X0Y1_E1END[3]),
    .X(net122));
 sky130_fd_sc_hd__buf_1 input123 (.A(Tile_X0Y1_E2END[0]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(Tile_X0Y1_E2END[1]),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(Tile_X0Y1_E2END[2]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 input126 (.A(Tile_X0Y1_E2END[3]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(Tile_X0Y1_E2END[4]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(Tile_X0Y1_E2END[5]),
    .X(net128));
 sky130_fd_sc_hd__buf_2 input129 (.A(Tile_X0Y1_E2END[6]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(Tile_X0Y1_E2END[7]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(Tile_X0Y1_E2MID[0]),
    .X(net131));
 sky130_fd_sc_hd__dlymetal6s2s_1 input132 (.A(Tile_X0Y1_E2MID[1]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(Tile_X0Y1_E2MID[2]),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 input134 (.A(Tile_X0Y1_E2MID[3]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(Tile_X0Y1_E2MID[4]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(Tile_X0Y1_E2MID[5]),
    .X(net136));
 sky130_fd_sc_hd__buf_2 input137 (.A(Tile_X0Y1_E2MID[6]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input138 (.A(Tile_X0Y1_E2MID[7]),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 input139 (.A(Tile_X0Y1_E6END[0]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input140 (.A(Tile_X0Y1_E6END[1]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 input141 (.A(Tile_X0Y1_EE4END[0]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(Tile_X0Y1_EE4END[1]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(Tile_X0Y1_EE4END[2]),
    .X(net143));
 sky130_fd_sc_hd__buf_1 input144 (.A(Tile_X0Y1_EE4END[3]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(Tile_X0Y1_FrameData[0]),
    .X(net145));
 sky130_fd_sc_hd__buf_2 input146 (.A(Tile_X0Y1_FrameData[10]),
    .X(net146));
 sky130_fd_sc_hd__buf_2 input147 (.A(Tile_X0Y1_FrameData[11]),
    .X(net147));
 sky130_fd_sc_hd__buf_2 input148 (.A(Tile_X0Y1_FrameData[12]),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input149 (.A(Tile_X0Y1_FrameData[13]),
    .X(net149));
 sky130_fd_sc_hd__buf_2 input150 (.A(Tile_X0Y1_FrameData[14]),
    .X(net150));
 sky130_fd_sc_hd__buf_2 input151 (.A(Tile_X0Y1_FrameData[15]),
    .X(net151));
 sky130_fd_sc_hd__buf_2 input152 (.A(Tile_X0Y1_FrameData[17]),
    .X(net152));
 sky130_fd_sc_hd__buf_2 input153 (.A(Tile_X0Y1_FrameData[18]),
    .X(net153));
 sky130_fd_sc_hd__buf_2 input154 (.A(Tile_X0Y1_FrameData[19]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 input155 (.A(Tile_X0Y1_FrameData[1]),
    .X(net155));
 sky130_fd_sc_hd__buf_2 input156 (.A(Tile_X0Y1_FrameData[20]),
    .X(net156));
 sky130_fd_sc_hd__buf_2 input157 (.A(Tile_X0Y1_FrameData[21]),
    .X(net157));
 sky130_fd_sc_hd__buf_2 input158 (.A(Tile_X0Y1_FrameData[22]),
    .X(net158));
 sky130_fd_sc_hd__buf_2 input159 (.A(Tile_X0Y1_FrameData[23]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input160 (.A(Tile_X0Y1_FrameData[24]),
    .X(net160));
 sky130_fd_sc_hd__buf_2 input161 (.A(Tile_X0Y1_FrameData[25]),
    .X(net161));
 sky130_fd_sc_hd__buf_2 input162 (.A(Tile_X0Y1_FrameData[26]),
    .X(net162));
 sky130_fd_sc_hd__buf_2 input163 (.A(Tile_X0Y1_FrameData[28]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 input164 (.A(Tile_X0Y1_FrameData[29]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 input165 (.A(Tile_X0Y1_FrameData[2]),
    .X(net165));
 sky130_fd_sc_hd__buf_2 input166 (.A(Tile_X0Y1_FrameData[3]),
    .X(net166));
 sky130_fd_sc_hd__buf_2 input167 (.A(Tile_X0Y1_FrameData[4]),
    .X(net167));
 sky130_fd_sc_hd__buf_2 input168 (.A(Tile_X0Y1_FrameData[5]),
    .X(net168));
 sky130_fd_sc_hd__buf_2 input169 (.A(Tile_X0Y1_FrameData[6]),
    .X(net169));
 sky130_fd_sc_hd__buf_2 input170 (.A(Tile_X0Y1_FrameData[7]),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(Tile_X0Y1_FrameData[8]),
    .X(net171));
 sky130_fd_sc_hd__buf_2 input172 (.A(Tile_X0Y1_FrameData[9]),
    .X(net172));
 sky130_fd_sc_hd__buf_4 input173 (.A(Tile_X0Y1_N1END[0]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 input174 (.A(Tile_X0Y1_N1END[1]),
    .X(net174));
 sky130_fd_sc_hd__buf_4 input175 (.A(Tile_X0Y1_N1END[2]),
    .X(net175));
 sky130_fd_sc_hd__buf_4 input176 (.A(Tile_X0Y1_N1END[3]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 input177 (.A(Tile_X0Y1_N2END[0]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 input178 (.A(Tile_X0Y1_N2END[1]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(Tile_X0Y1_N2END[2]),
    .X(net179));
 sky130_fd_sc_hd__buf_2 input180 (.A(Tile_X0Y1_N2END[3]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 input181 (.A(Tile_X0Y1_N2END[4]),
    .X(net181));
 sky130_fd_sc_hd__buf_2 input182 (.A(Tile_X0Y1_N2END[5]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 input183 (.A(Tile_X0Y1_N2END[6]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_4 input184 (.A(Tile_X0Y1_N2END[7]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_8 input185 (.A(Tile_X0Y1_N2MID[0]),
    .X(net185));
 sky130_fd_sc_hd__buf_4 input186 (.A(Tile_X0Y1_N2MID[1]),
    .X(net186));
 sky130_fd_sc_hd__buf_4 input187 (.A(Tile_X0Y1_N2MID[2]),
    .X(net187));
 sky130_fd_sc_hd__buf_4 input188 (.A(Tile_X0Y1_N2MID[3]),
    .X(net188));
 sky130_fd_sc_hd__buf_4 input189 (.A(Tile_X0Y1_N2MID[4]),
    .X(net189));
 sky130_fd_sc_hd__buf_4 input190 (.A(Tile_X0Y1_N2MID[5]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 input191 (.A(Tile_X0Y1_N2MID[6]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_8 input192 (.A(Tile_X0Y1_N2MID[7]),
    .X(net192));
 sky130_fd_sc_hd__dlymetal6s2s_1 input193 (.A(Tile_X0Y1_N4END[0]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 input194 (.A(Tile_X0Y1_N4END[1]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(Tile_X0Y1_N4END[2]),
    .X(net195));
 sky130_fd_sc_hd__buf_2 input196 (.A(Tile_X0Y1_N4END[3]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 input197 (.A(Tile_X0Y1_N4END[4]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 input198 (.A(Tile_X0Y1_N4END[5]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 input199 (.A(Tile_X0Y1_N4END[6]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_4 input200 (.A(Tile_X0Y1_N4END[7]),
    .X(net200));
 sky130_fd_sc_hd__dlymetal6s2s_1 input201 (.A(Tile_X0Y1_NN4END[0]),
    .X(net201));
 sky130_fd_sc_hd__dlymetal6s2s_1 input202 (.A(Tile_X0Y1_NN4END[1]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(Tile_X0Y1_NN4END[2]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 input204 (.A(Tile_X0Y1_NN4END[3]),
    .X(net204));
 sky130_fd_sc_hd__buf_2 input205 (.A(Tile_X0Y1_NN4END[4]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 input206 (.A(Tile_X0Y1_NN4END[5]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 input207 (.A(Tile_X0Y1_NN4END[6]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 input208 (.A(Tile_X0Y1_NN4END[7]),
    .X(net208));
 sky130_fd_sc_hd__buf_4 input209 (.A(Tile_X0Y1_W1END[0]),
    .X(net209));
 sky130_fd_sc_hd__buf_4 input210 (.A(Tile_X0Y1_W1END[1]),
    .X(net210));
 sky130_fd_sc_hd__buf_2 input211 (.A(Tile_X0Y1_W1END[2]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(Tile_X0Y1_W1END[3]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(Tile_X0Y1_W2END[0]),
    .X(net213));
 sky130_fd_sc_hd__buf_2 input214 (.A(Tile_X0Y1_W2END[1]),
    .X(net214));
 sky130_fd_sc_hd__buf_2 input215 (.A(Tile_X0Y1_W2END[2]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 input216 (.A(Tile_X0Y1_W2END[3]),
    .X(net216));
 sky130_fd_sc_hd__buf_2 input217 (.A(Tile_X0Y1_W2END[4]),
    .X(net217));
 sky130_fd_sc_hd__dlymetal6s2s_1 input218 (.A(Tile_X0Y1_W2END[5]),
    .X(net218));
 sky130_fd_sc_hd__dlymetal6s2s_1 input219 (.A(Tile_X0Y1_W2END[6]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 input220 (.A(Tile_X0Y1_W2END[7]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 input221 (.A(Tile_X0Y1_W2MID[0]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 input222 (.A(Tile_X0Y1_W2MID[1]),
    .X(net222));
 sky130_fd_sc_hd__buf_2 input223 (.A(Tile_X0Y1_W2MID[2]),
    .X(net223));
 sky130_fd_sc_hd__buf_2 input224 (.A(Tile_X0Y1_W2MID[3]),
    .X(net224));
 sky130_fd_sc_hd__buf_2 input225 (.A(Tile_X0Y1_W2MID[4]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 input226 (.A(Tile_X0Y1_W2MID[5]),
    .X(net226));
 sky130_fd_sc_hd__buf_2 input227 (.A(Tile_X0Y1_W2MID[6]),
    .X(net227));
 sky130_fd_sc_hd__buf_2 input228 (.A(Tile_X0Y1_W2MID[7]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 input229 (.A(Tile_X0Y1_W6END[0]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 input230 (.A(Tile_X0Y1_W6END[1]),
    .X(net230));
 sky130_fd_sc_hd__buf_2 input231 (.A(Tile_X0Y1_WW4END[0]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 input232 (.A(Tile_X0Y1_WW4END[1]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 input233 (.A(Tile_X0Y1_WW4END[2]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 input234 (.A(Tile_X0Y1_WW4END[3]),
    .X(net234));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(Tile_X0Y0_E1BEG[0]));
 sky130_fd_sc_hd__buf_4 output236 (.A(net236),
    .X(Tile_X0Y0_E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(Tile_X0Y0_E1BEG[2]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(Tile_X0Y0_E1BEG[3]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(Tile_X0Y0_E2BEG[0]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(Tile_X0Y0_E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net241),
    .X(Tile_X0Y0_E2BEG[2]));
 sky130_fd_sc_hd__buf_2 output242 (.A(net242),
    .X(Tile_X0Y0_E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(Tile_X0Y0_E2BEG[4]));
 sky130_fd_sc_hd__buf_6 output244 (.A(net244),
    .X(Tile_X0Y0_E2BEG[5]));
 sky130_fd_sc_hd__buf_2 output245 (.A(net245),
    .X(Tile_X0Y0_E2BEG[6]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .X(Tile_X0Y0_E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(Tile_X0Y0_E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(Tile_X0Y0_E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(Tile_X0Y0_E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output250 (.A(net250),
    .X(Tile_X0Y0_E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(Tile_X0Y0_E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(Tile_X0Y0_E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(Tile_X0Y0_E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(Tile_X0Y0_E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(Tile_X0Y0_E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(Tile_X0Y0_E6BEG[10]));
 sky130_fd_sc_hd__buf_6 output257 (.A(net257),
    .X(Tile_X0Y0_E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(Tile_X0Y0_E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(Tile_X0Y0_E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(Tile_X0Y0_E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(Tile_X0Y0_E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(Tile_X0Y0_E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(Tile_X0Y0_E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(Tile_X0Y0_E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(Tile_X0Y0_E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(Tile_X0Y0_E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(Tile_X0Y0_EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(Tile_X0Y0_EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(Tile_X0Y0_EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(Tile_X0Y0_EE4BEG[12]));
 sky130_fd_sc_hd__buf_6 output271 (.A(net271),
    .X(Tile_X0Y0_EE4BEG[13]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(Tile_X0Y0_EE4BEG[14]));
 sky130_fd_sc_hd__buf_6 output273 (.A(net273),
    .X(Tile_X0Y0_EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(Tile_X0Y0_EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(Tile_X0Y0_EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(Tile_X0Y0_EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(Tile_X0Y0_EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(Tile_X0Y0_EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(Tile_X0Y0_EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(Tile_X0Y0_EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(Tile_X0Y0_EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(Tile_X0Y0_EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(Tile_X0Y0_FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(Tile_X0Y0_FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(Tile_X0Y0_FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(Tile_X0Y0_FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(Tile_X0Y0_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(Tile_X0Y0_FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(Tile_X0Y0_FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(Tile_X0Y0_FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(Tile_X0Y0_FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(Tile_X0Y0_FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(Tile_X0Y0_FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .X(Tile_X0Y0_FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .X(Tile_X0Y0_FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .X(Tile_X0Y0_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(Tile_X0Y0_FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(Tile_X0Y0_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output299 (.A(net299),
    .X(Tile_X0Y0_FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .X(Tile_X0Y0_FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(Tile_X0Y0_FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(Tile_X0Y0_FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output303 (.A(net303),
    .X(Tile_X0Y0_FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(Tile_X0Y0_FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(Tile_X0Y0_FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(Tile_X0Y0_FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(Tile_X0Y0_FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(Tile_X0Y0_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(Tile_X0Y0_FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(Tile_X0Y0_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(Tile_X0Y0_FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(Tile_X0Y0_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(Tile_X0Y0_FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(Tile_X0Y0_FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(Tile_X0Y0_FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(Tile_X0Y0_FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(Tile_X0Y0_FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(Tile_X0Y0_FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .X(Tile_X0Y0_FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(Tile_X0Y0_FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(Tile_X0Y0_FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(Tile_X0Y0_FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(Tile_X0Y0_FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(Tile_X0Y0_FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(Tile_X0Y0_FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(Tile_X0Y0_FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(Tile_X0Y0_FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(Tile_X0Y0_FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(Tile_X0Y0_FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(Tile_X0Y0_FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(Tile_X0Y0_FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(Tile_X0Y0_FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output333 (.A(net333),
    .X(Tile_X0Y0_FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output334 (.A(net334),
    .X(Tile_X0Y0_FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output335 (.A(net335),
    .X(Tile_X0Y0_N1BEG[0]));
 sky130_fd_sc_hd__buf_8 output336 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ),
    .X(Tile_X0Y0_N1BEG[1]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .X(Tile_X0Y0_N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .X(Tile_X0Y0_N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(Tile_X0Y0_N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(Tile_X0Y0_N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(Tile_X0Y0_N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(Tile_X0Y0_N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(Tile_X0Y0_N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output344 (.A(net344),
    .X(Tile_X0Y0_N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net345),
    .X(Tile_X0Y0_N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(Tile_X0Y0_N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .X(Tile_X0Y0_N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output348 (.A(net348),
    .X(Tile_X0Y0_N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output349 (.A(net349),
    .X(Tile_X0Y0_N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output350 (.A(net350),
    .X(Tile_X0Y0_N2BEGb[3]));
 sky130_fd_sc_hd__buf_6 output351 (.A(net351),
    .X(Tile_X0Y0_N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output352 (.A(net352),
    .X(Tile_X0Y0_N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output353 (.A(net353),
    .X(Tile_X0Y0_N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output354 (.A(net354),
    .X(Tile_X0Y0_N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output355 (.A(net355),
    .X(Tile_X0Y0_N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output356 (.A(net356),
    .X(Tile_X0Y0_N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(Tile_X0Y0_N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(Tile_X0Y0_N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(Tile_X0Y0_N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(Tile_X0Y0_N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(Tile_X0Y0_N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(Tile_X0Y0_N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .X(Tile_X0Y0_N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(Tile_X0Y0_N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .X(Tile_X0Y0_N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output366 (.A(net366),
    .X(Tile_X0Y0_N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output367 (.A(net367),
    .X(Tile_X0Y0_N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .X(Tile_X0Y0_N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(Tile_X0Y0_N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .X(Tile_X0Y0_N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(Tile_X0Y0_NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(Tile_X0Y0_NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .X(Tile_X0Y0_NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .X(Tile_X0Y0_NN4BEG[12]));
 sky130_fd_sc_hd__buf_6 output375 (.A(net375),
    .X(Tile_X0Y0_NN4BEG[13]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .X(Tile_X0Y0_NN4BEG[14]));
 sky130_fd_sc_hd__buf_6 output377 (.A(net377),
    .X(Tile_X0Y0_NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net378),
    .X(Tile_X0Y0_NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(Tile_X0Y0_NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output380 (.A(net380),
    .X(Tile_X0Y0_NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net381),
    .X(Tile_X0Y0_NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output382 (.A(net382),
    .X(Tile_X0Y0_NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output383 (.A(net383),
    .X(Tile_X0Y0_NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output384 (.A(net384),
    .X(Tile_X0Y0_NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .X(Tile_X0Y0_NN4BEG[8]));
 sky130_fd_sc_hd__buf_6 output386 (.A(net386),
    .X(Tile_X0Y0_NN4BEG[9]));
 sky130_fd_sc_hd__buf_1 output387 (.A(net387),
    .X(Tile_X0Y0_UserCLKo));
 sky130_fd_sc_hd__buf_2 output388 (.A(net388),
    .X(Tile_X0Y0_W1BEG[0]));
 sky130_fd_sc_hd__buf_4 output389 (.A(net389),
    .X(Tile_X0Y0_W1BEG[1]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net390),
    .X(Tile_X0Y0_W1BEG[2]));
 sky130_fd_sc_hd__buf_2 output391 (.A(net391),
    .X(Tile_X0Y0_W1BEG[3]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .X(Tile_X0Y0_W2BEG[0]));
 sky130_fd_sc_hd__buf_2 output393 (.A(net393),
    .X(Tile_X0Y0_W2BEG[1]));
 sky130_fd_sc_hd__buf_2 output394 (.A(net394),
    .X(Tile_X0Y0_W2BEG[2]));
 sky130_fd_sc_hd__buf_2 output395 (.A(net395),
    .X(Tile_X0Y0_W2BEG[3]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net396),
    .X(Tile_X0Y0_W2BEG[4]));
 sky130_fd_sc_hd__buf_2 output397 (.A(net397),
    .X(Tile_X0Y0_W2BEG[5]));
 sky130_fd_sc_hd__buf_2 output398 (.A(net398),
    .X(Tile_X0Y0_W2BEG[6]));
 sky130_fd_sc_hd__buf_2 output399 (.A(net399),
    .X(Tile_X0Y0_W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output400 (.A(net400),
    .X(Tile_X0Y0_W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output401 (.A(net401),
    .X(Tile_X0Y0_W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output402 (.A(net402),
    .X(Tile_X0Y0_W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output403 (.A(net403),
    .X(Tile_X0Y0_W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output404 (.A(net404),
    .X(Tile_X0Y0_W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output405 (.A(net405),
    .X(Tile_X0Y0_W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output406 (.A(net406),
    .X(Tile_X0Y0_W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output407 (.A(net407),
    .X(Tile_X0Y0_W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output408 (.A(net408),
    .X(Tile_X0Y0_W6BEG[0]));
 sky130_fd_sc_hd__buf_2 output409 (.A(net409),
    .X(Tile_X0Y0_W6BEG[10]));
 sky130_fd_sc_hd__buf_6 output410 (.A(net410),
    .X(Tile_X0Y0_W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output411 (.A(net411),
    .X(Tile_X0Y0_W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output412 (.A(net412),
    .X(Tile_X0Y0_W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output413 (.A(net413),
    .X(Tile_X0Y0_W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output414 (.A(net414),
    .X(Tile_X0Y0_W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .X(Tile_X0Y0_W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output416 (.A(net416),
    .X(Tile_X0Y0_W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output417 (.A(net417),
    .X(Tile_X0Y0_W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output418 (.A(net418),
    .X(Tile_X0Y0_W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output419 (.A(net419),
    .X(Tile_X0Y0_W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output420 (.A(net420),
    .X(Tile_X0Y0_WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output421 (.A(net421),
    .X(Tile_X0Y0_WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output422 (.A(net422),
    .X(Tile_X0Y0_WW4BEG[11]));
 sky130_fd_sc_hd__buf_2 output423 (.A(net423),
    .X(Tile_X0Y0_WW4BEG[12]));
 sky130_fd_sc_hd__buf_6 output424 (.A(net424),
    .X(Tile_X0Y0_WW4BEG[13]));
 sky130_fd_sc_hd__buf_2 output425 (.A(net425),
    .X(Tile_X0Y0_WW4BEG[14]));
 sky130_fd_sc_hd__buf_6 output426 (.A(net426),
    .X(Tile_X0Y0_WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output427 (.A(net427),
    .X(Tile_X0Y0_WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output428 (.A(net428),
    .X(Tile_X0Y0_WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output429 (.A(net429),
    .X(Tile_X0Y0_WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output430 (.A(net430),
    .X(Tile_X0Y0_WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output431 (.A(net431),
    .X(Tile_X0Y0_WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output432 (.A(net432),
    .X(Tile_X0Y0_WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output433 (.A(net433),
    .X(Tile_X0Y0_WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output434 (.A(net434),
    .X(Tile_X0Y0_WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output435 (.A(net435),
    .X(Tile_X0Y0_WW4BEG[9]));
 sky130_fd_sc_hd__buf_2 output436 (.A(net436),
    .X(Tile_X0Y1_E1BEG[0]));
 sky130_fd_sc_hd__buf_2 output437 (.A(net437),
    .X(Tile_X0Y1_E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output438 (.A(net438),
    .X(Tile_X0Y1_E1BEG[2]));
 sky130_fd_sc_hd__buf_2 output439 (.A(net439),
    .X(Tile_X0Y1_E1BEG[3]));
 sky130_fd_sc_hd__buf_2 output440 (.A(net440),
    .X(Tile_X0Y1_E2BEG[0]));
 sky130_fd_sc_hd__buf_2 output441 (.A(net441),
    .X(Tile_X0Y1_E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output442 (.A(net442),
    .X(Tile_X0Y1_E2BEG[2]));
 sky130_fd_sc_hd__buf_2 output443 (.A(net443),
    .X(Tile_X0Y1_E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output444 (.A(net444),
    .X(Tile_X0Y1_E2BEG[4]));
 sky130_fd_sc_hd__buf_2 output445 (.A(net445),
    .X(Tile_X0Y1_E2BEG[5]));
 sky130_fd_sc_hd__buf_8 output446 (.A(net446),
    .X(Tile_X0Y1_E2BEG[6]));
 sky130_fd_sc_hd__buf_6 output447 (.A(net447),
    .X(Tile_X0Y1_E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output448 (.A(net448),
    .X(Tile_X0Y1_E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output449 (.A(net449),
    .X(Tile_X0Y1_E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output450 (.A(net450),
    .X(Tile_X0Y1_E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output451 (.A(net451),
    .X(Tile_X0Y1_E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output452 (.A(net452),
    .X(Tile_X0Y1_E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output453 (.A(net453),
    .X(Tile_X0Y1_E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output454 (.A(net454),
    .X(Tile_X0Y1_E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output455 (.A(net455),
    .X(Tile_X0Y1_E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output456 (.A(net456),
    .X(Tile_X0Y1_E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output457 (.A(net457),
    .X(Tile_X0Y1_E6BEG[10]));
 sky130_fd_sc_hd__buf_6 output458 (.A(net458),
    .X(Tile_X0Y1_E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output459 (.A(net459),
    .X(Tile_X0Y1_E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output460 (.A(net460),
    .X(Tile_X0Y1_E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output461 (.A(net461),
    .X(Tile_X0Y1_E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output462 (.A(net462),
    .X(Tile_X0Y1_E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output463 (.A(net463),
    .X(Tile_X0Y1_E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output464 (.A(net464),
    .X(Tile_X0Y1_E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output465 (.A(net465),
    .X(Tile_X0Y1_E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output466 (.A(net466),
    .X(Tile_X0Y1_E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output467 (.A(net467),
    .X(Tile_X0Y1_E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output468 (.A(net468),
    .X(Tile_X0Y1_EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output469 (.A(net469),
    .X(Tile_X0Y1_EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output470 (.A(net470),
    .X(Tile_X0Y1_EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output471 (.A(net471),
    .X(Tile_X0Y1_EE4BEG[12]));
 sky130_fd_sc_hd__buf_6 output472 (.A(net472),
    .X(Tile_X0Y1_EE4BEG[13]));
 sky130_fd_sc_hd__buf_6 output473 (.A(net473),
    .X(Tile_X0Y1_EE4BEG[14]));
 sky130_fd_sc_hd__buf_8 output474 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ),
    .X(Tile_X0Y1_EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output475 (.A(net475),
    .X(Tile_X0Y1_EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output476 (.A(net476),
    .X(Tile_X0Y1_EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output477 (.A(net477),
    .X(Tile_X0Y1_EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output478 (.A(net478),
    .X(Tile_X0Y1_EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output479 (.A(net479),
    .X(Tile_X0Y1_EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output480 (.A(net480),
    .X(Tile_X0Y1_EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output481 (.A(net481),
    .X(Tile_X0Y1_EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output482 (.A(net482),
    .X(Tile_X0Y1_EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output483 (.A(net483),
    .X(Tile_X0Y1_EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output484 (.A(net484),
    .X(Tile_X0Y1_FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output485 (.A(net485),
    .X(Tile_X0Y1_FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output486 (.A(net486),
    .X(Tile_X0Y1_FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output487 (.A(net487),
    .X(Tile_X0Y1_FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output488 (.A(net488),
    .X(Tile_X0Y1_FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output489 (.A(net489),
    .X(Tile_X0Y1_FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output490 (.A(net490),
    .X(Tile_X0Y1_FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output491 (.A(net491),
    .X(Tile_X0Y1_FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output492 (.A(net492),
    .X(Tile_X0Y1_FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output493 (.A(net493),
    .X(Tile_X0Y1_FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output494 (.A(net494),
    .X(Tile_X0Y1_FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output495 (.A(net495),
    .X(Tile_X0Y1_FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output496 (.A(net496),
    .X(Tile_X0Y1_FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output497 (.A(net497),
    .X(Tile_X0Y1_FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output498 (.A(net498),
    .X(Tile_X0Y1_FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output499 (.A(net499),
    .X(Tile_X0Y1_FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output500 (.A(net500),
    .X(Tile_X0Y1_FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output501 (.A(net501),
    .X(Tile_X0Y1_FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output502 (.A(net502),
    .X(Tile_X0Y1_FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output503 (.A(net503),
    .X(Tile_X0Y1_FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output504 (.A(net504),
    .X(Tile_X0Y1_FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output505 (.A(net505),
    .X(Tile_X0Y1_FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output506 (.A(net506),
    .X(Tile_X0Y1_FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output507 (.A(net507),
    .X(Tile_X0Y1_FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output508 (.A(net508),
    .X(Tile_X0Y1_FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output509 (.A(net509),
    .X(Tile_X0Y1_FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output510 (.A(net510),
    .X(Tile_X0Y1_FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output511 (.A(net511),
    .X(Tile_X0Y1_FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output512 (.A(net512),
    .X(Tile_X0Y1_FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output513 (.A(net513),
    .X(Tile_X0Y1_FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output514 (.A(net514),
    .X(Tile_X0Y1_FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output515 (.A(net515),
    .X(Tile_X0Y1_FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output516 (.A(net516),
    .X(Tile_X0Y1_S1BEG[0]));
 sky130_fd_sc_hd__buf_2 output517 (.A(net517),
    .X(Tile_X0Y1_S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output518 (.A(net518),
    .X(Tile_X0Y1_S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output519 (.A(net519),
    .X(Tile_X0Y1_S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output520 (.A(net520),
    .X(Tile_X0Y1_S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output521 (.A(net521),
    .X(Tile_X0Y1_S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output522 (.A(net522),
    .X(Tile_X0Y1_S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output523 (.A(net523),
    .X(Tile_X0Y1_S2BEG[3]));
 sky130_fd_sc_hd__buf_8 output524 (.A(net524),
    .X(Tile_X0Y1_S2BEG[4]));
 sky130_fd_sc_hd__buf_2 output525 (.A(net525),
    .X(Tile_X0Y1_S2BEG[5]));
 sky130_fd_sc_hd__buf_2 output526 (.A(net526),
    .X(Tile_X0Y1_S2BEG[6]));
 sky130_fd_sc_hd__buf_4 output527 (.A(net527),
    .X(Tile_X0Y1_S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output528 (.A(net528),
    .X(Tile_X0Y1_S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output529 (.A(net529),
    .X(Tile_X0Y1_S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output530 (.A(net530),
    .X(Tile_X0Y1_S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output531 (.A(net531),
    .X(Tile_X0Y1_S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output532 (.A(net532),
    .X(Tile_X0Y1_S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output533 (.A(net533),
    .X(Tile_X0Y1_S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output534 (.A(net534),
    .X(Tile_X0Y1_S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output535 (.A(net535),
    .X(Tile_X0Y1_S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output536 (.A(net536),
    .X(Tile_X0Y1_S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output537 (.A(net537),
    .X(Tile_X0Y1_S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output538 (.A(net538),
    .X(Tile_X0Y1_S4BEG[11]));
 sky130_fd_sc_hd__buf_2 output539 (.A(net539),
    .X(Tile_X0Y1_S4BEG[12]));
 sky130_fd_sc_hd__buf_2 output540 (.A(net540),
    .X(Tile_X0Y1_S4BEG[13]));
 sky130_fd_sc_hd__buf_2 output541 (.A(net541),
    .X(Tile_X0Y1_S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output542 (.A(net542),
    .X(Tile_X0Y1_S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output543 (.A(net543),
    .X(Tile_X0Y1_S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output544 (.A(net544),
    .X(Tile_X0Y1_S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output545 (.A(net545),
    .X(Tile_X0Y1_S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output546 (.A(net546),
    .X(Tile_X0Y1_S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output547 (.A(net547),
    .X(Tile_X0Y1_S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output548 (.A(net548),
    .X(Tile_X0Y1_S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output549 (.A(net549),
    .X(Tile_X0Y1_S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output550 (.A(net550),
    .X(Tile_X0Y1_S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output551 (.A(net551),
    .X(Tile_X0Y1_S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output552 (.A(net552),
    .X(Tile_X0Y1_SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output553 (.A(net553),
    .X(Tile_X0Y1_SS4BEG[10]));
 sky130_fd_sc_hd__buf_6 output554 (.A(net554),
    .X(Tile_X0Y1_SS4BEG[11]));
 sky130_fd_sc_hd__buf_2 output555 (.A(net555),
    .X(Tile_X0Y1_SS4BEG[12]));
 sky130_fd_sc_hd__buf_6 output556 (.A(net556),
    .X(Tile_X0Y1_SS4BEG[13]));
 sky130_fd_sc_hd__buf_2 output557 (.A(net557),
    .X(Tile_X0Y1_SS4BEG[14]));
 sky130_fd_sc_hd__buf_2 output558 (.A(net558),
    .X(Tile_X0Y1_SS4BEG[15]));
 sky130_fd_sc_hd__buf_2 output559 (.A(net559),
    .X(Tile_X0Y1_SS4BEG[1]));
 sky130_fd_sc_hd__buf_2 output560 (.A(net560),
    .X(Tile_X0Y1_SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output561 (.A(net561),
    .X(Tile_X0Y1_SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output562 (.A(net562),
    .X(Tile_X0Y1_SS4BEG[4]));
 sky130_fd_sc_hd__buf_2 output563 (.A(net563),
    .X(Tile_X0Y1_SS4BEG[5]));
 sky130_fd_sc_hd__buf_2 output564 (.A(net564),
    .X(Tile_X0Y1_SS4BEG[6]));
 sky130_fd_sc_hd__buf_2 output565 (.A(net565),
    .X(Tile_X0Y1_SS4BEG[7]));
 sky130_fd_sc_hd__buf_4 output566 (.A(net566),
    .X(Tile_X0Y1_SS4BEG[8]));
 sky130_fd_sc_hd__buf_6 output567 (.A(net567),
    .X(Tile_X0Y1_SS4BEG[9]));
 sky130_fd_sc_hd__buf_2 output568 (.A(net568),
    .X(Tile_X0Y1_W1BEG[0]));
 sky130_fd_sc_hd__buf_2 output569 (.A(net569),
    .X(Tile_X0Y1_W1BEG[1]));
 sky130_fd_sc_hd__buf_2 output570 (.A(net570),
    .X(Tile_X0Y1_W1BEG[2]));
 sky130_fd_sc_hd__buf_2 output571 (.A(net571),
    .X(Tile_X0Y1_W1BEG[3]));
 sky130_fd_sc_hd__buf_2 output572 (.A(net572),
    .X(Tile_X0Y1_W2BEG[0]));
 sky130_fd_sc_hd__buf_2 output573 (.A(net573),
    .X(Tile_X0Y1_W2BEG[1]));
 sky130_fd_sc_hd__buf_2 output574 (.A(net574),
    .X(Tile_X0Y1_W2BEG[2]));
 sky130_fd_sc_hd__buf_2 output575 (.A(net575),
    .X(Tile_X0Y1_W2BEG[3]));
 sky130_fd_sc_hd__buf_2 output576 (.A(net576),
    .X(Tile_X0Y1_W2BEG[4]));
 sky130_fd_sc_hd__buf_6 output577 (.A(net577),
    .X(Tile_X0Y1_W2BEG[5]));
 sky130_fd_sc_hd__buf_6 output578 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ),
    .X(Tile_X0Y1_W2BEG[6]));
 sky130_fd_sc_hd__buf_2 output579 (.A(net579),
    .X(Tile_X0Y1_W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output580 (.A(net580),
    .X(Tile_X0Y1_W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output581 (.A(net581),
    .X(Tile_X0Y1_W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output582 (.A(net582),
    .X(Tile_X0Y1_W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output583 (.A(net583),
    .X(Tile_X0Y1_W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output584 (.A(net584),
    .X(Tile_X0Y1_W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output585 (.A(net585),
    .X(Tile_X0Y1_W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output586 (.A(net586),
    .X(Tile_X0Y1_W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output587 (.A(net587),
    .X(Tile_X0Y1_W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output588 (.A(net588),
    .X(Tile_X0Y1_W6BEG[0]));
 sky130_fd_sc_hd__buf_2 output589 (.A(net589),
    .X(Tile_X0Y1_W6BEG[10]));
 sky130_fd_sc_hd__buf_6 output590 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ),
    .X(Tile_X0Y1_W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output591 (.A(net591),
    .X(Tile_X0Y1_W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output592 (.A(net592),
    .X(Tile_X0Y1_W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output593 (.A(net593),
    .X(Tile_X0Y1_W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output594 (.A(net594),
    .X(Tile_X0Y1_W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output595 (.A(net595),
    .X(Tile_X0Y1_W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output596 (.A(net596),
    .X(Tile_X0Y1_W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output597 (.A(net597),
    .X(Tile_X0Y1_W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output598 (.A(net598),
    .X(Tile_X0Y1_W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output599 (.A(net599),
    .X(Tile_X0Y1_W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output600 (.A(net600),
    .X(Tile_X0Y1_WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output601 (.A(net601),
    .X(Tile_X0Y1_WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output602 (.A(net602),
    .X(Tile_X0Y1_WW4BEG[11]));
 sky130_fd_sc_hd__buf_2 output603 (.A(net603),
    .X(Tile_X0Y1_WW4BEG[12]));
 sky130_fd_sc_hd__buf_6 output604 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ),
    .X(Tile_X0Y1_WW4BEG[13]));
 sky130_fd_sc_hd__buf_4 output605 (.A(net605),
    .X(Tile_X0Y1_WW4BEG[14]));
 sky130_fd_sc_hd__buf_6 output606 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ),
    .X(Tile_X0Y1_WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output607 (.A(net607),
    .X(Tile_X0Y1_WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output608 (.A(net608),
    .X(Tile_X0Y1_WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output609 (.A(net609),
    .X(Tile_X0Y1_WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output610 (.A(net610),
    .X(Tile_X0Y1_WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output611 (.A(net611),
    .X(Tile_X0Y1_WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output612 (.A(net612),
    .X(Tile_X0Y1_WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output613 (.A(net613),
    .X(Tile_X0Y1_WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output614 (.A(net614),
    .X(Tile_X0Y1_WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output615 (.A(net615),
    .X(Tile_X0Y1_WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_2 max_cap616 (.A(_1273_),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_4 wire617 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_Tile_X0Y1_UserCLK (.A(Tile_X0Y1_UserCLK),
    .X(Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_Tile_X0Y1_UserCLK (.A(Tile_X0Y1_UserCLK),
    .X(clknet_0_Tile_X0Y1_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_Tile_X0Y1_UserCLK (.A(clknet_0_Tile_X0Y1_UserCLK),
    .X(clknet_1_0__leaf_Tile_X0Y1_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_Tile_X0Y1_UserCLK_regs (.A(Tile_X0Y1_UserCLK_regs),
    .X(clknet_0_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_Tile_X0Y1_UserCLK_regs (.A(clknet_0_Tile_X0Y1_UserCLK_regs),
    .X(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_Tile_X0Y1_UserCLK_regs (.A(clknet_0_Tile_X0Y1_UserCLK_regs),
    .X(clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_Tile_X0Y1_UserCLK_regs (.A(clknet_0_Tile_X0Y1_UserCLK_regs),
    .X(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_Tile_X0Y1_UserCLK_regs (.A(clknet_0_Tile_X0Y1_UserCLK_regs),
    .X(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs));
 sky130_fd_sc_hd__mux4_2 clone1 (.A0(net980),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .A2(_0382_),
    .A3(net672),
    .S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ),
    .X(net618));
 sky130_fd_sc_hd__buf_6 rebuffer2 (.A(net684),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net619),
    .X(net620));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer4 (.A(net619),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_1158_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(_1158_),
    .X(net623));
 sky130_fd_sc_hd__o21ai_1 clone7 (.A1(\Tile_X0Y1_DSP_bot.A0 ),
    .A2(net1059),
    .B1(_0877_),
    .Y(net624));
 sky130_fd_sc_hd__o21ai_4 clone8 (.A1(net1061),
    .A2(\Tile_X0Y1_DSP_bot.B0 ),
    .B1(_0980_),
    .Y(net625));
 sky130_fd_sc_hd__o21ai_4 clone9 (.A1(\Tile_X0Y1_DSP_bot.B1 ),
    .A2(net1061),
    .B1(_0943_),
    .Y(net626));
 sky130_fd_sc_hd__buf_6 rebuffer10 (.A(_0394_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(_1158_),
    .X(net657));
 sky130_fd_sc_hd__mux2_4 clone41 (.A0(_0298_),
    .A1(_0295_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .X(net658));
 sky130_fd_sc_hd__o21ai_4 clone45 (.A1(net1059),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ),
    .B1(_0728_),
    .Y(net662));
 sky130_fd_sc_hd__clkbuf_2 rebuffer46 (.A(_0217_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net663),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .X(net666));
 sky130_fd_sc_hd__buf_6 rebuffer55 (.A(_0373_),
    .X(net672));
 sky130_fd_sc_hd__buf_6 rebuffer56 (.A(net702),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(net673),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(net673),
    .X(net675));
 sky130_fd_sc_hd__buf_8 clone59 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .X(net676));
 sky130_fd_sc_hd__buf_6 rebuffer67 (.A(net741),
    .X(net684));
 sky130_fd_sc_hd__buf_6 rebuffer71 (.A(_0373_),
    .X(net688));
 sky130_fd_sc_hd__buf_6 rebuffer72 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer73 (.A(net689),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_1 clone75 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_1 clone76 (.A(net742),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer77 (.A(net658),
    .X(net694));
 sky130_fd_sc_hd__buf_6 clone78 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_2 rebuffer85 (.A(_0383_),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer86 (.A(_0381_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer87 (.A(net731),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer88 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer89 (.A(net705),
    .X(net706));
 sky130_fd_sc_hd__buf_8 clone91 (.A(net1010),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_1 clone92 (.A(net1015),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer93 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_2 rebuffer94 (.A(_0213_),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer95 (.A(_0307_),
    .X(net712));
 sky130_fd_sc_hd__buf_8 clone97 (.A(net1001),
    .X(net714));
 sky130_fd_sc_hd__buf_6 clone98 (.A(net981),
    .X(net715));
 sky130_fd_sc_hd__buf_8 clone99 (.A(net994),
    .X(net716));
 sky130_fd_sc_hd__buf_6 rebuffer104 (.A(_0537_),
    .X(net721));
 sky130_fd_sc_hd__o21ai_4 clone105 (.A1(net1060),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ),
    .B1(_0542_),
    .Y(net722));
 sky130_fd_sc_hd__buf_6 clone107 (.A(net1048),
    .X(net724));
 sky130_fd_sc_hd__buf_6 rebuffer108 (.A(_0174_),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_2 rebuffer109 (.A(net746),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer110 (.A(net966),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer111 (.A(net966),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer112 (.A(net728),
    .X(net729));
 sky130_fd_sc_hd__buf_2 rebuffer113 (.A(net999),
    .X(net730));
 sky130_fd_sc_hd__buf_6 rebuffer114 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer115 (.A(net731),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_1 clone116 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__buf_6 clone117 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer118 (.A(\Tile_X0Y1_DSP_bot.A0 ),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_1 clone119 (.A(net1005),
    .X(net736));
 sky130_fd_sc_hd__buf_6 clone120 (.A(net1035),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer121 (.A(_0349_),
    .X(net738));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer122 (.A(_0307_),
    .X(net739));
 sky130_fd_sc_hd__buf_6 clone123 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_2 rebuffer124 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer125 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .X(net742));
 sky130_fd_sc_hd__buf_8 clone126 (.A(net977),
    .X(net743));
 sky130_fd_sc_hd__a22o_4 clone127 (.A1(net745),
    .A2(net725),
    .B1(_0197_),
    .B2(_0198_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer128 (.A(_0185_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer129 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_1 clone130 (.A(net999),
    .X(net747));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_404 ();
endmodule
