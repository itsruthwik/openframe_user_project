magic
tech sky130A
magscale 1 2
timestamp 1746698716
<< viali >>
rect 1593 8585 1627 8619
rect 1961 8585 1995 8619
rect 2329 8585 2363 8619
rect 2697 8585 2731 8619
rect 3065 8585 3099 8619
rect 3433 8585 3467 8619
rect 4169 8585 4203 8619
rect 4537 8585 4571 8619
rect 4905 8585 4939 8619
rect 5273 8585 5307 8619
rect 5641 8585 5675 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 7849 8585 7883 8619
rect 8217 8585 8251 8619
rect 11989 8585 12023 8619
rect 12357 8585 12391 8619
rect 12725 8585 12759 8619
rect 13001 8585 13035 8619
rect 13461 8585 13495 8619
rect 13829 8585 13863 8619
rect 14565 8585 14599 8619
rect 14933 8585 14967 8619
rect 15301 8585 15335 8619
rect 15669 8585 15703 8619
rect 16037 8585 16071 8619
rect 16405 8585 16439 8619
rect 16957 8585 16991 8619
rect 17233 8585 17267 8619
rect 17601 8585 17635 8619
rect 17969 8585 18003 8619
rect 18337 8585 18371 8619
rect 18705 8585 18739 8619
rect 19349 8585 19383 8619
rect 38485 8585 38519 8619
rect 39037 8585 39071 8619
rect 39405 8585 39439 8619
rect 40049 8585 40083 8619
rect 40785 8585 40819 8619
rect 41153 8585 41187 8619
rect 41521 8585 41555 8619
rect 42625 8585 42659 8619
rect 43729 8585 43763 8619
rect 44465 8585 44499 8619
rect 1777 8449 1811 8483
rect 2145 8449 2179 8483
rect 2513 8449 2547 8483
rect 2881 8449 2915 8483
rect 3249 8449 3283 8483
rect 3617 8449 3651 8483
rect 4353 8449 4387 8483
rect 4721 8449 4755 8483
rect 5089 8449 5123 8483
rect 5457 8449 5491 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 8033 8449 8067 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10253 8449 10287 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 11345 8449 11379 8483
rect 11805 8449 11839 8483
rect 12173 8449 12207 8483
rect 12541 8449 12575 8483
rect 13185 8449 13219 8483
rect 13277 8449 13311 8483
rect 13645 8449 13679 8483
rect 14381 8449 14415 8483
rect 14749 8449 14783 8483
rect 15117 8449 15151 8483
rect 15485 8449 15519 8483
rect 15853 8449 15887 8483
rect 16221 8449 16255 8483
rect 16773 8449 16807 8483
rect 17417 8449 17451 8483
rect 17785 8449 17819 8483
rect 18153 8449 18187 8483
rect 18521 8449 18555 8483
rect 18889 8449 18923 8483
rect 19533 8449 19567 8483
rect 38643 8449 38677 8483
rect 38841 8449 38875 8483
rect 39221 8449 39255 8483
rect 39865 8449 39899 8483
rect 40233 8449 40267 8483
rect 40601 8449 40635 8483
rect 40969 8449 41003 8483
rect 41337 8449 41371 8483
rect 41705 8449 41739 8483
rect 42441 8449 42475 8483
rect 42809 8449 42843 8483
rect 43177 8449 43211 8483
rect 43545 8449 43579 8483
rect 43913 8449 43947 8483
rect 44281 8449 44315 8483
rect 40417 8313 40451 8347
rect 41889 8313 41923 8347
rect 42993 8313 43027 8347
rect 43361 8313 43395 8347
rect 44097 8313 44131 8347
rect 8585 8245 8619 8279
rect 9321 8245 9355 8279
rect 9689 8245 9723 8279
rect 10057 8245 10091 8279
rect 10425 8245 10459 8279
rect 10793 8245 10827 8279
rect 11161 8245 11195 8279
rect 1501 8041 1535 8075
rect 3985 8041 4019 8075
rect 6561 8041 6595 8075
rect 9137 8041 9171 8075
rect 10149 8041 10183 8075
rect 10885 8041 10919 8075
rect 12357 8041 12391 8075
rect 14381 8041 14415 8075
rect 15945 8041 15979 8075
rect 16497 8041 16531 8075
rect 16957 8041 16991 8075
rect 17233 8041 17267 8075
rect 17877 8041 17911 8075
rect 25237 8041 25271 8075
rect 27629 8041 27663 8075
rect 30113 8041 30147 8075
rect 38025 8041 38059 8075
rect 40049 8041 40083 8075
rect 40785 8041 40819 8075
rect 42349 8041 42383 8075
rect 42717 8041 42751 8075
rect 43453 8041 43487 8075
rect 44189 8041 44223 8075
rect 1869 7973 1903 8007
rect 9873 7973 9907 8007
rect 10425 7973 10459 8007
rect 11897 7973 11931 8007
rect 12173 7973 12207 8007
rect 25605 7973 25639 8007
rect 26893 7973 26927 8007
rect 26985 7973 27019 8007
rect 28457 7973 28491 8007
rect 43085 7973 43119 8007
rect 26525 7905 26559 7939
rect 1685 7837 1719 7871
rect 2053 7837 2087 7871
rect 2421 7837 2455 7871
rect 4169 7837 4203 7871
rect 6745 7837 6779 7871
rect 9321 7837 9355 7871
rect 9597 7837 9631 7871
rect 9689 7837 9723 7871
rect 10149 7837 10183 7871
rect 10241 7837 10275 7871
rect 10885 7837 10919 7871
rect 10977 7837 11011 7871
rect 11897 7837 11931 7871
rect 11989 7837 12023 7871
rect 12541 7837 12575 7871
rect 14197 7837 14231 7871
rect 15761 7837 15795 7871
rect 16313 7837 16347 7871
rect 16957 7837 16991 7871
rect 17049 7837 17083 7871
rect 17785 7837 17819 7871
rect 18061 7837 18095 7871
rect 19257 7837 19291 7871
rect 19533 7837 19567 7871
rect 21649 7837 21683 7871
rect 21741 7837 21775 7871
rect 25421 7837 25455 7871
rect 25789 7837 25823 7871
rect 26709 7837 26743 7871
rect 27169 7837 27203 7871
rect 27813 7837 27847 7871
rect 28641 7837 28675 7871
rect 29929 7837 29963 7871
rect 36185 7837 36219 7871
rect 38209 7837 38243 7871
rect 39865 7837 39899 7871
rect 40601 7837 40635 7871
rect 41153 7837 41187 7871
rect 41797 7837 41831 7871
rect 42165 7837 42199 7871
rect 42533 7837 42567 7871
rect 42901 7837 42935 7871
rect 43269 7837 43303 7871
rect 43637 7837 43671 7871
rect 44005 7837 44039 7871
rect 5089 7769 5123 7803
rect 5273 7769 5307 7803
rect 2237 7701 2271 7735
rect 9597 7701 9631 7735
rect 11161 7701 11195 7735
rect 19441 7701 19475 7735
rect 21557 7701 21591 7735
rect 21925 7701 21959 7735
rect 36001 7701 36035 7735
rect 41337 7701 41371 7735
rect 41981 7701 42015 7735
rect 43821 7701 43855 7735
rect 1501 7497 1535 7531
rect 9597 7497 9631 7531
rect 12633 7497 12667 7531
rect 14749 7497 14783 7531
rect 15485 7497 15519 7531
rect 21373 7497 21407 7531
rect 36645 7497 36679 7531
rect 42257 7497 42291 7531
rect 42993 7497 43027 7531
rect 43361 7497 43395 7531
rect 43729 7497 43763 7531
rect 44097 7497 44131 7531
rect 44465 7497 44499 7531
rect 15209 7429 15243 7463
rect 41889 7429 41923 7463
rect 1685 7361 1719 7395
rect 9413 7361 9447 7395
rect 12449 7361 12483 7395
rect 14565 7361 14599 7395
rect 15301 7361 15335 7395
rect 21557 7361 21591 7395
rect 28457 7361 28491 7395
rect 34529 7361 34563 7395
rect 36369 7361 36403 7395
rect 36461 7361 36495 7395
rect 41061 7361 41095 7395
rect 42073 7361 42107 7395
rect 42533 7361 42567 7395
rect 42809 7361 42843 7395
rect 43177 7361 43211 7395
rect 43545 7361 43579 7395
rect 43913 7361 43947 7395
rect 44281 7361 44315 7395
rect 28273 7225 28307 7259
rect 34345 7225 34379 7259
rect 36185 7225 36219 7259
rect 41245 7225 41279 7259
rect 42717 7225 42751 7259
rect 41153 6953 41187 6987
rect 13553 6885 13587 6919
rect 43729 6885 43763 6919
rect 12541 6817 12575 6851
rect 13185 6817 13219 6851
rect 12633 6749 12667 6783
rect 12725 6749 12759 6783
rect 13277 6749 13311 6783
rect 13369 6749 13403 6783
rect 14105 6749 14139 6783
rect 20361 6749 20395 6783
rect 22661 6749 22695 6783
rect 25421 6749 25455 6783
rect 37565 6749 37599 6783
rect 40969 6749 41003 6783
rect 42533 6749 42567 6783
rect 42809 6749 42843 6783
rect 43177 6749 43211 6783
rect 43545 6749 43579 6783
rect 43913 6749 43947 6783
rect 44281 6749 44315 6783
rect 12909 6613 12943 6647
rect 14289 6613 14323 6647
rect 20177 6613 20211 6647
rect 22477 6613 22511 6647
rect 25237 6613 25271 6647
rect 37749 6613 37783 6647
rect 42717 6613 42751 6647
rect 42993 6613 43027 6647
rect 43361 6613 43395 6647
rect 44097 6613 44131 6647
rect 44465 6613 44499 6647
rect 22937 6409 22971 6443
rect 44097 6409 44131 6443
rect 44465 6409 44499 6443
rect 20085 6341 20119 6375
rect 16773 6273 16807 6307
rect 16865 6273 16899 6307
rect 19533 6273 19567 6307
rect 20177 6273 20211 6307
rect 20269 6273 20303 6307
rect 23121 6273 23155 6307
rect 27077 6273 27111 6307
rect 27353 6273 27387 6307
rect 28365 6273 28399 6307
rect 35173 6273 35207 6307
rect 36737 6273 36771 6307
rect 43545 6273 43579 6307
rect 43913 6273 43947 6307
rect 44281 6273 44315 6307
rect 34989 6205 35023 6239
rect 19349 6137 19383 6171
rect 28181 6137 28215 6171
rect 16681 6069 16715 6103
rect 17049 6069 17083 6103
rect 20453 6069 20487 6103
rect 27261 6069 27295 6103
rect 36553 6069 36587 6103
rect 43729 6069 43763 6103
rect 18613 5865 18647 5899
rect 44465 5865 44499 5899
rect 30573 5797 30607 5831
rect 34161 5797 34195 5831
rect 14841 5729 14875 5763
rect 18797 5661 18831 5695
rect 25421 5661 25455 5695
rect 29653 5661 29687 5695
rect 29745 5661 29779 5695
rect 30113 5661 30147 5695
rect 30297 5661 30331 5695
rect 30757 5661 30791 5695
rect 34345 5661 34379 5695
rect 43913 5661 43947 5695
rect 44281 5661 44315 5695
rect 14933 5593 14967 5627
rect 15117 5593 15151 5627
rect 15301 5593 15335 5627
rect 25237 5525 25271 5559
rect 29929 5525 29963 5559
rect 30481 5525 30515 5559
rect 44097 5525 44131 5559
rect 23213 5321 23247 5355
rect 44465 5321 44499 5355
rect 22937 5185 22971 5219
rect 23397 5185 23431 5219
rect 24225 5185 24259 5219
rect 31309 5185 31343 5219
rect 33701 5185 33735 5219
rect 43913 5185 43947 5219
rect 44281 5185 44315 5219
rect 23121 5049 23155 5083
rect 24041 5049 24075 5083
rect 33517 5049 33551 5083
rect 44097 5049 44131 5083
rect 31125 4981 31159 5015
rect 18613 4777 18647 4811
rect 41153 4777 41187 4811
rect 44465 4709 44499 4743
rect 18429 4573 18463 4607
rect 18797 4573 18831 4607
rect 19717 4573 19751 4607
rect 19809 4573 19843 4607
rect 33241 4573 33275 4607
rect 39221 4573 39255 4607
rect 40785 4573 40819 4607
rect 40969 4573 41003 4607
rect 43913 4573 43947 4607
rect 44281 4573 44315 4607
rect 18245 4437 18279 4471
rect 19625 4437 19659 4471
rect 19993 4437 20027 4471
rect 33057 4437 33091 4471
rect 39405 4437 39439 4471
rect 44097 4437 44131 4471
rect 16405 4097 16439 4131
rect 21925 4097 21959 4131
rect 22017 4097 22051 4131
rect 23397 4097 23431 4131
rect 23489 4097 23523 4131
rect 24317 4097 24351 4131
rect 24409 4097 24443 4131
rect 25697 4097 25731 4131
rect 25789 4097 25823 4131
rect 26985 4097 27019 4131
rect 27261 4097 27295 4131
rect 32321 4097 32355 4131
rect 43913 4097 43947 4131
rect 44281 4097 44315 4131
rect 16221 3961 16255 3995
rect 23673 3961 23707 3995
rect 27169 3961 27203 3995
rect 44097 3961 44131 3995
rect 44465 3961 44499 3995
rect 21833 3893 21867 3927
rect 22201 3893 22235 3927
rect 23305 3893 23339 3927
rect 24225 3893 24259 3927
rect 24593 3893 24627 3927
rect 25605 3893 25639 3927
rect 25973 3893 26007 3927
rect 32137 3893 32171 3927
rect 9229 3689 9263 3723
rect 11989 3689 12023 3723
rect 13645 3689 13679 3723
rect 14841 3689 14875 3723
rect 17969 3689 18003 3723
rect 44465 3621 44499 3655
rect 9413 3485 9447 3519
rect 12173 3485 12207 3519
rect 13829 3485 13863 3519
rect 15025 3485 15059 3519
rect 18153 3485 18187 3519
rect 19625 3485 19659 3519
rect 19717 3485 19751 3519
rect 19993 3485 20027 3519
rect 22753 3485 22787 3519
rect 43913 3485 43947 3519
rect 44281 3485 44315 3519
rect 19533 3349 19567 3383
rect 19901 3349 19935 3383
rect 20177 3349 20211 3383
rect 22937 3349 22971 3383
rect 44097 3349 44131 3383
rect 2145 3145 2179 3179
rect 9965 3145 9999 3179
rect 15025 3145 15059 3179
rect 21373 3145 21407 3179
rect 21649 3145 21683 3179
rect 24041 3145 24075 3179
rect 30849 3145 30883 3179
rect 36369 3145 36403 3179
rect 38301 3145 38335 3179
rect 44465 3145 44499 3179
rect 10793 3077 10827 3111
rect 11069 3077 11103 3111
rect 11253 3077 11287 3111
rect 2053 3009 2087 3043
rect 8033 3009 8067 3043
rect 9873 3009 9907 3043
rect 12357 3009 12391 3043
rect 14933 3009 14967 3043
rect 15853 3009 15887 3043
rect 15945 3009 15979 3043
rect 17785 3009 17819 3043
rect 17877 3009 17911 3043
rect 18153 3009 18187 3043
rect 20085 3009 20119 3043
rect 20269 3009 20303 3043
rect 21373 3009 21407 3043
rect 21465 3009 21499 3043
rect 23857 3009 23891 3043
rect 24225 3009 24259 3043
rect 24409 3009 24443 3043
rect 25513 3009 25547 3043
rect 26525 3009 26559 3043
rect 27813 3009 27847 3043
rect 27905 3009 27939 3043
rect 30665 3009 30699 3043
rect 36185 3009 36219 3043
rect 37289 3009 37323 3043
rect 38117 3009 38151 3043
rect 43545 3009 43579 3043
rect 43913 3009 43947 3043
rect 44281 3009 44315 3043
rect 8217 2941 8251 2975
rect 12541 2873 12575 2907
rect 37473 2873 37507 2907
rect 44097 2873 44131 2907
rect 15761 2805 15795 2839
rect 16129 2805 16163 2839
rect 17693 2805 17727 2839
rect 18061 2805 18095 2839
rect 18337 2805 18371 2839
rect 20453 2805 20487 2839
rect 24593 2805 24627 2839
rect 25697 2805 25731 2839
rect 26709 2805 26743 2839
rect 27721 2805 27755 2839
rect 28089 2805 28123 2839
rect 43729 2805 43763 2839
rect 42993 2533 43027 2567
rect 43729 2533 43763 2567
rect 44465 2533 44499 2567
rect 42815 2397 42849 2431
rect 43177 2397 43211 2431
rect 43545 2397 43579 2431
rect 43913 2397 43947 2431
rect 44281 2397 44315 2431
rect 43361 2261 43395 2295
rect 44097 2261 44131 2295
<< metal1 >>
rect 16574 11092 16580 11144
rect 16632 11132 16638 11144
rect 34606 11132 34612 11144
rect 16632 11104 34612 11132
rect 16632 11092 16638 11104
rect 34606 11092 34612 11104
rect 34664 11092 34670 11144
rect 18046 11024 18052 11076
rect 18104 11064 18110 11076
rect 33870 11064 33876 11076
rect 18104 11036 33876 11064
rect 18104 11024 18110 11036
rect 33870 11024 33876 11036
rect 33928 11024 33934 11076
rect 16390 10956 16396 11008
rect 16448 10996 16454 11008
rect 20714 10996 20720 11008
rect 16448 10968 20720 10996
rect 16448 10956 16454 10968
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 21358 10956 21364 11008
rect 21416 10996 21422 11008
rect 37274 10996 37280 11008
rect 21416 10968 37280 10996
rect 21416 10956 21422 10968
rect 37274 10956 37280 10968
rect 37332 10956 37338 11008
rect 15470 10888 15476 10940
rect 15528 10928 15534 10940
rect 27706 10928 27712 10940
rect 15528 10900 27712 10928
rect 15528 10888 15534 10900
rect 27706 10888 27712 10900
rect 27764 10888 27770 10940
rect 18782 10752 18788 10804
rect 18840 10792 18846 10804
rect 20346 10792 20352 10804
rect 18840 10764 20352 10792
rect 18840 10752 18846 10764
rect 20346 10752 20352 10764
rect 20404 10752 20410 10804
rect 37182 10004 37188 10056
rect 37240 10044 37246 10056
rect 38010 10044 38016 10056
rect 37240 10016 38016 10044
rect 37240 10004 37246 10016
rect 38010 10004 38016 10016
rect 38068 10004 38074 10056
rect 18598 9664 18604 9716
rect 18656 9704 18662 9716
rect 19610 9704 19616 9716
rect 18656 9676 19616 9704
rect 18656 9664 18662 9676
rect 19610 9664 19616 9676
rect 19668 9664 19674 9716
rect 1118 9392 1124 9444
rect 1176 9432 1182 9444
rect 40954 9432 40960 9444
rect 1176 9404 40960 9432
rect 1176 9392 1182 9404
rect 40954 9392 40960 9404
rect 41012 9392 41018 9444
rect 1026 9324 1032 9376
rect 1084 9364 1090 9376
rect 39666 9364 39672 9376
rect 1084 9336 39672 9364
rect 1084 9324 1090 9336
rect 39666 9324 39672 9336
rect 39724 9324 39730 9376
rect 9858 9256 9864 9308
rect 9916 9296 9922 9308
rect 31110 9296 31116 9308
rect 9916 9268 31116 9296
rect 9916 9256 9922 9268
rect 31110 9256 31116 9268
rect 31168 9256 31174 9308
rect 4338 9188 4344 9240
rect 4396 9228 4402 9240
rect 10318 9228 10324 9240
rect 4396 9200 10324 9228
rect 4396 9188 4402 9200
rect 10318 9188 10324 9200
rect 10376 9188 10382 9240
rect 16942 9188 16948 9240
rect 17000 9228 17006 9240
rect 34330 9228 34336 9240
rect 17000 9200 34336 9228
rect 17000 9188 17006 9200
rect 34330 9188 34336 9200
rect 34388 9188 34394 9240
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 21358 9160 21364 9172
rect 12492 9132 21364 9160
rect 12492 9120 12498 9132
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 27614 9120 27620 9172
rect 27672 9160 27678 9172
rect 39574 9160 39580 9172
rect 27672 9132 39580 9160
rect 27672 9120 27678 9132
rect 39574 9120 39580 9132
rect 39632 9120 39638 9172
rect 3602 9052 3608 9104
rect 3660 9092 3666 9104
rect 8294 9092 8300 9104
rect 3660 9064 8300 9092
rect 3660 9052 3666 9064
rect 8294 9052 8300 9064
rect 8352 9052 8358 9104
rect 17862 9092 17868 9104
rect 10612 9064 17868 9092
rect 1762 8984 1768 9036
rect 1820 9024 1826 9036
rect 1820 8996 2774 9024
rect 1820 8984 1826 8996
rect 2746 8956 2774 8996
rect 9646 8996 9904 9024
rect 9646 8956 9674 8996
rect 2746 8928 9674 8956
rect 9876 8956 9904 8996
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 10612 9024 10640 9064
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 19610 9052 19616 9104
rect 19668 9092 19674 9104
rect 22554 9092 22560 9104
rect 19668 9064 22560 9092
rect 19668 9052 19674 9064
rect 22554 9052 22560 9064
rect 22612 9052 22618 9104
rect 32674 9052 32680 9104
rect 32732 9092 32738 9104
rect 42794 9092 42800 9104
rect 32732 9064 42800 9092
rect 32732 9052 32738 9064
rect 42794 9052 42800 9064
rect 42852 9052 42858 9104
rect 10284 8996 10640 9024
rect 10284 8984 10290 8996
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 10928 8996 14412 9024
rect 10928 8984 10934 8996
rect 9876 8928 10456 8956
rect 2498 8848 2504 8900
rect 2556 8888 2562 8900
rect 5442 8888 5448 8900
rect 2556 8860 5448 8888
rect 2556 8848 2562 8860
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 10428 8888 10456 8928
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 14274 8956 14280 8968
rect 10560 8928 14280 8956
rect 10560 8916 10566 8928
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 14384 8956 14412 8996
rect 15654 8984 15660 9036
rect 15712 9024 15718 9036
rect 35434 9024 35440 9036
rect 15712 8996 35440 9024
rect 15712 8984 15718 8996
rect 35434 8984 35440 8996
rect 35492 8984 35498 9036
rect 37182 8956 37188 8968
rect 14384 8928 37188 8956
rect 37182 8916 37188 8928
rect 37240 8916 37246 8968
rect 40770 8916 40776 8968
rect 40828 8956 40834 8968
rect 43990 8956 43996 8968
rect 40828 8928 43996 8956
rect 40828 8916 40834 8928
rect 43990 8916 43996 8928
rect 44048 8916 44054 8968
rect 36446 8888 36452 8900
rect 10428 8860 36452 8888
rect 36446 8848 36452 8860
rect 36504 8848 36510 8900
rect 40034 8848 40040 8900
rect 40092 8888 40098 8900
rect 43530 8888 43536 8900
rect 40092 8860 43536 8888
rect 40092 8848 40098 8860
rect 43530 8848 43536 8860
rect 43588 8848 43594 8900
rect 3510 8780 3516 8832
rect 3568 8820 3574 8832
rect 11238 8820 11244 8832
rect 3568 8792 11244 8820
rect 3568 8780 3574 8792
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 13538 8820 13544 8832
rect 11388 8792 13544 8820
rect 11388 8780 11394 8792
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 33778 8780 33784 8832
rect 33836 8820 33842 8832
rect 42886 8820 42892 8832
rect 33836 8792 42892 8820
rect 33836 8780 33842 8792
rect 42886 8780 42892 8792
rect 42944 8780 42950 8832
rect 1104 8730 44896 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 44896 8730
rect 1104 8656 44896 8678
rect 1578 8576 1584 8628
rect 1636 8576 1642 8628
rect 1946 8576 1952 8628
rect 2004 8576 2010 8628
rect 2314 8576 2320 8628
rect 2372 8576 2378 8628
rect 2682 8576 2688 8628
rect 2740 8576 2746 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3053 8619 3111 8625
rect 3053 8616 3065 8619
rect 2924 8588 3065 8616
rect 2924 8576 2930 8588
rect 3053 8585 3065 8588
rect 3099 8585 3111 8619
rect 3053 8579 3111 8585
rect 3418 8576 3424 8628
rect 3476 8576 3482 8628
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 4522 8576 4528 8628
rect 4580 8576 4586 8628
rect 4890 8576 4896 8628
rect 4948 8576 4954 8628
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 6730 8576 6736 8628
rect 6788 8576 6794 8628
rect 7098 8576 7104 8628
rect 7156 8576 7162 8628
rect 7466 8576 7472 8628
rect 7524 8576 7530 8628
rect 7834 8576 7840 8628
rect 7892 8576 7898 8628
rect 8202 8576 8208 8628
rect 8260 8576 8266 8628
rect 11238 8616 11244 8628
rect 8312 8588 11244 8616
rect 8312 8548 8340 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11882 8576 11888 8628
rect 11940 8616 11946 8628
rect 11977 8619 12035 8625
rect 11977 8616 11989 8619
rect 11940 8588 11989 8616
rect 11940 8576 11946 8588
rect 11977 8585 11989 8588
rect 12023 8585 12035 8619
rect 11977 8579 12035 8585
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12345 8619 12403 8625
rect 12345 8616 12357 8619
rect 12308 8588 12357 8616
rect 12308 8576 12314 8588
rect 12345 8585 12357 8588
rect 12391 8585 12403 8619
rect 12345 8579 12403 8585
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 12713 8619 12771 8625
rect 12713 8616 12725 8619
rect 12676 8588 12725 8616
rect 12676 8576 12682 8588
rect 12713 8585 12725 8588
rect 12759 8585 12771 8619
rect 12713 8579 12771 8585
rect 12986 8576 12992 8628
rect 13044 8576 13050 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 13412 8588 13461 8616
rect 13412 8576 13418 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 13780 8588 13829 8616
rect 13780 8576 13786 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 13817 8579 13875 8585
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14516 8588 14565 8616
rect 14516 8576 14522 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14553 8579 14611 8585
rect 14826 8576 14832 8628
rect 14884 8616 14890 8628
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 14884 8588 14933 8616
rect 14884 8576 14890 8588
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 14921 8579 14979 8585
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15378 8616 15384 8628
rect 15335 8588 15384 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15620 8588 15669 8616
rect 15620 8576 15626 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15988 8588 16037 8616
rect 15988 8576 15994 8588
rect 16025 8585 16037 8588
rect 16071 8585 16083 8619
rect 16025 8579 16083 8585
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16393 8619 16451 8625
rect 16393 8616 16405 8619
rect 16356 8588 16405 8616
rect 16356 8576 16362 8588
rect 16393 8585 16405 8588
rect 16439 8585 16451 8619
rect 16393 8579 16451 8585
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 16724 8588 16957 8616
rect 16724 8576 16730 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 16945 8579 17003 8585
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 17092 8588 17233 8616
rect 17092 8576 17098 8588
rect 17221 8585 17233 8588
rect 17267 8585 17279 8619
rect 17221 8579 17279 8585
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 17589 8619 17647 8625
rect 17589 8616 17601 8619
rect 17460 8588 17601 8616
rect 17460 8576 17466 8588
rect 17589 8585 17601 8588
rect 17635 8585 17647 8619
rect 17589 8579 17647 8585
rect 17770 8576 17776 8628
rect 17828 8616 17834 8628
rect 17957 8619 18015 8625
rect 17957 8616 17969 8619
rect 17828 8588 17969 8616
rect 17828 8576 17834 8588
rect 17957 8585 17969 8588
rect 18003 8585 18015 8619
rect 17957 8579 18015 8585
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 18325 8619 18383 8625
rect 18325 8616 18337 8619
rect 18196 8588 18337 8616
rect 18196 8576 18202 8588
rect 18325 8585 18337 8588
rect 18371 8585 18383 8619
rect 18325 8579 18383 8585
rect 18506 8576 18512 8628
rect 18564 8616 18570 8628
rect 18693 8619 18751 8625
rect 18693 8616 18705 8619
rect 18564 8588 18705 8616
rect 18564 8576 18570 8588
rect 18693 8585 18705 8588
rect 18739 8585 18751 8619
rect 18693 8579 18751 8585
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 18932 8588 19349 8616
rect 18932 8576 18938 8588
rect 19337 8585 19349 8588
rect 19383 8585 19395 8619
rect 19337 8579 19395 8585
rect 38378 8576 38384 8628
rect 38436 8616 38442 8628
rect 38473 8619 38531 8625
rect 38473 8616 38485 8619
rect 38436 8588 38485 8616
rect 38436 8576 38442 8588
rect 38473 8585 38485 8588
rect 38519 8585 38531 8619
rect 38473 8579 38531 8585
rect 38562 8576 38568 8628
rect 38620 8616 38626 8628
rect 38654 8616 38660 8628
rect 38620 8588 38660 8616
rect 38620 8576 38626 8588
rect 38654 8576 38660 8588
rect 38712 8576 38718 8628
rect 38764 8588 38976 8616
rect 9582 8548 9588 8560
rect 2884 8520 8340 8548
rect 8404 8520 9588 8548
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 1780 8344 1808 8443
rect 2148 8412 2176 8443
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2884 8489 2912 8520
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8480 3295 8483
rect 3510 8480 3516 8492
rect 3283 8452 3516 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3602 8440 3608 8492
rect 3660 8440 3666 8492
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 5166 8412 5172 8424
rect 2148 8384 5172 8412
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 5460 8412 5488 8443
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6914 8440 6920 8492
rect 6972 8440 6978 8492
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 7834 8440 7840 8492
rect 7892 8480 7898 8492
rect 8404 8489 8432 8520
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 25774 8548 25780 8560
rect 9784 8520 12664 8548
rect 8021 8483 8079 8489
rect 8021 8480 8033 8483
rect 7892 8452 8033 8480
rect 7892 8440 7898 8452
rect 8021 8449 8033 8452
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8480 8815 8483
rect 9398 8480 9404 8492
rect 8803 8452 9404 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9674 8480 9680 8492
rect 9539 8452 9680 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 9784 8412 9812 8520
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10241 8483 10299 8489
rect 10241 8449 10253 8483
rect 10287 8480 10299 8483
rect 10502 8480 10508 8492
rect 10287 8452 10508 8480
rect 10287 8449 10299 8452
rect 10241 8443 10299 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 10594 8440 10600 8492
rect 10652 8440 10658 8492
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 11330 8440 11336 8492
rect 11388 8440 11394 8492
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 5460 8384 9812 8412
rect 10686 8372 10692 8424
rect 10744 8412 10750 8424
rect 11808 8412 11836 8443
rect 10744 8384 11836 8412
rect 10744 8372 10750 8384
rect 10226 8344 10232 8356
rect 1780 8316 10232 8344
rect 10226 8304 10232 8316
rect 10284 8304 10290 8356
rect 10502 8304 10508 8356
rect 10560 8344 10566 8356
rect 12176 8344 12204 8443
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 12308 8452 12541 8480
rect 12308 8440 12314 8452
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 12636 8412 12664 8520
rect 13188 8520 25780 8548
rect 13188 8489 13216 8520
rect 25774 8508 25780 8520
rect 25832 8508 25838 8560
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 13262 8440 13268 8492
rect 13320 8440 13326 8492
rect 13630 8440 13636 8492
rect 13688 8440 13694 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 13780 8452 14381 8480
rect 13780 8440 13786 8452
rect 14369 8449 14381 8452
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 14734 8440 14740 8492
rect 14792 8440 14798 8492
rect 14826 8440 14832 8492
rect 14884 8480 14890 8492
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14884 8452 15117 8480
rect 14884 8440 14890 8452
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 15378 8440 15384 8492
rect 15436 8480 15442 8492
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15436 8452 15485 8480
rect 15436 8440 15442 8452
rect 15473 8449 15485 8452
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 16206 8440 16212 8492
rect 16264 8440 16270 8492
rect 16482 8440 16488 8492
rect 16540 8480 16546 8492
rect 16761 8483 16819 8489
rect 16761 8480 16773 8483
rect 16540 8452 16773 8480
rect 16540 8440 16546 8452
rect 16761 8449 16773 8452
rect 16807 8449 16819 8483
rect 16761 8443 16819 8449
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17770 8440 17776 8492
rect 17828 8440 17834 8492
rect 18138 8440 18144 8492
rect 18196 8440 18202 8492
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18524 8412 18552 8443
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8480 19579 8483
rect 20622 8480 20628 8492
rect 19567 8452 20628 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 37274 8440 37280 8492
rect 37332 8480 37338 8492
rect 38631 8483 38689 8489
rect 38631 8480 38643 8483
rect 37332 8452 38643 8480
rect 37332 8440 37338 8452
rect 38631 8449 38643 8452
rect 38677 8449 38689 8483
rect 38631 8443 38689 8449
rect 19242 8412 19248 8424
rect 12636 8384 16574 8412
rect 18524 8384 19248 8412
rect 10560 8316 12204 8344
rect 10560 8304 10566 8316
rect 12894 8304 12900 8356
rect 12952 8344 12958 8356
rect 13722 8344 13728 8356
rect 12952 8316 13728 8344
rect 12952 8304 12958 8316
rect 13722 8304 13728 8316
rect 13780 8304 13786 8356
rect 16546 8344 16574 8384
rect 19242 8372 19248 8384
rect 19300 8372 19306 8424
rect 26694 8372 26700 8424
rect 26752 8412 26758 8424
rect 33778 8412 33784 8424
rect 26752 8384 33784 8412
rect 26752 8372 26758 8384
rect 33778 8372 33784 8384
rect 33836 8372 33842 8424
rect 38286 8372 38292 8424
rect 38344 8412 38350 8424
rect 38764 8412 38792 8588
rect 38948 8548 38976 8588
rect 39022 8576 39028 8628
rect 39080 8576 39086 8628
rect 39390 8576 39396 8628
rect 39448 8576 39454 8628
rect 39482 8576 39488 8628
rect 39540 8616 39546 8628
rect 40037 8619 40095 8625
rect 40037 8616 40049 8619
rect 39540 8588 40049 8616
rect 39540 8576 39546 8588
rect 40037 8585 40049 8588
rect 40083 8585 40095 8619
rect 40037 8579 40095 8585
rect 40218 8576 40224 8628
rect 40276 8616 40282 8628
rect 40773 8619 40831 8625
rect 40773 8616 40785 8619
rect 40276 8588 40785 8616
rect 40276 8576 40282 8588
rect 40773 8585 40785 8588
rect 40819 8585 40831 8619
rect 40773 8579 40831 8585
rect 40862 8576 40868 8628
rect 40920 8616 40926 8628
rect 41141 8619 41199 8625
rect 41141 8616 41153 8619
rect 40920 8588 41153 8616
rect 40920 8576 40926 8588
rect 41141 8585 41153 8588
rect 41187 8585 41199 8619
rect 41141 8579 41199 8585
rect 41230 8576 41236 8628
rect 41288 8616 41294 8628
rect 41509 8619 41567 8625
rect 41509 8616 41521 8619
rect 41288 8588 41521 8616
rect 41288 8576 41294 8588
rect 41509 8585 41521 8588
rect 41555 8585 41567 8619
rect 41509 8579 41567 8585
rect 41690 8576 41696 8628
rect 41748 8616 41754 8628
rect 42613 8619 42671 8625
rect 42613 8616 42625 8619
rect 41748 8588 42625 8616
rect 41748 8576 41754 8588
rect 42613 8585 42625 8588
rect 42659 8585 42671 8619
rect 42613 8579 42671 8585
rect 43254 8576 43260 8628
rect 43312 8616 43318 8628
rect 43717 8619 43775 8625
rect 43717 8616 43729 8619
rect 43312 8588 43729 8616
rect 43312 8576 43318 8588
rect 43717 8585 43729 8588
rect 43763 8585 43775 8619
rect 43717 8579 43775 8585
rect 44453 8619 44511 8625
rect 44453 8585 44465 8619
rect 44499 8585 44511 8619
rect 44453 8579 44511 8585
rect 38948 8520 39252 8548
rect 39224 8489 39252 8520
rect 43622 8508 43628 8560
rect 43680 8548 43686 8560
rect 44468 8548 44496 8579
rect 43680 8520 44496 8548
rect 43680 8508 43686 8520
rect 38829 8483 38887 8489
rect 38829 8449 38841 8483
rect 38875 8476 38887 8483
rect 39209 8483 39267 8489
rect 38829 8443 38844 8449
rect 38838 8424 38844 8443
rect 38896 8424 38902 8476
rect 39209 8449 39221 8483
rect 39255 8449 39267 8483
rect 39209 8443 39267 8449
rect 39574 8440 39580 8492
rect 39632 8480 39638 8492
rect 39853 8483 39911 8489
rect 39853 8480 39865 8483
rect 39632 8452 39865 8480
rect 39632 8440 39638 8452
rect 39853 8449 39865 8452
rect 39899 8449 39911 8483
rect 39853 8443 39911 8449
rect 40218 8440 40224 8492
rect 40276 8440 40282 8492
rect 40589 8483 40647 8489
rect 40589 8449 40601 8483
rect 40635 8449 40647 8483
rect 40589 8443 40647 8449
rect 40604 8412 40632 8443
rect 40862 8440 40868 8492
rect 40920 8480 40926 8492
rect 40957 8483 41015 8489
rect 40957 8480 40969 8483
rect 40920 8452 40969 8480
rect 40920 8440 40926 8452
rect 40957 8449 40969 8452
rect 41003 8449 41015 8483
rect 41325 8483 41383 8489
rect 41325 8480 41337 8483
rect 40957 8443 41015 8449
rect 41064 8452 41337 8480
rect 38344 8384 38792 8412
rect 39040 8384 40632 8412
rect 38344 8372 38350 8384
rect 23382 8344 23388 8356
rect 16546 8316 23388 8344
rect 23382 8304 23388 8316
rect 23440 8304 23446 8356
rect 35710 8304 35716 8356
rect 35768 8344 35774 8356
rect 35768 8316 38332 8344
rect 35768 8304 35774 8316
rect 8570 8236 8576 8288
rect 8628 8236 8634 8288
rect 9306 8236 9312 8288
rect 9364 8236 9370 8288
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 9677 8279 9735 8285
rect 9677 8276 9689 8279
rect 9548 8248 9689 8276
rect 9548 8236 9554 8248
rect 9677 8245 9689 8248
rect 9723 8245 9735 8279
rect 9677 8239 9735 8245
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10045 8279 10103 8285
rect 10045 8276 10057 8279
rect 10008 8248 10057 8276
rect 10008 8236 10014 8248
rect 10045 8245 10057 8248
rect 10091 8245 10103 8279
rect 10045 8239 10103 8245
rect 10410 8236 10416 8288
rect 10468 8236 10474 8288
rect 10778 8236 10784 8288
rect 10836 8236 10842 8288
rect 11146 8236 11152 8288
rect 11204 8236 11210 8288
rect 18138 8236 18144 8288
rect 18196 8276 18202 8288
rect 37826 8276 37832 8288
rect 18196 8248 37832 8276
rect 18196 8236 18202 8248
rect 37826 8236 37832 8248
rect 37884 8236 37890 8288
rect 38304 8276 38332 8316
rect 38378 8304 38384 8356
rect 38436 8344 38442 8356
rect 38654 8344 38660 8356
rect 38436 8316 38660 8344
rect 38436 8304 38442 8316
rect 38654 8304 38660 8316
rect 38712 8304 38718 8356
rect 39040 8344 39068 8384
rect 40678 8372 40684 8424
rect 40736 8412 40742 8424
rect 41064 8412 41092 8452
rect 41325 8449 41337 8452
rect 41371 8449 41383 8483
rect 41325 8443 41383 8449
rect 41690 8440 41696 8492
rect 41748 8440 41754 8492
rect 42429 8483 42487 8489
rect 42429 8449 42441 8483
rect 42475 8449 42487 8483
rect 42429 8443 42487 8449
rect 42444 8412 42472 8443
rect 42794 8440 42800 8492
rect 42852 8440 42858 8492
rect 42886 8440 42892 8492
rect 42944 8480 42950 8492
rect 43165 8483 43223 8489
rect 43165 8480 43177 8483
rect 42944 8452 43177 8480
rect 42944 8440 42950 8452
rect 43165 8449 43177 8452
rect 43211 8449 43223 8483
rect 43165 8443 43223 8449
rect 43254 8440 43260 8492
rect 43312 8480 43318 8492
rect 43312 8452 43484 8480
rect 43312 8440 43318 8452
rect 40736 8384 41092 8412
rect 41156 8384 42472 8412
rect 40736 8372 40742 8384
rect 38948 8316 39068 8344
rect 38948 8276 38976 8316
rect 39850 8304 39856 8356
rect 39908 8344 39914 8356
rect 40405 8347 40463 8353
rect 40405 8344 40417 8347
rect 39908 8316 40417 8344
rect 39908 8304 39914 8316
rect 40405 8313 40417 8316
rect 40451 8313 40463 8347
rect 41156 8344 41184 8384
rect 42518 8372 42524 8424
rect 42576 8412 42582 8424
rect 43456 8412 43484 8452
rect 43530 8440 43536 8492
rect 43588 8440 43594 8492
rect 43901 8483 43959 8489
rect 43901 8449 43913 8483
rect 43947 8449 43959 8483
rect 43901 8443 43959 8449
rect 43916 8412 43944 8443
rect 43990 8440 43996 8492
rect 44048 8480 44054 8492
rect 44269 8483 44327 8489
rect 44269 8480 44281 8483
rect 44048 8452 44281 8480
rect 44048 8440 44054 8452
rect 44269 8449 44281 8452
rect 44315 8449 44327 8483
rect 44269 8443 44327 8449
rect 42576 8384 43392 8412
rect 43456 8384 43944 8412
rect 42576 8372 42582 8384
rect 40405 8307 40463 8313
rect 40512 8316 41184 8344
rect 38304 8248 38976 8276
rect 39942 8236 39948 8288
rect 40000 8276 40006 8288
rect 40512 8276 40540 8316
rect 41322 8304 41328 8356
rect 41380 8344 41386 8356
rect 41877 8347 41935 8353
rect 41877 8344 41889 8347
rect 41380 8316 41889 8344
rect 41380 8304 41386 8316
rect 41877 8313 41889 8316
rect 41923 8313 41935 8347
rect 41877 8307 41935 8313
rect 42058 8304 42064 8356
rect 42116 8344 42122 8356
rect 43364 8353 43392 8384
rect 42981 8347 43039 8353
rect 42981 8344 42993 8347
rect 42116 8316 42993 8344
rect 42116 8304 42122 8316
rect 42981 8313 42993 8316
rect 43027 8313 43039 8347
rect 42981 8307 43039 8313
rect 43349 8347 43407 8353
rect 43349 8313 43361 8347
rect 43395 8313 43407 8347
rect 43349 8307 43407 8313
rect 43438 8304 43444 8356
rect 43496 8344 43502 8356
rect 44085 8347 44143 8353
rect 44085 8344 44097 8347
rect 43496 8316 44097 8344
rect 43496 8304 43502 8316
rect 44085 8313 44097 8316
rect 44131 8313 44143 8347
rect 44085 8307 44143 8313
rect 40000 8248 40540 8276
rect 40000 8236 40006 8248
rect 42334 8236 42340 8288
rect 42392 8276 42398 8288
rect 44634 8276 44640 8288
rect 42392 8248 44640 8276
rect 42392 8236 42398 8248
rect 44634 8236 44640 8248
rect 44692 8236 44698 8288
rect 1104 8186 44896 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 43950 8186
rect 44002 8134 44014 8186
rect 44066 8134 44078 8186
rect 44130 8134 44142 8186
rect 44194 8134 44206 8186
rect 44258 8134 44896 8186
rect 1104 8112 44896 8134
rect 1210 8032 1216 8084
rect 1268 8072 1274 8084
rect 1489 8075 1547 8081
rect 1489 8072 1501 8075
rect 1268 8044 1501 8072
rect 1268 8032 1274 8044
rect 1489 8041 1501 8044
rect 1535 8041 1547 8075
rect 1489 8035 1547 8041
rect 3786 8032 3792 8084
rect 3844 8072 3850 8084
rect 3973 8075 4031 8081
rect 3973 8072 3985 8075
rect 3844 8044 3985 8072
rect 3844 8032 3850 8044
rect 3973 8041 3985 8044
rect 4019 8041 4031 8075
rect 3973 8035 4031 8041
rect 6362 8032 6368 8084
rect 6420 8072 6426 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 6420 8044 6561 8072
rect 6420 8032 6426 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8904 8044 9137 8072
rect 8904 8032 8910 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 10134 8032 10140 8084
rect 10192 8032 10198 8084
rect 10502 8072 10508 8084
rect 10336 8044 10508 8072
rect 106 7964 112 8016
rect 164 8004 170 8016
rect 1857 8007 1915 8013
rect 1857 8004 1869 8007
rect 164 7976 1869 8004
rect 164 7964 170 7976
rect 1857 7973 1869 7976
rect 1903 7973 1915 8007
rect 1857 7967 1915 7973
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 8004 9919 8007
rect 10336 8004 10364 8044
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10870 8032 10876 8084
rect 10928 8032 10934 8084
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 11572 8044 12357 8072
rect 11572 8032 11578 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 13630 8072 13636 8084
rect 12345 8035 12403 8041
rect 12452 8044 13636 8072
rect 9907 7976 10364 8004
rect 10413 8007 10471 8013
rect 9907 7973 9919 7976
rect 9861 7967 9919 7973
rect 10413 7973 10425 8007
rect 10459 7973 10471 8007
rect 10413 7967 10471 7973
rect 11885 8007 11943 8013
rect 11885 7973 11897 8007
rect 11931 8004 11943 8007
rect 11974 8004 11980 8016
rect 11931 7976 11980 8004
rect 11931 7973 11943 7976
rect 11885 7967 11943 7973
rect 8846 7936 8852 7948
rect 1688 7908 8852 7936
rect 1688 7877 1716 7908
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 10428 7936 10456 7967
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 12161 8007 12219 8013
rect 12161 7973 12173 8007
rect 12207 8004 12219 8007
rect 12452 8004 12480 8044
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 14366 8032 14372 8084
rect 14424 8032 14430 8084
rect 15933 8075 15991 8081
rect 15933 8041 15945 8075
rect 15979 8072 15991 8075
rect 16206 8072 16212 8084
rect 15979 8044 16212 8072
rect 15979 8041 15991 8044
rect 15933 8035 15991 8041
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 16482 8032 16488 8084
rect 16540 8032 16546 8084
rect 16942 8032 16948 8084
rect 17000 8032 17006 8084
rect 17221 8075 17279 8081
rect 17221 8041 17233 8075
rect 17267 8072 17279 8075
rect 17402 8072 17408 8084
rect 17267 8044 17408 8072
rect 17267 8041 17279 8044
rect 17221 8035 17279 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 17770 8032 17776 8084
rect 17828 8072 17834 8084
rect 17865 8075 17923 8081
rect 17865 8072 17877 8075
rect 17828 8044 17877 8072
rect 17828 8032 17834 8044
rect 17865 8041 17877 8044
rect 17911 8041 17923 8075
rect 17865 8035 17923 8041
rect 21376 8044 24900 8072
rect 21376 8004 21404 8044
rect 12207 7976 12480 8004
rect 12544 7976 21404 8004
rect 12207 7973 12219 7976
rect 12161 7967 12219 7973
rect 12250 7936 12256 7948
rect 10428 7908 12256 7936
rect 12250 7896 12256 7908
rect 12308 7896 12314 7948
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 2314 7868 2320 7880
rect 2087 7840 2320 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 2406 7828 2412 7880
rect 2464 7828 2470 7880
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 9490 7868 9496 7880
rect 9355 7840 9496 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 3970 7760 3976 7812
rect 4028 7800 4034 7812
rect 5077 7803 5135 7809
rect 5077 7800 5089 7803
rect 4028 7772 5089 7800
rect 4028 7760 4034 7772
rect 5077 7769 5089 7772
rect 5123 7769 5135 7803
rect 5077 7763 5135 7769
rect 5258 7760 5264 7812
rect 5316 7760 5322 7812
rect 6748 7800 6776 7831
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 12544 7877 12572 7976
rect 22002 7964 22008 8016
rect 22060 8004 22066 8016
rect 24872 8004 24900 8044
rect 25222 8032 25228 8084
rect 25280 8032 25286 8084
rect 27617 8075 27675 8081
rect 27617 8072 27629 8075
rect 25332 8044 27629 8072
rect 25332 8004 25360 8044
rect 27617 8041 27629 8044
rect 27663 8041 27675 8075
rect 27617 8035 27675 8041
rect 30101 8075 30159 8081
rect 30101 8041 30113 8075
rect 30147 8072 30159 8075
rect 36630 8072 36636 8084
rect 30147 8044 36636 8072
rect 30147 8041 30159 8044
rect 30101 8035 30159 8041
rect 36630 8032 36636 8044
rect 36688 8032 36694 8084
rect 37826 8032 37832 8084
rect 37884 8072 37890 8084
rect 38013 8075 38071 8081
rect 38013 8072 38025 8075
rect 37884 8044 38025 8072
rect 37884 8032 37890 8044
rect 38013 8041 38025 8044
rect 38059 8041 38071 8075
rect 38013 8035 38071 8041
rect 40034 8032 40040 8084
rect 40092 8032 40098 8084
rect 40770 8032 40776 8084
rect 40828 8032 40834 8084
rect 42334 8032 42340 8084
rect 42392 8032 42398 8084
rect 42702 8032 42708 8084
rect 42760 8032 42766 8084
rect 43441 8075 43499 8081
rect 43441 8041 43453 8075
rect 43487 8072 43499 8075
rect 43530 8072 43536 8084
rect 43487 8044 43536 8072
rect 43487 8041 43499 8044
rect 43441 8035 43499 8041
rect 43530 8032 43536 8044
rect 43588 8032 43594 8084
rect 43714 8032 43720 8084
rect 43772 8072 43778 8084
rect 44177 8075 44235 8081
rect 44177 8072 44189 8075
rect 43772 8044 44189 8072
rect 43772 8032 43778 8044
rect 44177 8041 44189 8044
rect 44223 8041 44235 8075
rect 44177 8035 44235 8041
rect 22060 7976 24808 8004
rect 24872 7976 25360 8004
rect 22060 7964 22066 7976
rect 16574 7936 16580 7948
rect 16546 7896 16580 7936
rect 16632 7896 16638 7948
rect 16758 7896 16764 7948
rect 16816 7936 16822 7948
rect 16816 7908 19288 7936
rect 16816 7896 16822 7908
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7868 9643 7871
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9631 7840 9689 7868
rect 9631 7837 9643 7840
rect 9585 7831 9643 7837
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7868 10195 7871
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 10183 7840 10241 7868
rect 10183 7837 10195 7840
rect 10137 7831 10195 7837
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10873 7871 10931 7877
rect 10873 7837 10885 7871
rect 10919 7868 10931 7871
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 10919 7840 10977 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11931 7840 11989 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 12529 7871 12587 7877
rect 12529 7837 12541 7871
rect 12575 7837 12587 7871
rect 12529 7831 12587 7837
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 12676 7840 14197 7868
rect 12676 7828 12682 7840
rect 14185 7837 14197 7840
rect 14231 7837 14243 7871
rect 14185 7831 14243 7837
rect 15746 7828 15752 7880
rect 15804 7828 15810 7880
rect 16301 7871 16359 7877
rect 16301 7837 16313 7871
rect 16347 7868 16359 7871
rect 16546 7868 16574 7896
rect 16347 7840 16574 7868
rect 16945 7871 17003 7877
rect 16347 7837 16359 7840
rect 16301 7831 16359 7837
rect 16945 7837 16957 7871
rect 16991 7868 17003 7871
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16991 7840 17049 7868
rect 16991 7837 17003 7840
rect 16945 7831 17003 7837
rect 17037 7837 17049 7840
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7868 17831 7871
rect 18046 7868 18052 7880
rect 17819 7840 18052 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 19260 7877 19288 7908
rect 19334 7896 19340 7948
rect 19392 7936 19398 7948
rect 19392 7908 24716 7936
rect 19392 7896 19398 7908
rect 19245 7871 19303 7877
rect 19245 7837 19257 7871
rect 19291 7868 19303 7871
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 19291 7840 19533 7868
rect 19291 7837 19303 7840
rect 19245 7831 19303 7837
rect 19521 7837 19533 7840
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 21637 7871 21695 7877
rect 21637 7837 21649 7871
rect 21683 7868 21695 7871
rect 21729 7871 21787 7877
rect 21729 7868 21741 7871
rect 21683 7840 21741 7868
rect 21683 7837 21695 7840
rect 21637 7831 21695 7837
rect 21729 7837 21741 7840
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 9766 7800 9772 7812
rect 6748 7772 9772 7800
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 13262 7800 13268 7812
rect 11164 7772 13268 7800
rect 842 7692 848 7744
rect 900 7732 906 7744
rect 2225 7735 2283 7741
rect 2225 7732 2237 7735
rect 900 7704 2237 7732
rect 900 7692 906 7704
rect 2225 7701 2237 7704
rect 2271 7701 2283 7735
rect 2225 7695 2283 7701
rect 9585 7735 9643 7741
rect 9585 7701 9597 7735
rect 9631 7732 9643 7735
rect 11054 7732 11060 7744
rect 9631 7704 11060 7732
rect 9631 7701 9643 7704
rect 9585 7695 9643 7701
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 11164 7741 11192 7772
rect 13262 7760 13268 7772
rect 13320 7760 13326 7812
rect 13538 7760 13544 7812
rect 13596 7800 13602 7812
rect 22002 7800 22008 7812
rect 13596 7772 22008 7800
rect 13596 7760 13602 7772
rect 22002 7760 22008 7772
rect 22060 7760 22066 7812
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7701 11207 7735
rect 11149 7695 11207 7701
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 15470 7732 15476 7744
rect 11940 7704 15476 7732
rect 11940 7692 11946 7704
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 19426 7692 19432 7744
rect 19484 7692 19490 7744
rect 21542 7692 21548 7744
rect 21600 7692 21606 7744
rect 21910 7692 21916 7744
rect 21968 7692 21974 7744
rect 24688 7732 24716 7908
rect 24780 7800 24808 7976
rect 25590 7964 25596 8016
rect 25648 7964 25654 8016
rect 25774 7964 25780 8016
rect 25832 8004 25838 8016
rect 26786 8004 26792 8016
rect 25832 7976 26792 8004
rect 25832 7964 25838 7976
rect 26786 7964 26792 7976
rect 26844 7964 26850 8016
rect 26881 8007 26939 8013
rect 26881 7973 26893 8007
rect 26927 7973 26939 8007
rect 26881 7967 26939 7973
rect 25866 7936 25872 7948
rect 25424 7908 25872 7936
rect 25424 7877 25452 7908
rect 25866 7896 25872 7908
rect 25924 7896 25930 7948
rect 26510 7896 26516 7948
rect 26568 7896 26574 7948
rect 25409 7871 25467 7877
rect 25409 7837 25421 7871
rect 25455 7837 25467 7871
rect 25409 7831 25467 7837
rect 25777 7871 25835 7877
rect 25777 7837 25789 7871
rect 25823 7868 25835 7871
rect 26326 7868 26332 7880
rect 25823 7840 26332 7868
rect 25823 7837 25835 7840
rect 25777 7831 25835 7837
rect 26326 7828 26332 7840
rect 26384 7828 26390 7880
rect 26528 7868 26556 7896
rect 26896 7880 26924 7967
rect 26970 7964 26976 8016
rect 27028 7964 27034 8016
rect 28445 8007 28503 8013
rect 28445 8004 28457 8007
rect 27264 7976 28457 8004
rect 26697 7871 26755 7877
rect 26697 7868 26709 7871
rect 26528 7840 26709 7868
rect 26697 7837 26709 7840
rect 26743 7837 26755 7871
rect 26697 7831 26755 7837
rect 26878 7828 26884 7880
rect 26936 7828 26942 7880
rect 27062 7828 27068 7880
rect 27120 7868 27126 7880
rect 27157 7871 27215 7877
rect 27157 7868 27169 7871
rect 27120 7840 27169 7868
rect 27120 7828 27126 7840
rect 27157 7837 27169 7840
rect 27203 7837 27215 7871
rect 27157 7831 27215 7837
rect 27264 7800 27292 7976
rect 28445 7973 28457 7976
rect 28491 7973 28503 8007
rect 28445 7967 28503 7973
rect 36170 7964 36176 8016
rect 36228 8004 36234 8016
rect 36228 7976 40724 8004
rect 36228 7964 36234 7976
rect 33594 7896 33600 7948
rect 33652 7936 33658 7948
rect 33652 7908 38240 7936
rect 33652 7896 33658 7908
rect 27801 7871 27859 7877
rect 27801 7837 27813 7871
rect 27847 7868 27859 7871
rect 28074 7868 28080 7880
rect 27847 7840 28080 7868
rect 27847 7837 27859 7840
rect 27801 7831 27859 7837
rect 28074 7828 28080 7840
rect 28132 7828 28138 7880
rect 28442 7828 28448 7880
rect 28500 7868 28506 7880
rect 28629 7871 28687 7877
rect 28629 7868 28641 7871
rect 28500 7840 28641 7868
rect 28500 7828 28506 7840
rect 28629 7837 28641 7840
rect 28675 7837 28687 7871
rect 28629 7831 28687 7837
rect 29917 7871 29975 7877
rect 29917 7837 29929 7871
rect 29963 7868 29975 7871
rect 33410 7868 33416 7880
rect 29963 7840 33416 7868
rect 29963 7837 29975 7840
rect 29917 7831 29975 7837
rect 33410 7828 33416 7840
rect 33468 7828 33474 7880
rect 33502 7828 33508 7880
rect 33560 7868 33566 7880
rect 38212 7877 38240 7908
rect 36173 7871 36231 7877
rect 36173 7868 36185 7871
rect 33560 7840 36185 7868
rect 33560 7828 33566 7840
rect 36173 7837 36185 7840
rect 36219 7837 36231 7871
rect 36173 7831 36231 7837
rect 38197 7871 38255 7877
rect 38197 7837 38209 7871
rect 38243 7837 38255 7871
rect 38197 7831 38255 7837
rect 39853 7871 39911 7877
rect 39853 7837 39865 7871
rect 39899 7837 39911 7871
rect 39853 7831 39911 7837
rect 24780 7772 27292 7800
rect 35802 7760 35808 7812
rect 35860 7800 35866 7812
rect 35860 7772 36124 7800
rect 35860 7760 35866 7772
rect 35989 7735 36047 7741
rect 35989 7732 36001 7735
rect 24688 7704 36001 7732
rect 35989 7701 36001 7704
rect 36035 7701 36047 7735
rect 36096 7732 36124 7772
rect 39868 7732 39896 7831
rect 40586 7828 40592 7880
rect 40644 7828 40650 7880
rect 40696 7868 40724 7976
rect 41138 7964 41144 8016
rect 41196 8004 41202 8016
rect 43073 8007 43131 8013
rect 41196 7976 43024 8004
rect 41196 7964 41202 7976
rect 40770 7896 40776 7948
rect 40828 7936 40834 7948
rect 40828 7908 42564 7936
rect 40828 7896 40834 7908
rect 41141 7871 41199 7877
rect 41141 7868 41153 7871
rect 40696 7840 41153 7868
rect 41141 7837 41153 7840
rect 41187 7837 41199 7871
rect 41141 7831 41199 7837
rect 41230 7828 41236 7880
rect 41288 7868 41294 7880
rect 41785 7871 41843 7877
rect 41785 7868 41797 7871
rect 41288 7840 41797 7868
rect 41288 7828 41294 7840
rect 41785 7837 41797 7840
rect 41831 7837 41843 7871
rect 41785 7831 41843 7837
rect 42150 7828 42156 7880
rect 42208 7828 42214 7880
rect 42536 7877 42564 7908
rect 42521 7871 42579 7877
rect 42521 7837 42533 7871
rect 42567 7837 42579 7871
rect 42521 7831 42579 7837
rect 42610 7828 42616 7880
rect 42668 7868 42674 7880
rect 42889 7871 42947 7877
rect 42889 7868 42901 7871
rect 42668 7840 42901 7868
rect 42668 7828 42674 7840
rect 42889 7837 42901 7840
rect 42935 7837 42947 7871
rect 42996 7868 43024 7976
rect 43073 7973 43085 8007
rect 43119 8004 43131 8007
rect 43119 7976 43852 8004
rect 43119 7973 43131 7976
rect 43073 7967 43131 7973
rect 43438 7896 43444 7948
rect 43496 7936 43502 7948
rect 43824 7936 43852 7976
rect 44450 7936 44456 7948
rect 43496 7908 43668 7936
rect 43824 7908 44456 7936
rect 43496 7896 43502 7908
rect 43640 7877 43668 7908
rect 44450 7896 44456 7908
rect 44508 7896 44514 7948
rect 43257 7871 43315 7877
rect 43257 7868 43269 7871
rect 42996 7840 43269 7868
rect 42889 7831 42947 7837
rect 43257 7837 43269 7840
rect 43303 7837 43315 7871
rect 43257 7831 43315 7837
rect 43625 7871 43683 7877
rect 43625 7837 43637 7871
rect 43671 7837 43683 7871
rect 43993 7871 44051 7877
rect 43993 7868 44005 7871
rect 43625 7831 43683 7837
rect 43732 7840 44005 7868
rect 43732 7800 43760 7840
rect 43993 7837 44005 7840
rect 44039 7837 44051 7871
rect 43993 7831 44051 7837
rect 44818 7800 44824 7812
rect 41340 7772 43760 7800
rect 43916 7772 44824 7800
rect 41340 7741 41368 7772
rect 36096 7704 39896 7732
rect 41325 7735 41383 7741
rect 35989 7695 36047 7701
rect 41325 7701 41337 7735
rect 41371 7701 41383 7735
rect 41325 7695 41383 7701
rect 41969 7735 42027 7741
rect 41969 7701 41981 7735
rect 42015 7732 42027 7735
rect 42058 7732 42064 7744
rect 42015 7704 42064 7732
rect 42015 7701 42027 7704
rect 41969 7695 42027 7701
rect 42058 7692 42064 7704
rect 42116 7692 42122 7744
rect 43809 7735 43867 7741
rect 43809 7701 43821 7735
rect 43855 7732 43867 7735
rect 43916 7732 43944 7772
rect 44818 7760 44824 7772
rect 44876 7760 44882 7812
rect 43855 7704 43944 7732
rect 43855 7701 43867 7704
rect 43809 7695 43867 7701
rect 1104 7642 44896 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 44896 7642
rect 1104 7568 44896 7590
rect 474 7488 480 7540
rect 532 7528 538 7540
rect 1489 7531 1547 7537
rect 1489 7528 1501 7531
rect 532 7500 1501 7528
rect 532 7488 538 7500
rect 1489 7497 1501 7500
rect 1535 7497 1547 7531
rect 1489 7491 1547 7497
rect 9585 7531 9643 7537
rect 9585 7497 9597 7531
rect 9631 7528 9643 7531
rect 10686 7528 10692 7540
rect 9631 7500 10692 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 12618 7488 12624 7540
rect 12676 7488 12682 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 15378 7528 15384 7540
rect 14783 7500 15384 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 15473 7531 15531 7537
rect 15473 7497 15485 7531
rect 15519 7528 15531 7531
rect 15838 7528 15844 7540
rect 15519 7500 15844 7528
rect 15519 7497 15531 7500
rect 15473 7491 15531 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 17862 7488 17868 7540
rect 17920 7528 17926 7540
rect 21361 7531 21419 7537
rect 21361 7528 21373 7531
rect 17920 7500 21373 7528
rect 17920 7488 17926 7500
rect 21361 7497 21373 7500
rect 21407 7497 21419 7531
rect 21361 7491 21419 7497
rect 26878 7488 26884 7540
rect 26936 7528 26942 7540
rect 36633 7531 36691 7537
rect 26936 7500 36584 7528
rect 26936 7488 26942 7500
rect 12066 7460 12072 7472
rect 2746 7432 12072 7460
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 2746 7392 2774 7432
rect 12066 7420 12072 7432
rect 12124 7420 12130 7472
rect 15197 7463 15255 7469
rect 15197 7429 15209 7463
rect 15243 7460 15255 7463
rect 15654 7460 15660 7472
rect 15243 7432 15660 7460
rect 15243 7429 15255 7432
rect 15197 7423 15255 7429
rect 1719 7364 2774 7392
rect 9401 7395 9459 7401
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 11882 7392 11888 7404
rect 9447 7364 11888 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 12434 7352 12440 7404
rect 12492 7352 12498 7404
rect 13722 7352 13728 7404
rect 13780 7392 13786 7404
rect 14366 7392 14372 7404
rect 13780 7364 14372 7392
rect 13780 7352 13786 7364
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 14550 7352 14556 7404
rect 14608 7352 14614 7404
rect 15304 7401 15332 7432
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 32858 7420 32864 7472
rect 32916 7460 32922 7472
rect 36556 7460 36584 7500
rect 36633 7497 36645 7531
rect 36679 7528 36691 7531
rect 42245 7531 42303 7537
rect 36679 7500 42196 7528
rect 36679 7497 36691 7500
rect 36633 7491 36691 7497
rect 40770 7460 40776 7472
rect 32916 7432 36400 7460
rect 36556 7432 40776 7460
rect 32916 7420 32922 7432
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7392 15347 7395
rect 21545 7395 21603 7401
rect 15335 7364 15369 7392
rect 15335 7361 15347 7364
rect 15289 7355 15347 7361
rect 21545 7361 21557 7395
rect 21591 7392 21603 7395
rect 23290 7392 23296 7404
rect 21591 7364 23296 7392
rect 21591 7361 21603 7364
rect 21545 7355 21603 7361
rect 23290 7352 23296 7364
rect 23348 7352 23354 7404
rect 28445 7395 28503 7401
rect 28445 7361 28457 7395
rect 28491 7392 28503 7395
rect 28810 7392 28816 7404
rect 28491 7364 28816 7392
rect 28491 7361 28503 7364
rect 28445 7355 28503 7361
rect 28810 7352 28816 7364
rect 28868 7352 28874 7404
rect 32398 7352 32404 7404
rect 32456 7392 32462 7404
rect 36372 7401 36400 7432
rect 40770 7420 40776 7432
rect 40828 7420 40834 7472
rect 41874 7420 41880 7472
rect 41932 7420 41938 7472
rect 34517 7395 34575 7401
rect 34517 7392 34529 7395
rect 32456 7364 34529 7392
rect 32456 7352 32462 7364
rect 34517 7361 34529 7364
rect 34563 7361 34575 7395
rect 34517 7355 34575 7361
rect 36357 7395 36415 7401
rect 36357 7361 36369 7395
rect 36403 7361 36415 7395
rect 36357 7355 36415 7361
rect 36446 7352 36452 7404
rect 36504 7352 36510 7404
rect 39850 7352 39856 7404
rect 39908 7392 39914 7404
rect 41049 7395 41107 7401
rect 41049 7392 41061 7395
rect 39908 7364 41061 7392
rect 39908 7352 39914 7364
rect 41049 7361 41061 7364
rect 41095 7361 41107 7395
rect 41892 7392 41920 7420
rect 42061 7395 42119 7401
rect 42061 7392 42073 7395
rect 41892 7364 42073 7392
rect 41049 7355 41107 7361
rect 42061 7361 42073 7364
rect 42107 7361 42119 7395
rect 42168 7392 42196 7500
rect 42245 7497 42257 7531
rect 42291 7528 42303 7531
rect 42610 7528 42616 7540
rect 42291 7500 42616 7528
rect 42291 7497 42303 7500
rect 42245 7491 42303 7497
rect 42610 7488 42616 7500
rect 42668 7488 42674 7540
rect 42978 7488 42984 7540
rect 43036 7488 43042 7540
rect 43346 7488 43352 7540
rect 43404 7488 43410 7540
rect 43717 7531 43775 7537
rect 43717 7497 43729 7531
rect 43763 7528 43775 7531
rect 43806 7528 43812 7540
rect 43763 7500 43812 7528
rect 43763 7497 43775 7500
rect 43717 7491 43775 7497
rect 43806 7488 43812 7500
rect 43864 7488 43870 7540
rect 44085 7531 44143 7537
rect 44085 7497 44097 7531
rect 44131 7528 44143 7531
rect 44358 7528 44364 7540
rect 44131 7500 44364 7528
rect 44131 7497 44143 7500
rect 44085 7491 44143 7497
rect 44358 7488 44364 7500
rect 44416 7488 44422 7540
rect 44450 7488 44456 7540
rect 44508 7488 44514 7540
rect 42426 7392 42432 7404
rect 42168 7364 42432 7392
rect 42061 7355 42119 7361
rect 42426 7352 42432 7364
rect 42484 7352 42490 7404
rect 42521 7395 42579 7401
rect 42521 7361 42533 7395
rect 42567 7361 42579 7395
rect 42521 7355 42579 7361
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 17954 7324 17960 7336
rect 4212 7296 17960 7324
rect 4212 7284 4218 7296
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 18932 7296 36216 7324
rect 18932 7284 18938 7296
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 28261 7259 28319 7265
rect 28261 7256 28273 7259
rect 11020 7228 28273 7256
rect 11020 7216 11026 7228
rect 28261 7225 28273 7228
rect 28307 7225 28319 7259
rect 28261 7219 28319 7225
rect 34330 7216 34336 7268
rect 34388 7216 34394 7268
rect 36188 7265 36216 7296
rect 41966 7284 41972 7336
rect 42024 7324 42030 7336
rect 42536 7324 42564 7355
rect 42794 7352 42800 7404
rect 42852 7352 42858 7404
rect 43162 7352 43168 7404
rect 43220 7352 43226 7404
rect 43254 7352 43260 7404
rect 43312 7392 43318 7404
rect 43533 7395 43591 7401
rect 43533 7392 43545 7395
rect 43312 7364 43545 7392
rect 43312 7352 43318 7364
rect 43533 7361 43545 7364
rect 43579 7361 43591 7395
rect 43533 7355 43591 7361
rect 43901 7395 43959 7401
rect 43901 7361 43913 7395
rect 43947 7361 43959 7395
rect 43901 7355 43959 7361
rect 44269 7395 44327 7401
rect 44269 7361 44281 7395
rect 44315 7392 44327 7395
rect 44358 7392 44364 7404
rect 44315 7364 44364 7392
rect 44315 7361 44327 7364
rect 44269 7355 44327 7361
rect 43806 7324 43812 7336
rect 42024 7296 42564 7324
rect 42720 7296 43812 7324
rect 42024 7284 42030 7296
rect 36173 7259 36231 7265
rect 36173 7225 36185 7259
rect 36219 7225 36231 7259
rect 36173 7219 36231 7225
rect 41230 7216 41236 7268
rect 41288 7216 41294 7268
rect 42610 7256 42616 7268
rect 41340 7228 42616 7256
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 14642 7188 14648 7200
rect 14332 7160 14648 7188
rect 14332 7148 14338 7160
rect 14642 7148 14648 7160
rect 14700 7148 14706 7200
rect 36630 7148 36636 7200
rect 36688 7188 36694 7200
rect 41340 7188 41368 7228
rect 42610 7216 42616 7228
rect 42668 7216 42674 7268
rect 42720 7265 42748 7296
rect 43806 7284 43812 7296
rect 43864 7284 43870 7336
rect 42705 7259 42763 7265
rect 42705 7225 42717 7259
rect 42751 7225 42763 7259
rect 42705 7219 42763 7225
rect 42794 7216 42800 7268
rect 42852 7256 42858 7268
rect 43916 7256 43944 7355
rect 44358 7352 44364 7364
rect 44416 7352 44422 7404
rect 42852 7228 43944 7256
rect 42852 7216 42858 7228
rect 36688 7160 41368 7188
rect 36688 7148 36694 7160
rect 42058 7148 42064 7200
rect 42116 7188 42122 7200
rect 45002 7188 45008 7200
rect 42116 7160 45008 7188
rect 42116 7148 42122 7160
rect 45002 7148 45008 7160
rect 45060 7148 45066 7200
rect 1104 7098 44896 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 43950 7098
rect 44002 7046 44014 7098
rect 44066 7046 44078 7098
rect 44130 7046 44142 7098
rect 44194 7046 44206 7098
rect 44258 7046 44896 7098
rect 1104 7024 44896 7046
rect 2406 6944 2412 6996
rect 2464 6984 2470 6996
rect 11974 6984 11980 6996
rect 2464 6956 11980 6984
rect 2464 6944 2470 6956
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 14366 6984 14372 6996
rect 12406 6956 14372 6984
rect 2314 6876 2320 6928
rect 2372 6916 2378 6928
rect 12406 6916 12434 6956
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 14550 6944 14556 6996
rect 14608 6984 14614 6996
rect 32766 6984 32772 6996
rect 14608 6956 32772 6984
rect 14608 6944 14614 6956
rect 32766 6944 32772 6956
rect 32824 6944 32830 6996
rect 41141 6987 41199 6993
rect 41141 6953 41153 6987
rect 41187 6984 41199 6987
rect 43438 6984 43444 6996
rect 41187 6956 43444 6984
rect 41187 6953 41199 6956
rect 41141 6947 41199 6953
rect 43438 6944 43444 6956
rect 43496 6944 43502 6996
rect 43806 6944 43812 6996
rect 43864 6984 43870 6996
rect 44266 6984 44272 6996
rect 43864 6956 44272 6984
rect 43864 6944 43870 6956
rect 44266 6944 44272 6956
rect 44324 6944 44330 6996
rect 2372 6888 12434 6916
rect 13541 6919 13599 6925
rect 2372 6876 2378 6888
rect 13541 6885 13553 6919
rect 13587 6914 13599 6919
rect 13587 6886 13621 6914
rect 13587 6885 13599 6886
rect 13541 6879 13599 6885
rect 12526 6808 12532 6860
rect 12584 6808 12590 6860
rect 13170 6808 13176 6860
rect 13228 6808 13234 6860
rect 13556 6848 13584 6879
rect 14274 6876 14280 6928
rect 14332 6916 14338 6928
rect 19150 6916 19156 6928
rect 14332 6888 19156 6916
rect 14332 6876 14338 6888
rect 19150 6876 19156 6888
rect 19208 6876 19214 6928
rect 36078 6876 36084 6928
rect 36136 6916 36142 6928
rect 40862 6916 40868 6928
rect 36136 6888 40868 6916
rect 36136 6876 36142 6888
rect 40862 6876 40868 6888
rect 40920 6876 40926 6928
rect 43717 6919 43775 6925
rect 43717 6885 43729 6919
rect 43763 6916 43775 6919
rect 43763 6888 43944 6916
rect 43763 6885 43775 6888
rect 43717 6879 43775 6885
rect 14734 6848 14740 6860
rect 13556 6820 14740 6848
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 14918 6808 14924 6860
rect 14976 6848 14982 6860
rect 34146 6848 34152 6860
rect 14976 6820 34152 6848
rect 14976 6808 14982 6820
rect 34146 6808 34152 6820
rect 34204 6808 34210 6860
rect 43806 6848 43812 6860
rect 42536 6820 43812 6848
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6780 12679 6783
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12667 6752 12725 6780
rect 12667 6749 12679 6752
rect 12621 6743 12679 6749
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 13357 6783 13415 6789
rect 13357 6780 13369 6783
rect 13311 6752 13369 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13357 6749 13369 6752
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 20349 6783 20407 6789
rect 14139 6752 20300 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 5166 6672 5172 6724
rect 5224 6712 5230 6724
rect 5224 6684 20208 6712
rect 5224 6672 5230 6684
rect 12894 6604 12900 6656
rect 12952 6604 12958 6656
rect 14277 6647 14335 6653
rect 14277 6613 14289 6647
rect 14323 6644 14335 6647
rect 14826 6644 14832 6656
rect 14323 6616 14832 6644
rect 14323 6613 14335 6616
rect 14277 6607 14335 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 20180 6653 20208 6684
rect 20165 6647 20223 6653
rect 20165 6613 20177 6647
rect 20211 6613 20223 6647
rect 20272 6644 20300 6752
rect 20349 6749 20361 6783
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6780 22707 6783
rect 23658 6780 23664 6792
rect 22695 6752 23664 6780
rect 22695 6749 22707 6752
rect 22649 6743 22707 6749
rect 20364 6712 20392 6743
rect 23658 6740 23664 6752
rect 23716 6740 23722 6792
rect 25409 6783 25467 6789
rect 25409 6749 25421 6783
rect 25455 6780 25467 6783
rect 25498 6780 25504 6792
rect 25455 6752 25504 6780
rect 25455 6749 25467 6752
rect 25409 6743 25467 6749
rect 25498 6740 25504 6752
rect 25556 6740 25562 6792
rect 37553 6783 37611 6789
rect 37553 6749 37565 6783
rect 37599 6780 37611 6783
rect 37734 6780 37740 6792
rect 37599 6752 37740 6780
rect 37599 6749 37611 6752
rect 37553 6743 37611 6749
rect 37734 6740 37740 6752
rect 37792 6740 37798 6792
rect 40954 6740 40960 6792
rect 41012 6740 41018 6792
rect 42536 6789 42564 6820
rect 43806 6808 43812 6820
rect 43864 6808 43870 6860
rect 43916 6848 43944 6888
rect 45738 6848 45744 6860
rect 43916 6820 45744 6848
rect 45738 6808 45744 6820
rect 45796 6808 45802 6860
rect 42521 6783 42579 6789
rect 42521 6749 42533 6783
rect 42567 6749 42579 6783
rect 42521 6743 42579 6749
rect 42797 6783 42855 6789
rect 42797 6749 42809 6783
rect 42843 6749 42855 6783
rect 42797 6743 42855 6749
rect 22922 6712 22928 6724
rect 20364 6684 22928 6712
rect 22922 6672 22928 6684
rect 22980 6672 22986 6724
rect 25682 6672 25688 6724
rect 25740 6712 25746 6724
rect 42812 6712 42840 6743
rect 43162 6740 43168 6792
rect 43220 6740 43226 6792
rect 43533 6783 43591 6789
rect 43533 6749 43545 6783
rect 43579 6749 43591 6783
rect 43533 6743 43591 6749
rect 43548 6712 43576 6743
rect 43898 6740 43904 6792
rect 43956 6740 43962 6792
rect 43990 6740 43996 6792
rect 44048 6780 44054 6792
rect 44269 6783 44327 6789
rect 44269 6780 44281 6783
rect 44048 6752 44281 6780
rect 44048 6740 44054 6752
rect 44269 6749 44281 6752
rect 44315 6749 44327 6783
rect 44269 6743 44327 6749
rect 25740 6684 42840 6712
rect 42904 6684 43576 6712
rect 25740 6672 25746 6684
rect 22370 6644 22376 6656
rect 20272 6616 22376 6644
rect 20165 6607 20223 6613
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 22462 6604 22468 6656
rect 22520 6604 22526 6656
rect 23382 6604 23388 6656
rect 23440 6644 23446 6656
rect 25225 6647 25283 6653
rect 25225 6644 25237 6647
rect 23440 6616 25237 6644
rect 23440 6604 23446 6616
rect 25225 6613 25237 6616
rect 25271 6613 25283 6647
rect 25225 6607 25283 6613
rect 37737 6647 37795 6653
rect 37737 6613 37749 6647
rect 37783 6644 37795 6647
rect 42150 6644 42156 6656
rect 37783 6616 42156 6644
rect 37783 6613 37795 6616
rect 37737 6607 37795 6613
rect 42150 6604 42156 6616
rect 42208 6604 42214 6656
rect 42705 6647 42763 6653
rect 42705 6613 42717 6647
rect 42751 6644 42763 6647
rect 42904 6644 42932 6684
rect 43622 6672 43628 6724
rect 43680 6712 43686 6724
rect 43680 6684 44128 6712
rect 43680 6672 43686 6684
rect 42751 6616 42932 6644
rect 42751 6613 42763 6616
rect 42705 6607 42763 6613
rect 42978 6604 42984 6656
rect 43036 6604 43042 6656
rect 43346 6604 43352 6656
rect 43404 6604 43410 6656
rect 44100 6653 44128 6684
rect 44085 6647 44143 6653
rect 44085 6613 44097 6647
rect 44131 6613 44143 6647
rect 44085 6607 44143 6613
rect 44450 6604 44456 6656
rect 44508 6604 44514 6656
rect 1104 6554 44896 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 44896 6554
rect 1104 6480 44896 6502
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 14918 6440 14924 6452
rect 9732 6412 14924 6440
rect 9732 6400 9738 6412
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 22925 6443 22983 6449
rect 22925 6440 22937 6443
rect 16546 6412 22937 6440
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 16546 6372 16574 6412
rect 22925 6409 22937 6412
rect 22971 6409 22983 6443
rect 22925 6403 22983 6409
rect 32490 6400 32496 6452
rect 32548 6440 32554 6452
rect 32548 6412 36768 6440
rect 32548 6400 32554 6412
rect 6972 6344 16574 6372
rect 6972 6332 6978 6344
rect 19150 6332 19156 6384
rect 19208 6372 19214 6384
rect 20073 6375 20131 6381
rect 20073 6372 20085 6375
rect 19208 6344 20085 6372
rect 19208 6332 19214 6344
rect 20073 6341 20085 6344
rect 20119 6341 20131 6375
rect 20073 6335 20131 6341
rect 23934 6332 23940 6384
rect 23992 6372 23998 6384
rect 23992 6344 36584 6372
rect 23992 6332 23998 6344
rect 16761 6307 16819 6313
rect 16761 6273 16773 6307
rect 16807 6304 16819 6307
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16807 6276 16865 6304
rect 16807 6273 16819 6276
rect 16761 6267 16819 6273
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 19521 6307 19579 6313
rect 19521 6273 19533 6307
rect 19567 6304 19579 6307
rect 19610 6304 19616 6316
rect 19567 6276 19616 6304
rect 19567 6273 19579 6276
rect 19521 6267 19579 6273
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6304 20223 6307
rect 20257 6307 20315 6313
rect 20257 6304 20269 6307
rect 20211 6276 20269 6304
rect 20211 6273 20223 6276
rect 20165 6267 20223 6273
rect 20257 6273 20269 6276
rect 20303 6273 20315 6307
rect 20257 6267 20315 6273
rect 23109 6307 23167 6313
rect 23109 6273 23121 6307
rect 23155 6304 23167 6307
rect 24026 6304 24032 6316
rect 23155 6276 24032 6304
rect 23155 6273 23167 6276
rect 23109 6267 23167 6273
rect 24026 6264 24032 6276
rect 24084 6264 24090 6316
rect 24670 6264 24676 6316
rect 24728 6304 24734 6316
rect 27065 6307 27123 6313
rect 27065 6304 27077 6307
rect 24728 6276 27077 6304
rect 24728 6264 24734 6276
rect 27065 6273 27077 6276
rect 27111 6304 27123 6307
rect 27341 6307 27399 6313
rect 27341 6304 27353 6307
rect 27111 6276 27353 6304
rect 27111 6273 27123 6276
rect 27065 6267 27123 6273
rect 27341 6273 27353 6276
rect 27387 6273 27399 6307
rect 27341 6267 27399 6273
rect 28353 6307 28411 6313
rect 28353 6273 28365 6307
rect 28399 6304 28411 6307
rect 29178 6304 29184 6316
rect 28399 6276 29184 6304
rect 28399 6273 28411 6276
rect 28353 6267 28411 6273
rect 29178 6264 29184 6276
rect 29236 6264 29242 6316
rect 31754 6264 31760 6316
rect 31812 6304 31818 6316
rect 35161 6307 35219 6313
rect 35161 6304 35173 6307
rect 31812 6276 35173 6304
rect 31812 6264 31818 6276
rect 35161 6273 35173 6276
rect 35207 6273 35219 6307
rect 35161 6267 35219 6273
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 5500 6208 19380 6236
rect 5500 6196 5506 6208
rect 10594 6128 10600 6180
rect 10652 6168 10658 6180
rect 19352 6177 19380 6208
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 34514 6236 34520 6248
rect 20680 6208 34520 6236
rect 20680 6196 20686 6208
rect 34514 6196 34520 6208
rect 34572 6196 34578 6248
rect 34974 6196 34980 6248
rect 35032 6196 35038 6248
rect 36556 6236 36584 6344
rect 36740 6313 36768 6412
rect 44082 6400 44088 6452
rect 44140 6400 44146 6452
rect 44453 6443 44511 6449
rect 44453 6409 44465 6443
rect 44499 6440 44511 6443
rect 45370 6440 45376 6452
rect 44499 6412 45376 6440
rect 44499 6409 44511 6412
rect 44453 6403 44511 6409
rect 45370 6400 45376 6412
rect 45428 6400 45434 6452
rect 42794 6332 42800 6384
rect 42852 6372 42858 6384
rect 43990 6372 43996 6384
rect 42852 6344 43996 6372
rect 42852 6332 42858 6344
rect 43990 6332 43996 6344
rect 44048 6332 44054 6384
rect 36725 6307 36783 6313
rect 36725 6273 36737 6307
rect 36771 6273 36783 6307
rect 36725 6267 36783 6273
rect 43530 6264 43536 6316
rect 43588 6264 43594 6316
rect 43622 6264 43628 6316
rect 43680 6304 43686 6316
rect 43901 6307 43959 6313
rect 43901 6304 43913 6307
rect 43680 6276 43913 6304
rect 43680 6264 43686 6276
rect 43901 6273 43913 6276
rect 43947 6273 43959 6307
rect 43901 6267 43959 6273
rect 44266 6264 44272 6316
rect 44324 6264 44330 6316
rect 44358 6236 44364 6248
rect 36556 6208 44364 6236
rect 44358 6196 44364 6208
rect 44416 6196 44422 6248
rect 19337 6171 19395 6177
rect 10652 6140 19196 6168
rect 10652 6128 10658 6140
rect 16666 6060 16672 6112
rect 16724 6060 16730 6112
rect 17037 6103 17095 6109
rect 17037 6069 17049 6103
rect 17083 6100 17095 6103
rect 19058 6100 19064 6112
rect 17083 6072 19064 6100
rect 17083 6069 17095 6072
rect 17037 6063 17095 6069
rect 19058 6060 19064 6072
rect 19116 6060 19122 6112
rect 19168 6100 19196 6140
rect 19337 6137 19349 6171
rect 19383 6137 19395 6171
rect 28169 6171 28227 6177
rect 28169 6168 28181 6171
rect 19337 6131 19395 6137
rect 19444 6140 28181 6168
rect 19444 6100 19472 6140
rect 28169 6137 28181 6140
rect 28215 6137 28227 6171
rect 28169 6131 28227 6137
rect 34422 6128 34428 6180
rect 34480 6168 34486 6180
rect 43898 6168 43904 6180
rect 34480 6140 43904 6168
rect 34480 6128 34486 6140
rect 43898 6128 43904 6140
rect 43956 6128 43962 6180
rect 19168 6072 19472 6100
rect 20438 6060 20444 6112
rect 20496 6060 20502 6112
rect 27246 6060 27252 6112
rect 27304 6060 27310 6112
rect 29914 6060 29920 6112
rect 29972 6100 29978 6112
rect 34238 6100 34244 6112
rect 29972 6072 34244 6100
rect 29972 6060 29978 6072
rect 34238 6060 34244 6072
rect 34296 6060 34302 6112
rect 34514 6060 34520 6112
rect 34572 6100 34578 6112
rect 36541 6103 36599 6109
rect 36541 6100 36553 6103
rect 34572 6072 36553 6100
rect 34572 6060 34578 6072
rect 36541 6069 36553 6072
rect 36587 6069 36599 6103
rect 36541 6063 36599 6069
rect 43714 6060 43720 6112
rect 43772 6060 43778 6112
rect 1104 6010 44896 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 43950 6010
rect 44002 5958 44014 6010
rect 44066 5958 44078 6010
rect 44130 5958 44142 6010
rect 44194 5958 44206 6010
rect 44258 5958 44896 6010
rect 1104 5936 44896 5958
rect 18601 5899 18659 5905
rect 18601 5896 18613 5899
rect 14844 5868 18613 5896
rect 11238 5788 11244 5840
rect 11296 5828 11302 5840
rect 14844 5828 14872 5868
rect 18601 5865 18613 5868
rect 18647 5865 18659 5899
rect 18601 5859 18659 5865
rect 20438 5856 20444 5908
rect 20496 5896 20502 5908
rect 20496 5868 43944 5896
rect 20496 5856 20502 5868
rect 11296 5800 14872 5828
rect 11296 5788 11302 5800
rect 15010 5788 15016 5840
rect 15068 5828 15074 5840
rect 30561 5831 30619 5837
rect 30561 5828 30573 5831
rect 15068 5800 30573 5828
rect 15068 5788 15074 5800
rect 30561 5797 30573 5800
rect 30607 5797 30619 5831
rect 30561 5791 30619 5797
rect 34146 5788 34152 5840
rect 34204 5788 34210 5840
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 14829 5763 14887 5769
rect 14829 5760 14841 5763
rect 13780 5732 14841 5760
rect 13780 5720 13786 5732
rect 14829 5729 14841 5732
rect 14875 5729 14887 5763
rect 14829 5723 14887 5729
rect 19426 5720 19432 5772
rect 19484 5760 19490 5772
rect 26142 5760 26148 5772
rect 19484 5732 26148 5760
rect 19484 5720 19490 5732
rect 26142 5720 26148 5732
rect 26200 5720 26206 5772
rect 27246 5720 27252 5772
rect 27304 5760 27310 5772
rect 43530 5760 43536 5772
rect 27304 5732 43536 5760
rect 27304 5720 27310 5732
rect 43530 5720 43536 5732
rect 43588 5720 43594 5772
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 18785 5695 18843 5701
rect 5868 5664 16574 5692
rect 5868 5652 5874 5664
rect 14921 5627 14979 5633
rect 14921 5593 14933 5627
rect 14967 5624 14979 5627
rect 15105 5627 15163 5633
rect 15105 5624 15117 5627
rect 14967 5596 15117 5624
rect 14967 5593 14979 5596
rect 14921 5587 14979 5593
rect 15105 5593 15117 5596
rect 15151 5593 15163 5627
rect 15105 5587 15163 5593
rect 15286 5584 15292 5636
rect 15344 5584 15350 5636
rect 16546 5624 16574 5664
rect 18785 5661 18797 5695
rect 18831 5692 18843 5695
rect 22186 5692 22192 5704
rect 18831 5664 22192 5692
rect 18831 5661 18843 5664
rect 18785 5655 18843 5661
rect 22186 5652 22192 5664
rect 22244 5652 22250 5704
rect 25130 5652 25136 5704
rect 25188 5692 25194 5704
rect 25409 5695 25467 5701
rect 25409 5692 25421 5695
rect 25188 5664 25421 5692
rect 25188 5652 25194 5664
rect 25409 5661 25421 5664
rect 25455 5661 25467 5695
rect 25409 5655 25467 5661
rect 29546 5652 29552 5704
rect 29604 5652 29610 5704
rect 29638 5652 29644 5704
rect 29696 5692 29702 5704
rect 29733 5695 29791 5701
rect 29733 5692 29745 5695
rect 29696 5664 29745 5692
rect 29696 5652 29702 5664
rect 29733 5661 29745 5664
rect 29779 5661 29791 5695
rect 29733 5655 29791 5661
rect 30098 5652 30104 5704
rect 30156 5692 30162 5704
rect 30285 5695 30343 5701
rect 30285 5692 30297 5695
rect 30156 5664 30297 5692
rect 30156 5652 30162 5664
rect 30285 5661 30297 5664
rect 30331 5661 30343 5695
rect 30745 5695 30803 5701
rect 30745 5692 30757 5695
rect 30285 5655 30343 5661
rect 30392 5664 30757 5692
rect 29564 5624 29592 5652
rect 30392 5624 30420 5664
rect 30745 5661 30757 5664
rect 30791 5661 30803 5695
rect 30745 5655 30803 5661
rect 31386 5652 31392 5704
rect 31444 5692 31450 5704
rect 43916 5701 43944 5868
rect 44450 5856 44456 5908
rect 44508 5856 44514 5908
rect 34333 5695 34391 5701
rect 34333 5692 34345 5695
rect 31444 5664 34345 5692
rect 31444 5652 31450 5664
rect 34333 5661 34345 5664
rect 34379 5661 34391 5695
rect 34333 5655 34391 5661
rect 43901 5695 43959 5701
rect 43901 5661 43913 5695
rect 43947 5661 43959 5695
rect 43901 5655 43959 5661
rect 44266 5652 44272 5704
rect 44324 5652 44330 5704
rect 43254 5624 43260 5636
rect 16546 5596 25268 5624
rect 29564 5596 30420 5624
rect 30484 5596 43260 5624
rect 7282 5516 7288 5568
rect 7340 5556 7346 5568
rect 22462 5556 22468 5568
rect 7340 5528 22468 5556
rect 7340 5516 7346 5528
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 25240 5565 25268 5596
rect 25225 5559 25283 5565
rect 25225 5525 25237 5559
rect 25271 5525 25283 5559
rect 25225 5519 25283 5525
rect 29914 5516 29920 5568
rect 29972 5516 29978 5568
rect 30484 5565 30512 5596
rect 43254 5584 43260 5596
rect 43312 5584 43318 5636
rect 30469 5559 30527 5565
rect 30469 5525 30481 5559
rect 30515 5525 30527 5559
rect 30469 5519 30527 5525
rect 31018 5516 31024 5568
rect 31076 5556 31082 5568
rect 33502 5556 33508 5568
rect 31076 5528 33508 5556
rect 31076 5516 31082 5528
rect 33502 5516 33508 5528
rect 33560 5516 33566 5568
rect 33594 5516 33600 5568
rect 33652 5556 33658 5568
rect 36170 5556 36176 5568
rect 33652 5528 36176 5556
rect 33652 5516 33658 5528
rect 36170 5516 36176 5528
rect 36228 5516 36234 5568
rect 44085 5559 44143 5565
rect 44085 5525 44097 5559
rect 44131 5556 44143 5559
rect 44358 5556 44364 5568
rect 44131 5528 44364 5556
rect 44131 5525 44143 5528
rect 44085 5519 44143 5525
rect 44358 5516 44364 5528
rect 44416 5516 44422 5568
rect 1104 5466 44896 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 44896 5466
rect 1104 5392 44896 5414
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 23201 5355 23259 5361
rect 23201 5352 23213 5355
rect 9824 5324 23213 5352
rect 9824 5312 9830 5324
rect 23201 5321 23213 5324
rect 23247 5321 23259 5355
rect 31202 5352 31208 5364
rect 23201 5315 23259 5321
rect 23308 5324 31208 5352
rect 19058 5244 19064 5296
rect 19116 5284 19122 5296
rect 23308 5284 23336 5324
rect 31202 5312 31208 5324
rect 31260 5312 31266 5364
rect 33502 5312 33508 5364
rect 33560 5352 33566 5364
rect 33560 5324 44312 5352
rect 33560 5312 33566 5324
rect 24394 5284 24400 5296
rect 19116 5256 23336 5284
rect 23400 5256 24400 5284
rect 19116 5244 19122 5256
rect 20714 5176 20720 5228
rect 20772 5216 20778 5228
rect 23400 5225 23428 5256
rect 24394 5244 24400 5256
rect 24452 5244 24458 5296
rect 26142 5244 26148 5296
rect 26200 5284 26206 5296
rect 31018 5284 31024 5296
rect 26200 5256 31024 5284
rect 26200 5244 26206 5256
rect 31018 5244 31024 5256
rect 31076 5244 31082 5296
rect 31570 5244 31576 5296
rect 31628 5284 31634 5296
rect 31628 5256 31754 5284
rect 31628 5244 31634 5256
rect 22925 5219 22983 5225
rect 22925 5216 22937 5219
rect 20772 5188 22937 5216
rect 20772 5176 20778 5188
rect 22925 5185 22937 5188
rect 22971 5185 22983 5219
rect 22925 5179 22983 5185
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 24213 5219 24271 5225
rect 24213 5185 24225 5219
rect 24259 5216 24271 5219
rect 24762 5216 24768 5228
rect 24259 5188 24768 5216
rect 24259 5185 24271 5188
rect 24213 5179 24271 5185
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 30006 5176 30012 5228
rect 30064 5216 30070 5228
rect 31297 5219 31355 5225
rect 31297 5216 31309 5219
rect 30064 5188 31309 5216
rect 30064 5176 30070 5188
rect 31297 5185 31309 5188
rect 31343 5185 31355 5219
rect 31726 5216 31754 5256
rect 44284 5225 44312 5324
rect 44450 5312 44456 5364
rect 44508 5312 44514 5364
rect 33689 5219 33747 5225
rect 33689 5216 33701 5219
rect 31726 5188 33701 5216
rect 31297 5179 31355 5185
rect 33689 5185 33701 5188
rect 33735 5185 33747 5219
rect 43901 5219 43959 5225
rect 43901 5216 43913 5219
rect 33689 5179 33747 5185
rect 41386 5188 43913 5216
rect 23124 5120 28994 5148
rect 23124 5089 23152 5120
rect 23109 5083 23167 5089
rect 23109 5049 23121 5083
rect 23155 5049 23167 5083
rect 23109 5043 23167 5049
rect 23198 5040 23204 5092
rect 23256 5080 23262 5092
rect 24029 5083 24087 5089
rect 24029 5080 24041 5083
rect 23256 5052 24041 5080
rect 23256 5040 23262 5052
rect 24029 5049 24041 5052
rect 24075 5049 24087 5083
rect 28966 5080 28994 5120
rect 31128 5120 31340 5148
rect 31128 5080 31156 5120
rect 28966 5052 31156 5080
rect 24029 5043 24087 5049
rect 6178 4972 6184 5024
rect 6236 5012 6242 5024
rect 22922 5012 22928 5024
rect 6236 4984 22928 5012
rect 6236 4972 6242 4984
rect 22922 4972 22928 4984
rect 22980 4972 22986 5024
rect 31110 4972 31116 5024
rect 31168 4972 31174 5024
rect 31312 5012 31340 5120
rect 31386 5108 31392 5160
rect 31444 5148 31450 5160
rect 41386 5148 41414 5188
rect 43901 5185 43913 5188
rect 43947 5185 43959 5219
rect 43901 5179 43959 5185
rect 44269 5219 44327 5225
rect 44269 5185 44281 5219
rect 44315 5185 44327 5219
rect 44269 5179 44327 5185
rect 31444 5120 41414 5148
rect 31444 5108 31450 5120
rect 33502 5040 33508 5092
rect 33560 5040 33566 5092
rect 44082 5040 44088 5092
rect 44140 5040 44146 5092
rect 41046 5012 41052 5024
rect 31312 4984 41052 5012
rect 41046 4972 41052 4984
rect 41104 4972 41110 5024
rect 1104 4922 44896 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 43950 4922
rect 44002 4870 44014 4922
rect 44066 4870 44078 4922
rect 44130 4870 44142 4922
rect 44194 4870 44206 4922
rect 44258 4870 44896 4922
rect 1104 4848 44896 4870
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 8386 4808 8392 4820
rect 7708 4780 8392 4808
rect 7708 4768 7714 4780
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 18601 4811 18659 4817
rect 18601 4808 18613 4811
rect 11480 4780 18613 4808
rect 11480 4768 11486 4780
rect 18601 4777 18613 4780
rect 18647 4777 18659 4811
rect 18601 4771 18659 4777
rect 41138 4768 41144 4820
rect 41196 4768 41202 4820
rect 21450 4740 21456 4752
rect 18432 4712 21456 4740
rect 18432 4613 18460 4712
rect 21450 4700 21456 4712
rect 21508 4700 21514 4752
rect 23382 4700 23388 4752
rect 23440 4740 23446 4752
rect 43622 4740 43628 4752
rect 23440 4712 43628 4740
rect 23440 4700 23446 4712
rect 43622 4700 43628 4712
rect 43680 4700 43686 4752
rect 44450 4700 44456 4752
rect 44508 4700 44514 4752
rect 21818 4672 21824 4684
rect 18800 4644 21824 4672
rect 18800 4613 18828 4644
rect 21818 4632 21824 4644
rect 21876 4632 21882 4684
rect 21910 4632 21916 4684
rect 21968 4672 21974 4684
rect 21968 4644 44312 4672
rect 21968 4632 21974 4644
rect 18417 4607 18475 4613
rect 18417 4573 18429 4607
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 18785 4607 18843 4613
rect 18785 4573 18797 4607
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 19797 4607 19855 4613
rect 19797 4604 19809 4607
rect 19751 4576 19809 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 19797 4573 19809 4576
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 30650 4564 30656 4616
rect 30708 4604 30714 4616
rect 33229 4607 33287 4613
rect 33229 4604 33241 4607
rect 30708 4576 33241 4604
rect 30708 4564 30714 4576
rect 33229 4573 33241 4576
rect 33275 4573 33287 4607
rect 33229 4567 33287 4573
rect 39209 4607 39267 4613
rect 39209 4573 39221 4607
rect 39255 4604 39267 4607
rect 39666 4604 39672 4616
rect 39255 4576 39672 4604
rect 39255 4573 39267 4576
rect 39209 4567 39267 4573
rect 39666 4564 39672 4576
rect 39724 4564 39730 4616
rect 40770 4564 40776 4616
rect 40828 4604 40834 4616
rect 40957 4607 41015 4613
rect 40957 4604 40969 4607
rect 40828 4576 40969 4604
rect 40828 4564 40834 4576
rect 40957 4573 40969 4576
rect 41003 4573 41015 4607
rect 40957 4567 41015 4573
rect 41046 4564 41052 4616
rect 41104 4604 41110 4616
rect 44284 4613 44312 4644
rect 43901 4607 43959 4613
rect 43901 4604 43913 4607
rect 41104 4576 43913 4604
rect 41104 4564 41110 4576
rect 43901 4573 43913 4576
rect 43947 4573 43959 4607
rect 43901 4567 43959 4573
rect 44269 4607 44327 4613
rect 44269 4573 44281 4607
rect 44315 4573 44327 4607
rect 44269 4567 44327 4573
rect 9490 4496 9496 4548
rect 9548 4536 9554 4548
rect 42794 4536 42800 4548
rect 9548 4508 22094 4536
rect 9548 4496 9554 4508
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 18233 4471 18291 4477
rect 18233 4468 18245 4471
rect 8352 4440 18245 4468
rect 8352 4428 8358 4440
rect 18233 4437 18245 4440
rect 18279 4437 18291 4471
rect 18233 4431 18291 4437
rect 19610 4428 19616 4480
rect 19668 4428 19674 4480
rect 19978 4428 19984 4480
rect 20036 4428 20042 4480
rect 22066 4468 22094 4508
rect 39408 4508 42800 4536
rect 39408 4477 39436 4508
rect 42794 4496 42800 4508
rect 42852 4496 42858 4548
rect 33045 4471 33103 4477
rect 33045 4468 33057 4471
rect 22066 4440 33057 4468
rect 33045 4437 33057 4440
rect 33091 4437 33103 4471
rect 33045 4431 33103 4437
rect 39393 4471 39451 4477
rect 39393 4437 39405 4471
rect 39439 4437 39451 4471
rect 39393 4431 39451 4437
rect 44082 4428 44088 4480
rect 44140 4428 44146 4480
rect 1104 4378 44896 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 44896 4378
rect 1104 4304 44896 4326
rect 19978 4224 19984 4276
rect 20036 4264 20042 4276
rect 44358 4264 44364 4276
rect 20036 4236 44364 4264
rect 20036 4224 20042 4236
rect 44358 4224 44364 4236
rect 44416 4224 44422 4276
rect 14274 4156 14280 4208
rect 14332 4196 14338 4208
rect 19610 4196 19616 4208
rect 14332 4168 19616 4196
rect 14332 4156 14338 4168
rect 19610 4156 19616 4168
rect 19668 4156 19674 4208
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16393 4131 16451 4137
rect 16393 4128 16405 4131
rect 16356 4100 16405 4128
rect 16356 4088 16362 4100
rect 16393 4097 16405 4100
rect 16439 4097 16451 4131
rect 16393 4091 16451 4097
rect 21913 4131 21971 4137
rect 21913 4097 21925 4131
rect 21959 4128 21971 4131
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21959 4100 22017 4128
rect 21959 4097 21971 4100
rect 21913 4091 21971 4097
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 23385 4131 23443 4137
rect 23385 4097 23397 4131
rect 23431 4128 23443 4131
rect 23477 4131 23535 4137
rect 23477 4128 23489 4131
rect 23431 4100 23489 4128
rect 23431 4097 23443 4100
rect 23385 4091 23443 4097
rect 23477 4097 23489 4100
rect 23523 4097 23535 4131
rect 23477 4091 23535 4097
rect 24305 4131 24363 4137
rect 24305 4097 24317 4131
rect 24351 4128 24363 4131
rect 24397 4131 24455 4137
rect 24397 4128 24409 4131
rect 24351 4100 24409 4128
rect 24351 4097 24363 4100
rect 24305 4091 24363 4097
rect 24397 4097 24409 4100
rect 24443 4097 24455 4131
rect 24397 4091 24455 4097
rect 25685 4131 25743 4137
rect 25685 4097 25697 4131
rect 25731 4128 25743 4131
rect 25777 4131 25835 4137
rect 25777 4128 25789 4131
rect 25731 4100 25789 4128
rect 25731 4097 25743 4100
rect 25685 4091 25743 4097
rect 25777 4097 25789 4100
rect 25823 4097 25835 4131
rect 25777 4091 25835 4097
rect 26878 4088 26884 4140
rect 26936 4128 26942 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 26936 4100 26985 4128
rect 26936 4088 26942 4100
rect 26973 4097 26985 4100
rect 27019 4128 27031 4131
rect 27249 4131 27307 4137
rect 27249 4128 27261 4131
rect 27019 4100 27261 4128
rect 27019 4097 27031 4100
rect 26973 4091 27031 4097
rect 27249 4097 27261 4100
rect 27295 4097 27307 4131
rect 27249 4091 27307 4097
rect 30374 4088 30380 4140
rect 30432 4128 30438 4140
rect 32309 4131 32367 4137
rect 32309 4128 32321 4131
rect 30432 4100 32321 4128
rect 30432 4088 30438 4100
rect 32309 4097 32321 4100
rect 32355 4097 32367 4131
rect 32309 4091 32367 4097
rect 42610 4088 42616 4140
rect 42668 4128 42674 4140
rect 43901 4131 43959 4137
rect 43901 4128 43913 4131
rect 42668 4100 43913 4128
rect 42668 4088 42674 4100
rect 43901 4097 43913 4100
rect 43947 4097 43959 4131
rect 43901 4091 43959 4097
rect 44269 4131 44327 4137
rect 44269 4097 44281 4131
rect 44315 4097 44327 4131
rect 44269 4091 44327 4097
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 9916 4032 26740 4060
rect 9916 4020 9922 4032
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 16209 3995 16267 4001
rect 16209 3992 16221 3995
rect 10376 3964 16221 3992
rect 10376 3952 10382 3964
rect 16209 3961 16221 3964
rect 16255 3961 16267 3995
rect 16209 3955 16267 3961
rect 17678 3952 17684 4004
rect 17736 3992 17742 4004
rect 23382 3992 23388 4004
rect 17736 3964 23388 3992
rect 17736 3952 17742 3964
rect 23382 3952 23388 3964
rect 23440 3952 23446 4004
rect 23658 3952 23664 4004
rect 23716 3952 23722 4004
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 14182 3924 14188 3936
rect 9456 3896 14188 3924
rect 9456 3884 9462 3896
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 17494 3884 17500 3936
rect 17552 3924 17558 3936
rect 18782 3924 18788 3936
rect 17552 3896 18788 3924
rect 17552 3884 17558 3896
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 20496 3896 21833 3924
rect 20496 3884 20502 3896
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 21821 3887 21879 3893
rect 22186 3884 22192 3936
rect 22244 3884 22250 3936
rect 23290 3884 23296 3936
rect 23348 3884 23354 3936
rect 24210 3884 24216 3936
rect 24268 3884 24274 3936
rect 24578 3884 24584 3936
rect 24636 3884 24642 3936
rect 25590 3884 25596 3936
rect 25648 3884 25654 3936
rect 25866 3884 25872 3936
rect 25924 3924 25930 3936
rect 25961 3927 26019 3933
rect 25961 3924 25973 3927
rect 25924 3896 25973 3924
rect 25924 3884 25930 3896
rect 25961 3893 25973 3896
rect 26007 3893 26019 3927
rect 26712 3924 26740 4032
rect 42794 4020 42800 4072
rect 42852 4060 42858 4072
rect 44284 4060 44312 4091
rect 42852 4032 44312 4060
rect 42852 4020 42858 4032
rect 27157 3995 27215 4001
rect 27157 3961 27169 3995
rect 27203 3992 27215 3995
rect 36538 3992 36544 4004
rect 27203 3964 36544 3992
rect 27203 3961 27215 3964
rect 27157 3955 27215 3961
rect 36538 3952 36544 3964
rect 36596 3952 36602 4004
rect 44082 3952 44088 4004
rect 44140 3952 44146 4004
rect 44450 3952 44456 4004
rect 44508 3952 44514 4004
rect 32125 3927 32183 3933
rect 32125 3924 32137 3927
rect 26712 3896 32137 3924
rect 25961 3887 26019 3893
rect 32125 3893 32137 3896
rect 32171 3893 32183 3927
rect 32125 3887 32183 3893
rect 1104 3834 44896 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 43950 3834
rect 44002 3782 44014 3834
rect 44066 3782 44078 3834
rect 44130 3782 44142 3834
rect 44194 3782 44206 3834
rect 44258 3782 44896 3834
rect 1104 3760 44896 3782
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 9217 3723 9275 3729
rect 9217 3720 9229 3723
rect 8904 3692 9229 3720
rect 8904 3680 8910 3692
rect 9217 3689 9229 3692
rect 9263 3689 9275 3723
rect 9217 3683 9275 3689
rect 11974 3680 11980 3732
rect 12032 3680 12038 3732
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 12124 3692 13645 3720
rect 12124 3680 12130 3692
rect 13633 3689 13645 3692
rect 13679 3689 13691 3723
rect 13633 3683 13691 3689
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 14424 3692 14841 3720
rect 14424 3680 14430 3692
rect 14829 3689 14841 3692
rect 14875 3689 14887 3723
rect 14829 3683 14887 3689
rect 17954 3680 17960 3732
rect 18012 3680 18018 3732
rect 20898 3680 20904 3732
rect 20956 3720 20962 3732
rect 27614 3720 27620 3732
rect 20956 3692 27620 3720
rect 20956 3680 20962 3692
rect 27614 3680 27620 3692
rect 27672 3680 27678 3732
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 38562 3652 38568 3664
rect 10008 3624 38568 3652
rect 10008 3612 10014 3624
rect 38562 3612 38568 3624
rect 38620 3612 38626 3664
rect 44450 3612 44456 3664
rect 44508 3612 44514 3664
rect 20990 3584 20996 3596
rect 12406 3556 17632 3584
rect 9398 3476 9404 3528
rect 9456 3476 9462 3528
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 12406 3516 12434 3556
rect 12207 3488 12434 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 13814 3476 13820 3528
rect 13872 3476 13878 3528
rect 15013 3519 15071 3525
rect 15013 3485 15025 3519
rect 15059 3516 15071 3519
rect 17494 3516 17500 3528
rect 15059 3488 17500 3516
rect 15059 3485 15071 3488
rect 15013 3479 15071 3485
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17604 3448 17632 3556
rect 18156 3556 20996 3584
rect 18156 3525 18184 3556
rect 20990 3544 20996 3556
rect 21048 3544 21054 3596
rect 22646 3544 22652 3596
rect 22704 3584 22710 3596
rect 40678 3584 40684 3596
rect 22704 3556 40684 3584
rect 22704 3544 22710 3556
rect 40678 3544 40684 3556
rect 40736 3544 40742 3596
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3516 19671 3519
rect 19705 3519 19763 3525
rect 19705 3516 19717 3519
rect 19659 3488 19717 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 19705 3485 19717 3488
rect 19751 3485 19763 3519
rect 19705 3479 19763 3485
rect 19981 3519 20039 3525
rect 19981 3485 19993 3519
rect 20027 3485 20039 3519
rect 19981 3479 20039 3485
rect 18598 3448 18604 3460
rect 2746 3420 16574 3448
rect 17604 3420 18604 3448
rect 2130 3340 2136 3392
rect 2188 3380 2194 3392
rect 2746 3380 2774 3420
rect 2188 3352 2774 3380
rect 16546 3380 16574 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 18690 3408 18696 3460
rect 18748 3448 18754 3460
rect 19996 3448 20024 3479
rect 20806 3476 20812 3528
rect 20864 3516 20870 3528
rect 22741 3519 22799 3525
rect 22741 3516 22753 3519
rect 20864 3488 22753 3516
rect 20864 3476 20870 3488
rect 22741 3485 22753 3488
rect 22787 3485 22799 3519
rect 33778 3516 33784 3528
rect 22741 3479 22799 3485
rect 28966 3488 33784 3516
rect 28966 3448 28994 3488
rect 33778 3476 33784 3488
rect 33836 3476 33842 3528
rect 36538 3476 36544 3528
rect 36596 3516 36602 3528
rect 43901 3519 43959 3525
rect 43901 3516 43913 3519
rect 36596 3488 43913 3516
rect 36596 3476 36602 3488
rect 43901 3485 43913 3488
rect 43947 3485 43959 3519
rect 43901 3479 43959 3485
rect 44269 3519 44327 3525
rect 44269 3485 44281 3519
rect 44315 3516 44327 3519
rect 44358 3516 44364 3528
rect 44315 3488 44364 3516
rect 44315 3485 44327 3488
rect 44269 3479 44327 3485
rect 44358 3476 44364 3488
rect 44416 3476 44422 3528
rect 31570 3448 31576 3460
rect 18748 3420 20024 3448
rect 20180 3420 28994 3448
rect 31496 3420 31576 3448
rect 18748 3408 18754 3420
rect 19426 3380 19432 3392
rect 16546 3352 19432 3380
rect 2188 3340 2194 3352
rect 19426 3340 19432 3352
rect 19484 3340 19490 3392
rect 19518 3340 19524 3392
rect 19576 3340 19582 3392
rect 19794 3340 19800 3392
rect 19852 3380 19858 3392
rect 20180 3389 20208 3420
rect 19889 3383 19947 3389
rect 19889 3380 19901 3383
rect 19852 3352 19901 3380
rect 19852 3340 19858 3352
rect 19889 3349 19901 3352
rect 19935 3349 19947 3383
rect 19889 3343 19947 3349
rect 20165 3383 20223 3389
rect 20165 3349 20177 3383
rect 20211 3349 20223 3383
rect 20165 3343 20223 3349
rect 20254 3340 20260 3392
rect 20312 3380 20318 3392
rect 22646 3380 22652 3392
rect 20312 3352 22652 3380
rect 20312 3340 20318 3352
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 22925 3383 22983 3389
rect 22925 3349 22937 3383
rect 22971 3380 22983 3383
rect 31496 3380 31524 3420
rect 31570 3408 31576 3420
rect 31628 3408 31634 3460
rect 31754 3408 31760 3460
rect 31812 3448 31818 3460
rect 39942 3448 39948 3460
rect 31812 3420 39948 3448
rect 31812 3408 31818 3420
rect 39942 3408 39948 3420
rect 40000 3408 40006 3460
rect 22971 3352 31524 3380
rect 22971 3349 22983 3352
rect 22925 3343 22983 3349
rect 33778 3340 33784 3392
rect 33836 3380 33842 3392
rect 41690 3380 41696 3392
rect 33836 3352 41696 3380
rect 33836 3340 33842 3352
rect 41690 3340 41696 3352
rect 41748 3340 41754 3392
rect 44082 3340 44088 3392
rect 44140 3340 44146 3392
rect 1104 3290 44896 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 44896 3290
rect 1104 3216 44896 3238
rect 2130 3136 2136 3188
rect 2188 3136 2194 3188
rect 9950 3136 9956 3188
rect 10008 3136 10014 3188
rect 15013 3179 15071 3185
rect 15013 3145 15025 3179
rect 15059 3176 15071 3179
rect 15059 3148 21312 3176
rect 15059 3145 15071 3148
rect 15013 3139 15071 3145
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 10781 3111 10839 3117
rect 10781 3108 10793 3111
rect 9640 3080 10793 3108
rect 9640 3068 9646 3080
rect 10781 3077 10793 3080
rect 10827 3108 10839 3111
rect 11057 3111 11115 3117
rect 11057 3108 11069 3111
rect 10827 3080 11069 3108
rect 10827 3077 10839 3080
rect 10781 3071 10839 3077
rect 11057 3077 11069 3080
rect 11103 3077 11115 3111
rect 11057 3071 11115 3077
rect 11241 3111 11299 3117
rect 11241 3077 11253 3111
rect 11287 3108 11299 3111
rect 16114 3108 16120 3120
rect 11287 3080 16120 3108
rect 11287 3077 11299 3080
rect 11241 3071 11299 3077
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 20898 3108 20904 3120
rect 16224 3080 20904 3108
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 2041 3043 2099 3049
rect 2041 3040 2053 3043
rect 1452 3012 2053 3040
rect 1452 3000 1458 3012
rect 2041 3009 2053 3012
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 7892 3012 8033 3040
rect 7892 3000 7898 3012
rect 8021 3009 8033 3012
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3040 9919 3043
rect 10226 3040 10232 3052
rect 9907 3012 10232 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 12342 3000 12348 3052
rect 12400 3000 12406 3052
rect 14458 3000 14464 3052
rect 14516 3040 14522 3052
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14516 3012 14933 3040
rect 14516 3000 14522 3012
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3040 15899 3043
rect 15933 3043 15991 3049
rect 15933 3040 15945 3043
rect 15887 3012 15945 3040
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 15933 3009 15945 3012
rect 15979 3009 15991 3043
rect 15933 3003 15991 3009
rect 8205 2975 8263 2981
rect 8205 2941 8217 2975
rect 8251 2972 8263 2975
rect 16224 2972 16252 3080
rect 20898 3068 20904 3080
rect 20956 3068 20962 3120
rect 16298 3000 16304 3052
rect 16356 3040 16362 3052
rect 17678 3040 17684 3052
rect 16356 3012 17684 3040
rect 16356 3000 16362 3012
rect 17678 3000 17684 3012
rect 17736 3000 17742 3052
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3040 17831 3043
rect 17865 3043 17923 3049
rect 17865 3040 17877 3043
rect 17819 3012 17877 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 17865 3009 17877 3012
rect 17911 3009 17923 3043
rect 17865 3003 17923 3009
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3009 18199 3043
rect 18141 3003 18199 3009
rect 8251 2944 16252 2972
rect 8251 2941 8263 2944
rect 8205 2935 8263 2941
rect 16574 2932 16580 2984
rect 16632 2972 16638 2984
rect 18156 2972 18184 3003
rect 19702 3000 19708 3052
rect 19760 3040 19766 3052
rect 20073 3043 20131 3049
rect 20073 3040 20085 3043
rect 19760 3012 20085 3040
rect 19760 3000 19766 3012
rect 20073 3009 20085 3012
rect 20119 3040 20131 3043
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 20119 3012 20269 3040
rect 20119 3009 20131 3012
rect 20073 3003 20131 3009
rect 20257 3009 20269 3012
rect 20303 3009 20315 3043
rect 20257 3003 20315 3009
rect 21284 2972 21312 3148
rect 21358 3136 21364 3188
rect 21416 3136 21422 3188
rect 21637 3179 21695 3185
rect 21637 3145 21649 3179
rect 21683 3176 21695 3179
rect 23934 3176 23940 3188
rect 21683 3148 23940 3176
rect 21683 3145 21695 3148
rect 21637 3139 21695 3145
rect 23934 3136 23940 3148
rect 23992 3136 23998 3188
rect 24029 3179 24087 3185
rect 24029 3145 24041 3179
rect 24075 3176 24087 3179
rect 30837 3179 30895 3185
rect 24075 3148 27936 3176
rect 24075 3145 24087 3148
rect 24029 3139 24087 3145
rect 25038 3068 25044 3120
rect 25096 3108 25102 3120
rect 27908 3108 27936 3148
rect 30837 3145 30849 3179
rect 30883 3176 30895 3179
rect 36357 3179 36415 3185
rect 30883 3148 36308 3176
rect 30883 3145 30895 3148
rect 30837 3139 30895 3145
rect 32674 3108 32680 3120
rect 25096 3080 26556 3108
rect 27908 3080 32680 3108
rect 25096 3068 25102 3080
rect 21361 3043 21419 3049
rect 21361 3009 21373 3043
rect 21407 3040 21419 3043
rect 21453 3043 21511 3049
rect 21453 3040 21465 3043
rect 21407 3012 21465 3040
rect 21407 3009 21419 3012
rect 21361 3003 21419 3009
rect 21453 3009 21465 3012
rect 21499 3009 21511 3043
rect 21453 3003 21511 3009
rect 23474 3000 23480 3052
rect 23532 3040 23538 3052
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 23532 3012 23857 3040
rect 23532 3000 23538 3012
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 24210 3000 24216 3052
rect 24268 3040 24274 3052
rect 24397 3043 24455 3049
rect 24397 3040 24409 3043
rect 24268 3012 24409 3040
rect 24268 3000 24274 3012
rect 24397 3009 24409 3012
rect 24443 3009 24455 3043
rect 24397 3003 24455 3009
rect 25498 3000 25504 3052
rect 25556 3000 25562 3052
rect 26528 3049 26556 3080
rect 32674 3068 32680 3080
rect 32732 3068 32738 3120
rect 26513 3043 26571 3049
rect 26513 3009 26525 3043
rect 26559 3009 26571 3043
rect 26513 3003 26571 3009
rect 27801 3043 27859 3049
rect 27801 3009 27813 3043
rect 27847 3040 27859 3043
rect 27893 3043 27951 3049
rect 27893 3040 27905 3043
rect 27847 3012 27905 3040
rect 27847 3009 27859 3012
rect 27801 3003 27859 3009
rect 27893 3009 27905 3012
rect 27939 3009 27951 3043
rect 27893 3003 27951 3009
rect 29270 3000 29276 3052
rect 29328 3040 29334 3052
rect 30653 3043 30711 3049
rect 30653 3040 30665 3043
rect 29328 3012 30665 3040
rect 29328 3000 29334 3012
rect 30653 3009 30665 3012
rect 30699 3009 30711 3043
rect 30653 3003 30711 3009
rect 36170 3000 36176 3052
rect 36228 3000 36234 3052
rect 36078 2972 36084 2984
rect 16632 2944 18184 2972
rect 18248 2944 18460 2972
rect 21284 2944 36084 2972
rect 16632 2932 16638 2944
rect 12529 2907 12587 2913
rect 12529 2873 12541 2907
rect 12575 2904 12587 2907
rect 18248 2904 18276 2944
rect 12575 2876 18276 2904
rect 18432 2904 18460 2944
rect 36078 2932 36084 2944
rect 36136 2932 36142 2984
rect 36280 2972 36308 3148
rect 36357 3145 36369 3179
rect 36403 3176 36415 3179
rect 37274 3176 37280 3188
rect 36403 3148 37280 3176
rect 36403 3145 36415 3148
rect 36357 3139 36415 3145
rect 37274 3136 37280 3148
rect 37332 3136 37338 3188
rect 38286 3136 38292 3188
rect 38344 3136 38350 3188
rect 42886 3136 42892 3188
rect 42944 3176 42950 3188
rect 42944 3148 44312 3176
rect 42944 3136 42950 3148
rect 40034 3068 40040 3120
rect 40092 3108 40098 3120
rect 40092 3080 43944 3108
rect 40092 3068 40098 3080
rect 37274 3000 37280 3052
rect 37332 3000 37338 3052
rect 37366 3000 37372 3052
rect 37424 3040 37430 3052
rect 38105 3043 38163 3049
rect 38105 3040 38117 3043
rect 37424 3012 38117 3040
rect 37424 3000 37430 3012
rect 38105 3009 38117 3012
rect 38151 3009 38163 3043
rect 38105 3003 38163 3009
rect 40126 3000 40132 3052
rect 40184 3040 40190 3052
rect 43916 3049 43944 3080
rect 44284 3049 44312 3148
rect 44450 3136 44456 3188
rect 44508 3136 44514 3188
rect 43533 3043 43591 3049
rect 43533 3040 43545 3043
rect 40184 3012 43545 3040
rect 40184 3000 40190 3012
rect 43533 3009 43545 3012
rect 43579 3009 43591 3043
rect 43533 3003 43591 3009
rect 43901 3043 43959 3049
rect 43901 3009 43913 3043
rect 43947 3009 43959 3043
rect 43901 3003 43959 3009
rect 44269 3043 44327 3049
rect 44269 3009 44281 3043
rect 44315 3009 44327 3043
rect 44269 3003 44327 3009
rect 43070 2972 43076 2984
rect 36280 2944 43076 2972
rect 43070 2932 43076 2944
rect 43128 2932 43134 2984
rect 35710 2904 35716 2916
rect 18432 2876 35716 2904
rect 12575 2873 12587 2876
rect 12529 2867 12587 2873
rect 35710 2864 35716 2876
rect 35768 2864 35774 2916
rect 37461 2907 37519 2913
rect 37461 2873 37473 2907
rect 37507 2904 37519 2907
rect 38378 2904 38384 2916
rect 37507 2876 38384 2904
rect 37507 2873 37519 2876
rect 37461 2867 37519 2873
rect 38378 2864 38384 2876
rect 38436 2864 38442 2916
rect 44082 2864 44088 2916
rect 44140 2864 44146 2916
rect 15746 2796 15752 2848
rect 15804 2796 15810 2848
rect 16114 2796 16120 2848
rect 16172 2796 16178 2848
rect 17678 2796 17684 2848
rect 17736 2796 17742 2848
rect 18046 2796 18052 2848
rect 18104 2796 18110 2848
rect 18325 2839 18383 2845
rect 18325 2805 18337 2839
rect 18371 2836 18383 2839
rect 20254 2836 20260 2848
rect 18371 2808 20260 2836
rect 18371 2805 18383 2808
rect 18325 2799 18383 2805
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 20441 2839 20499 2845
rect 20441 2805 20453 2839
rect 20487 2836 20499 2839
rect 20530 2836 20536 2848
rect 20487 2808 20536 2836
rect 20487 2805 20499 2808
rect 20441 2799 20499 2805
rect 20530 2796 20536 2808
rect 20588 2796 20594 2848
rect 24581 2839 24639 2845
rect 24581 2805 24593 2839
rect 24627 2836 24639 2839
rect 24854 2836 24860 2848
rect 24627 2808 24860 2836
rect 24627 2805 24639 2808
rect 24581 2799 24639 2805
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 25682 2796 25688 2848
rect 25740 2796 25746 2848
rect 26694 2796 26700 2848
rect 26752 2796 26758 2848
rect 27706 2796 27712 2848
rect 27764 2796 27770 2848
rect 28077 2839 28135 2845
rect 28077 2805 28089 2839
rect 28123 2836 28135 2839
rect 30282 2836 30288 2848
rect 28123 2808 30288 2836
rect 28123 2805 28135 2808
rect 28077 2799 28135 2805
rect 30282 2796 30288 2808
rect 30340 2796 30346 2848
rect 43717 2839 43775 2845
rect 43717 2805 43729 2839
rect 43763 2836 43775 2839
rect 44818 2836 44824 2848
rect 43763 2808 44824 2836
rect 43763 2805 43775 2808
rect 43717 2799 43775 2805
rect 44818 2796 44824 2808
rect 44876 2796 44882 2848
rect 1104 2746 44896 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 43950 2746
rect 44002 2694 44014 2746
rect 44066 2694 44078 2746
rect 44130 2694 44142 2746
rect 44194 2694 44206 2746
rect 44258 2694 44896 2746
rect 1104 2672 44896 2694
rect 19426 2592 19432 2644
rect 19484 2632 19490 2644
rect 43530 2632 43536 2644
rect 19484 2604 43536 2632
rect 19484 2592 19490 2604
rect 43530 2592 43536 2604
rect 43588 2592 43594 2644
rect 19794 2524 19800 2576
rect 19852 2564 19858 2576
rect 36722 2564 36728 2576
rect 19852 2536 36728 2564
rect 19852 2524 19858 2536
rect 36722 2524 36728 2536
rect 36780 2524 36786 2576
rect 36998 2524 37004 2576
rect 37056 2564 37062 2576
rect 37056 2536 42932 2564
rect 37056 2524 37062 2536
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18104 2468 33824 2496
rect 18104 2456 18110 2468
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 33796 2428 33824 2468
rect 36906 2456 36912 2508
rect 36964 2496 36970 2508
rect 42904 2496 42932 2536
rect 42978 2524 42984 2576
rect 43036 2524 43042 2576
rect 43717 2567 43775 2573
rect 43717 2533 43729 2567
rect 43763 2564 43775 2567
rect 44358 2564 44364 2576
rect 43763 2536 44364 2564
rect 43763 2533 43775 2536
rect 43717 2527 43775 2533
rect 44358 2524 44364 2536
rect 44416 2524 44422 2576
rect 44450 2524 44456 2576
rect 44508 2524 44514 2576
rect 36964 2468 42840 2496
rect 42904 2468 43944 2496
rect 36964 2456 36970 2468
rect 36998 2428 37004 2440
rect 16172 2400 31754 2428
rect 33796 2400 37004 2428
rect 16172 2388 16178 2400
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 26878 2360 26884 2372
rect 12492 2332 26884 2360
rect 12492 2320 12498 2332
rect 26878 2320 26884 2332
rect 26936 2320 26942 2372
rect 31726 2360 31754 2400
rect 36998 2388 37004 2400
rect 37056 2388 37062 2440
rect 42812 2437 42840 2468
rect 42803 2431 42861 2437
rect 42803 2397 42815 2431
rect 42849 2397 42861 2431
rect 42803 2391 42861 2397
rect 43165 2431 43223 2437
rect 43165 2397 43177 2431
rect 43211 2397 43223 2431
rect 43165 2391 43223 2397
rect 43180 2360 43208 2391
rect 43530 2388 43536 2440
rect 43588 2388 43594 2440
rect 43916 2437 43944 2468
rect 43901 2431 43959 2437
rect 43901 2397 43913 2431
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 44269 2431 44327 2437
rect 44269 2397 44281 2431
rect 44315 2397 44327 2431
rect 44269 2391 44327 2397
rect 44284 2360 44312 2391
rect 31726 2332 43208 2360
rect 43272 2332 44312 2360
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 25498 2292 25504 2304
rect 5592 2264 25504 2292
rect 5592 2252 5598 2264
rect 25498 2252 25504 2264
rect 25556 2252 25562 2304
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 43272 2292 43300 2332
rect 30340 2264 43300 2292
rect 30340 2252 30346 2264
rect 43346 2252 43352 2304
rect 43404 2252 43410 2304
rect 44082 2252 44088 2304
rect 44140 2252 44146 2304
rect 1104 2202 44896 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 44896 2202
rect 1104 2128 44896 2150
rect 31386 212 31392 264
rect 31444 252 31450 264
rect 40586 252 40592 264
rect 31444 224 40592 252
rect 31444 212 31450 224
rect 40586 212 40592 224
rect 40644 212 40650 264
rect 3878 144 3884 196
rect 3936 144 3942 196
rect 5994 144 6000 196
rect 6052 184 6058 196
rect 37366 184 37372 196
rect 6052 156 37372 184
rect 6052 144 6058 156
rect 37366 144 37372 156
rect 37424 144 37430 196
rect 3896 116 3924 144
rect 37274 116 37280 128
rect 3896 88 37280 116
rect 37274 76 37280 88
rect 37332 76 37338 128
rect 1854 8 1860 60
rect 1912 48 1918 60
rect 36170 48 36176 60
rect 1912 20 36176 48
rect 1912 8 1918 20
rect 36170 8 36176 20
rect 36228 8 36234 60
<< via1 >>
rect 16580 11092 16632 11144
rect 34612 11092 34664 11144
rect 18052 11024 18104 11076
rect 33876 11024 33928 11076
rect 16396 10956 16448 11008
rect 20720 10956 20772 11008
rect 21364 10956 21416 11008
rect 37280 10956 37332 11008
rect 15476 10888 15528 10940
rect 27712 10888 27764 10940
rect 18788 10752 18840 10804
rect 20352 10752 20404 10804
rect 37188 10004 37240 10056
rect 38016 10004 38068 10056
rect 18604 9664 18656 9716
rect 19616 9664 19668 9716
rect 1124 9392 1176 9444
rect 40960 9392 41012 9444
rect 1032 9324 1084 9376
rect 39672 9324 39724 9376
rect 9864 9256 9916 9308
rect 31116 9256 31168 9308
rect 4344 9188 4396 9240
rect 10324 9188 10376 9240
rect 16948 9188 17000 9240
rect 34336 9188 34388 9240
rect 12440 9120 12492 9172
rect 21364 9120 21416 9172
rect 27620 9120 27672 9172
rect 39580 9120 39632 9172
rect 3608 9052 3660 9104
rect 8300 9052 8352 9104
rect 1768 8984 1820 9036
rect 10232 8984 10284 9036
rect 17868 9052 17920 9104
rect 19616 9052 19668 9104
rect 22560 9052 22612 9104
rect 32680 9052 32732 9104
rect 42800 9052 42852 9104
rect 10876 8984 10928 9036
rect 2504 8848 2556 8900
rect 5448 8848 5500 8900
rect 10508 8916 10560 8968
rect 14280 8916 14332 8968
rect 15660 8984 15712 9036
rect 35440 8984 35492 9036
rect 37188 8916 37240 8968
rect 40776 8916 40828 8968
rect 43996 8916 44048 8968
rect 36452 8848 36504 8900
rect 40040 8848 40092 8900
rect 43536 8848 43588 8900
rect 3516 8780 3568 8832
rect 11244 8780 11296 8832
rect 11336 8780 11388 8832
rect 13544 8780 13596 8832
rect 33784 8780 33836 8832
rect 42892 8780 42944 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 2872 8576 2924 8628
rect 3424 8619 3476 8628
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 4160 8619 4212 8628
rect 4160 8585 4169 8619
rect 4169 8585 4203 8619
rect 4203 8585 4212 8619
rect 4160 8576 4212 8585
rect 4528 8619 4580 8628
rect 4528 8585 4537 8619
rect 4537 8585 4571 8619
rect 4571 8585 4580 8619
rect 4528 8576 4580 8585
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 6000 8619 6052 8628
rect 6000 8585 6009 8619
rect 6009 8585 6043 8619
rect 6043 8585 6052 8619
rect 6000 8576 6052 8585
rect 6736 8619 6788 8628
rect 6736 8585 6745 8619
rect 6745 8585 6779 8619
rect 6779 8585 6788 8619
rect 6736 8576 6788 8585
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 7472 8619 7524 8628
rect 7472 8585 7481 8619
rect 7481 8585 7515 8619
rect 7515 8585 7524 8619
rect 7472 8576 7524 8585
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 11244 8576 11296 8628
rect 11888 8576 11940 8628
rect 12256 8576 12308 8628
rect 12624 8576 12676 8628
rect 12992 8619 13044 8628
rect 12992 8585 13001 8619
rect 13001 8585 13035 8619
rect 13035 8585 13044 8619
rect 12992 8576 13044 8585
rect 13360 8576 13412 8628
rect 13728 8576 13780 8628
rect 14464 8576 14516 8628
rect 14832 8576 14884 8628
rect 15384 8576 15436 8628
rect 15568 8576 15620 8628
rect 15936 8576 15988 8628
rect 16304 8576 16356 8628
rect 16672 8576 16724 8628
rect 17040 8576 17092 8628
rect 17408 8576 17460 8628
rect 17776 8576 17828 8628
rect 18144 8576 18196 8628
rect 18512 8576 18564 8628
rect 18880 8576 18932 8628
rect 38384 8576 38436 8628
rect 38568 8576 38620 8628
rect 38660 8576 38712 8628
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 3516 8440 3568 8492
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 5172 8372 5224 8424
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 7840 8440 7892 8492
rect 9588 8508 9640 8560
rect 9404 8440 9456 8492
rect 9680 8440 9732 8492
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10508 8440 10560 8492
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 10692 8372 10744 8424
rect 10232 8304 10284 8356
rect 10508 8304 10560 8356
rect 12256 8440 12308 8492
rect 25780 8508 25832 8560
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 13268 8440 13320 8449
rect 13636 8483 13688 8492
rect 13636 8449 13645 8483
rect 13645 8449 13679 8483
rect 13679 8449 13688 8483
rect 13636 8440 13688 8449
rect 13728 8440 13780 8492
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 14832 8440 14884 8492
rect 15384 8440 15436 8492
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16212 8483 16264 8492
rect 16212 8449 16221 8483
rect 16221 8449 16255 8483
rect 16255 8449 16264 8483
rect 16212 8440 16264 8449
rect 16488 8440 16540 8492
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 20628 8440 20680 8492
rect 37280 8440 37332 8492
rect 12900 8304 12952 8356
rect 13728 8304 13780 8356
rect 19248 8372 19300 8424
rect 26700 8372 26752 8424
rect 33784 8372 33836 8424
rect 38292 8372 38344 8424
rect 39028 8619 39080 8628
rect 39028 8585 39037 8619
rect 39037 8585 39071 8619
rect 39071 8585 39080 8619
rect 39028 8576 39080 8585
rect 39396 8619 39448 8628
rect 39396 8585 39405 8619
rect 39405 8585 39439 8619
rect 39439 8585 39448 8619
rect 39396 8576 39448 8585
rect 39488 8576 39540 8628
rect 40224 8576 40276 8628
rect 40868 8576 40920 8628
rect 41236 8576 41288 8628
rect 41696 8576 41748 8628
rect 43260 8576 43312 8628
rect 43628 8508 43680 8560
rect 38844 8449 38875 8476
rect 38875 8449 38896 8476
rect 38844 8424 38896 8449
rect 39580 8440 39632 8492
rect 40224 8483 40276 8492
rect 40224 8449 40233 8483
rect 40233 8449 40267 8483
rect 40267 8449 40276 8483
rect 40224 8440 40276 8449
rect 40868 8440 40920 8492
rect 23388 8304 23440 8356
rect 35716 8304 35768 8356
rect 8576 8279 8628 8288
rect 8576 8245 8585 8279
rect 8585 8245 8619 8279
rect 8619 8245 8628 8279
rect 8576 8236 8628 8245
rect 9312 8279 9364 8288
rect 9312 8245 9321 8279
rect 9321 8245 9355 8279
rect 9355 8245 9364 8279
rect 9312 8236 9364 8245
rect 9496 8236 9548 8288
rect 9956 8236 10008 8288
rect 10416 8279 10468 8288
rect 10416 8245 10425 8279
rect 10425 8245 10459 8279
rect 10459 8245 10468 8279
rect 10416 8236 10468 8245
rect 10784 8279 10836 8288
rect 10784 8245 10793 8279
rect 10793 8245 10827 8279
rect 10827 8245 10836 8279
rect 10784 8236 10836 8245
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 18144 8236 18196 8288
rect 37832 8236 37884 8288
rect 38384 8304 38436 8356
rect 38660 8304 38712 8356
rect 40684 8372 40736 8424
rect 41696 8483 41748 8492
rect 41696 8449 41705 8483
rect 41705 8449 41739 8483
rect 41739 8449 41748 8483
rect 41696 8440 41748 8449
rect 42800 8483 42852 8492
rect 42800 8449 42809 8483
rect 42809 8449 42843 8483
rect 42843 8449 42852 8483
rect 42800 8440 42852 8449
rect 42892 8440 42944 8492
rect 43260 8440 43312 8492
rect 39856 8304 39908 8356
rect 42524 8372 42576 8424
rect 43536 8483 43588 8492
rect 43536 8449 43545 8483
rect 43545 8449 43579 8483
rect 43579 8449 43588 8483
rect 43536 8440 43588 8449
rect 43996 8440 44048 8492
rect 39948 8236 40000 8288
rect 41328 8304 41380 8356
rect 42064 8304 42116 8356
rect 43444 8304 43496 8356
rect 42340 8236 42392 8288
rect 44640 8236 44692 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 43950 8134 44002 8186
rect 44014 8134 44066 8186
rect 44078 8134 44130 8186
rect 44142 8134 44194 8186
rect 44206 8134 44258 8186
rect 1216 8032 1268 8084
rect 3792 8032 3844 8084
rect 6368 8032 6420 8084
rect 8852 8032 8904 8084
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 112 7964 164 8016
rect 10508 8032 10560 8084
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 11520 8032 11572 8084
rect 8852 7896 8904 7948
rect 11980 7964 12032 8016
rect 13636 8032 13688 8084
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 16212 8032 16264 8084
rect 16488 8075 16540 8084
rect 16488 8041 16497 8075
rect 16497 8041 16531 8075
rect 16531 8041 16540 8075
rect 16488 8032 16540 8041
rect 16948 8075 17000 8084
rect 16948 8041 16957 8075
rect 16957 8041 16991 8075
rect 16991 8041 17000 8075
rect 16948 8032 17000 8041
rect 17408 8032 17460 8084
rect 17776 8032 17828 8084
rect 12256 7896 12308 7948
rect 2320 7828 2372 7880
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 3976 7760 4028 7812
rect 5264 7803 5316 7812
rect 5264 7769 5273 7803
rect 5273 7769 5307 7803
rect 5307 7769 5316 7803
rect 5264 7760 5316 7769
rect 9496 7828 9548 7880
rect 22008 7964 22060 8016
rect 25228 8075 25280 8084
rect 25228 8041 25237 8075
rect 25237 8041 25271 8075
rect 25271 8041 25280 8075
rect 25228 8032 25280 8041
rect 36636 8032 36688 8084
rect 37832 8032 37884 8084
rect 40040 8075 40092 8084
rect 40040 8041 40049 8075
rect 40049 8041 40083 8075
rect 40083 8041 40092 8075
rect 40040 8032 40092 8041
rect 40776 8075 40828 8084
rect 40776 8041 40785 8075
rect 40785 8041 40819 8075
rect 40819 8041 40828 8075
rect 40776 8032 40828 8041
rect 42340 8075 42392 8084
rect 42340 8041 42349 8075
rect 42349 8041 42383 8075
rect 42383 8041 42392 8075
rect 42340 8032 42392 8041
rect 42708 8075 42760 8084
rect 42708 8041 42717 8075
rect 42717 8041 42751 8075
rect 42751 8041 42760 8075
rect 42708 8032 42760 8041
rect 43536 8032 43588 8084
rect 43720 8032 43772 8084
rect 16580 7896 16632 7948
rect 16764 7896 16816 7948
rect 12624 7828 12676 7880
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 19340 7896 19392 7948
rect 9772 7760 9824 7812
rect 848 7692 900 7744
rect 11060 7692 11112 7744
rect 13268 7760 13320 7812
rect 13544 7760 13596 7812
rect 22008 7760 22060 7812
rect 11888 7692 11940 7744
rect 15476 7692 15528 7744
rect 19432 7735 19484 7744
rect 19432 7701 19441 7735
rect 19441 7701 19475 7735
rect 19475 7701 19484 7735
rect 19432 7692 19484 7701
rect 21548 7735 21600 7744
rect 21548 7701 21557 7735
rect 21557 7701 21591 7735
rect 21591 7701 21600 7735
rect 21548 7692 21600 7701
rect 21916 7735 21968 7744
rect 21916 7701 21925 7735
rect 21925 7701 21959 7735
rect 21959 7701 21968 7735
rect 21916 7692 21968 7701
rect 25596 8007 25648 8016
rect 25596 7973 25605 8007
rect 25605 7973 25639 8007
rect 25639 7973 25648 8007
rect 25596 7964 25648 7973
rect 25780 7964 25832 8016
rect 26792 7964 26844 8016
rect 25872 7896 25924 7948
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 26332 7828 26384 7880
rect 26976 8007 27028 8016
rect 26976 7973 26985 8007
rect 26985 7973 27019 8007
rect 27019 7973 27028 8007
rect 26976 7964 27028 7973
rect 26884 7828 26936 7880
rect 27068 7828 27120 7880
rect 36176 7964 36228 8016
rect 33600 7896 33652 7948
rect 28080 7828 28132 7880
rect 28448 7828 28500 7880
rect 33416 7828 33468 7880
rect 33508 7828 33560 7880
rect 35808 7760 35860 7812
rect 40592 7871 40644 7880
rect 40592 7837 40601 7871
rect 40601 7837 40635 7871
rect 40635 7837 40644 7871
rect 40592 7828 40644 7837
rect 41144 7964 41196 8016
rect 40776 7896 40828 7948
rect 41236 7828 41288 7880
rect 42156 7871 42208 7880
rect 42156 7837 42165 7871
rect 42165 7837 42199 7871
rect 42199 7837 42208 7871
rect 42156 7828 42208 7837
rect 42616 7828 42668 7880
rect 43444 7896 43496 7948
rect 44456 7896 44508 7948
rect 42064 7692 42116 7744
rect 44824 7760 44876 7812
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 480 7488 532 7540
rect 10692 7488 10744 7540
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 15384 7488 15436 7540
rect 15844 7488 15896 7540
rect 17868 7488 17920 7540
rect 26884 7488 26936 7540
rect 12072 7420 12124 7472
rect 11888 7352 11940 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 13728 7352 13780 7404
rect 14372 7352 14424 7404
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 15660 7420 15712 7472
rect 32864 7420 32916 7472
rect 23296 7352 23348 7404
rect 28816 7352 28868 7404
rect 32404 7352 32456 7404
rect 40776 7420 40828 7472
rect 41880 7463 41932 7472
rect 41880 7429 41889 7463
rect 41889 7429 41923 7463
rect 41923 7429 41932 7463
rect 41880 7420 41932 7429
rect 36452 7395 36504 7404
rect 36452 7361 36461 7395
rect 36461 7361 36495 7395
rect 36495 7361 36504 7395
rect 36452 7352 36504 7361
rect 39856 7352 39908 7404
rect 42616 7488 42668 7540
rect 42984 7531 43036 7540
rect 42984 7497 42993 7531
rect 42993 7497 43027 7531
rect 43027 7497 43036 7531
rect 42984 7488 43036 7497
rect 43352 7531 43404 7540
rect 43352 7497 43361 7531
rect 43361 7497 43395 7531
rect 43395 7497 43404 7531
rect 43352 7488 43404 7497
rect 43812 7488 43864 7540
rect 44364 7488 44416 7540
rect 44456 7531 44508 7540
rect 44456 7497 44465 7531
rect 44465 7497 44499 7531
rect 44499 7497 44508 7531
rect 44456 7488 44508 7497
rect 42432 7352 42484 7404
rect 4160 7284 4212 7336
rect 17960 7284 18012 7336
rect 18880 7284 18932 7336
rect 10968 7216 11020 7268
rect 34336 7259 34388 7268
rect 34336 7225 34345 7259
rect 34345 7225 34379 7259
rect 34379 7225 34388 7259
rect 34336 7216 34388 7225
rect 41972 7284 42024 7336
rect 42800 7395 42852 7404
rect 42800 7361 42809 7395
rect 42809 7361 42843 7395
rect 42843 7361 42852 7395
rect 42800 7352 42852 7361
rect 43168 7395 43220 7404
rect 43168 7361 43177 7395
rect 43177 7361 43211 7395
rect 43211 7361 43220 7395
rect 43168 7352 43220 7361
rect 43260 7352 43312 7404
rect 41236 7259 41288 7268
rect 41236 7225 41245 7259
rect 41245 7225 41279 7259
rect 41279 7225 41288 7259
rect 41236 7216 41288 7225
rect 14280 7148 14332 7200
rect 14648 7148 14700 7200
rect 36636 7148 36688 7200
rect 42616 7216 42668 7268
rect 43812 7284 43864 7336
rect 42800 7216 42852 7268
rect 44364 7352 44416 7404
rect 42064 7148 42116 7200
rect 45008 7148 45060 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 43950 7046 44002 7098
rect 44014 7046 44066 7098
rect 44078 7046 44130 7098
rect 44142 7046 44194 7098
rect 44206 7046 44258 7098
rect 2412 6944 2464 6996
rect 11980 6944 12032 6996
rect 2320 6876 2372 6928
rect 14372 6944 14424 6996
rect 14556 6944 14608 6996
rect 32772 6944 32824 6996
rect 43444 6944 43496 6996
rect 43812 6944 43864 6996
rect 44272 6944 44324 6996
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 13176 6851 13228 6860
rect 13176 6817 13185 6851
rect 13185 6817 13219 6851
rect 13219 6817 13228 6851
rect 13176 6808 13228 6817
rect 14280 6876 14332 6928
rect 19156 6876 19208 6928
rect 36084 6876 36136 6928
rect 40868 6876 40920 6928
rect 14740 6808 14792 6860
rect 14924 6808 14976 6860
rect 34152 6808 34204 6860
rect 5172 6672 5224 6724
rect 12900 6647 12952 6656
rect 12900 6613 12909 6647
rect 12909 6613 12943 6647
rect 12943 6613 12952 6647
rect 12900 6604 12952 6613
rect 14832 6604 14884 6656
rect 23664 6740 23716 6792
rect 25504 6740 25556 6792
rect 37740 6740 37792 6792
rect 40960 6783 41012 6792
rect 40960 6749 40969 6783
rect 40969 6749 41003 6783
rect 41003 6749 41012 6783
rect 40960 6740 41012 6749
rect 43812 6808 43864 6860
rect 45744 6808 45796 6860
rect 22928 6672 22980 6724
rect 25688 6672 25740 6724
rect 43168 6783 43220 6792
rect 43168 6749 43177 6783
rect 43177 6749 43211 6783
rect 43211 6749 43220 6783
rect 43168 6740 43220 6749
rect 43904 6783 43956 6792
rect 43904 6749 43913 6783
rect 43913 6749 43947 6783
rect 43947 6749 43956 6783
rect 43904 6740 43956 6749
rect 43996 6740 44048 6792
rect 22376 6604 22428 6656
rect 22468 6647 22520 6656
rect 22468 6613 22477 6647
rect 22477 6613 22511 6647
rect 22511 6613 22520 6647
rect 22468 6604 22520 6613
rect 23388 6604 23440 6656
rect 42156 6604 42208 6656
rect 43628 6672 43680 6724
rect 42984 6647 43036 6656
rect 42984 6613 42993 6647
rect 42993 6613 43027 6647
rect 43027 6613 43036 6647
rect 42984 6604 43036 6613
rect 43352 6647 43404 6656
rect 43352 6613 43361 6647
rect 43361 6613 43395 6647
rect 43395 6613 43404 6647
rect 43352 6604 43404 6613
rect 44456 6647 44508 6656
rect 44456 6613 44465 6647
rect 44465 6613 44499 6647
rect 44499 6613 44508 6647
rect 44456 6604 44508 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 9680 6400 9732 6452
rect 14924 6400 14976 6452
rect 6920 6332 6972 6384
rect 32496 6400 32548 6452
rect 19156 6332 19208 6384
rect 23940 6332 23992 6384
rect 19616 6264 19668 6316
rect 24032 6264 24084 6316
rect 24676 6264 24728 6316
rect 29184 6264 29236 6316
rect 31760 6264 31812 6316
rect 5448 6196 5500 6248
rect 10600 6128 10652 6180
rect 20628 6196 20680 6248
rect 34520 6196 34572 6248
rect 34980 6239 35032 6248
rect 34980 6205 34989 6239
rect 34989 6205 35023 6239
rect 35023 6205 35032 6239
rect 34980 6196 35032 6205
rect 44088 6443 44140 6452
rect 44088 6409 44097 6443
rect 44097 6409 44131 6443
rect 44131 6409 44140 6443
rect 44088 6400 44140 6409
rect 45376 6400 45428 6452
rect 42800 6332 42852 6384
rect 43996 6332 44048 6384
rect 43536 6307 43588 6316
rect 43536 6273 43545 6307
rect 43545 6273 43579 6307
rect 43579 6273 43588 6307
rect 43536 6264 43588 6273
rect 43628 6264 43680 6316
rect 44272 6307 44324 6316
rect 44272 6273 44281 6307
rect 44281 6273 44315 6307
rect 44315 6273 44324 6307
rect 44272 6264 44324 6273
rect 44364 6196 44416 6248
rect 16672 6103 16724 6112
rect 16672 6069 16681 6103
rect 16681 6069 16715 6103
rect 16715 6069 16724 6103
rect 16672 6060 16724 6069
rect 19064 6060 19116 6112
rect 34428 6128 34480 6180
rect 43904 6128 43956 6180
rect 20444 6103 20496 6112
rect 20444 6069 20453 6103
rect 20453 6069 20487 6103
rect 20487 6069 20496 6103
rect 20444 6060 20496 6069
rect 27252 6103 27304 6112
rect 27252 6069 27261 6103
rect 27261 6069 27295 6103
rect 27295 6069 27304 6103
rect 27252 6060 27304 6069
rect 29920 6060 29972 6112
rect 34244 6060 34296 6112
rect 34520 6060 34572 6112
rect 43720 6103 43772 6112
rect 43720 6069 43729 6103
rect 43729 6069 43763 6103
rect 43763 6069 43772 6103
rect 43720 6060 43772 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 43950 5958 44002 6010
rect 44014 5958 44066 6010
rect 44078 5958 44130 6010
rect 44142 5958 44194 6010
rect 44206 5958 44258 6010
rect 11244 5788 11296 5840
rect 20444 5856 20496 5908
rect 15016 5788 15068 5840
rect 34152 5831 34204 5840
rect 34152 5797 34161 5831
rect 34161 5797 34195 5831
rect 34195 5797 34204 5831
rect 34152 5788 34204 5797
rect 13728 5720 13780 5772
rect 19432 5720 19484 5772
rect 26148 5720 26200 5772
rect 27252 5720 27304 5772
rect 43536 5720 43588 5772
rect 5816 5652 5868 5704
rect 15292 5627 15344 5636
rect 15292 5593 15301 5627
rect 15301 5593 15335 5627
rect 15335 5593 15344 5627
rect 15292 5584 15344 5593
rect 22192 5652 22244 5704
rect 25136 5652 25188 5704
rect 29552 5652 29604 5704
rect 29644 5695 29696 5704
rect 29644 5661 29653 5695
rect 29653 5661 29687 5695
rect 29687 5661 29696 5695
rect 29644 5652 29696 5661
rect 30104 5695 30156 5704
rect 30104 5661 30113 5695
rect 30113 5661 30147 5695
rect 30147 5661 30156 5695
rect 30104 5652 30156 5661
rect 31392 5652 31444 5704
rect 44456 5899 44508 5908
rect 44456 5865 44465 5899
rect 44465 5865 44499 5899
rect 44499 5865 44508 5899
rect 44456 5856 44508 5865
rect 44272 5695 44324 5704
rect 44272 5661 44281 5695
rect 44281 5661 44315 5695
rect 44315 5661 44324 5695
rect 44272 5652 44324 5661
rect 7288 5516 7340 5568
rect 22468 5516 22520 5568
rect 29920 5559 29972 5568
rect 29920 5525 29929 5559
rect 29929 5525 29963 5559
rect 29963 5525 29972 5559
rect 29920 5516 29972 5525
rect 43260 5584 43312 5636
rect 31024 5516 31076 5568
rect 33508 5516 33560 5568
rect 33600 5516 33652 5568
rect 36176 5516 36228 5568
rect 44364 5516 44416 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 9772 5312 9824 5364
rect 19064 5244 19116 5296
rect 31208 5312 31260 5364
rect 33508 5312 33560 5364
rect 20720 5176 20772 5228
rect 24400 5244 24452 5296
rect 26148 5244 26200 5296
rect 31024 5244 31076 5296
rect 31576 5244 31628 5296
rect 24768 5176 24820 5228
rect 30012 5176 30064 5228
rect 44456 5355 44508 5364
rect 44456 5321 44465 5355
rect 44465 5321 44499 5355
rect 44499 5321 44508 5355
rect 44456 5312 44508 5321
rect 23204 5040 23256 5092
rect 6184 4972 6236 5024
rect 22928 4972 22980 5024
rect 31116 5015 31168 5024
rect 31116 4981 31125 5015
rect 31125 4981 31159 5015
rect 31159 4981 31168 5015
rect 31116 4972 31168 4981
rect 31392 5108 31444 5160
rect 33508 5083 33560 5092
rect 33508 5049 33517 5083
rect 33517 5049 33551 5083
rect 33551 5049 33560 5083
rect 33508 5040 33560 5049
rect 44088 5083 44140 5092
rect 44088 5049 44097 5083
rect 44097 5049 44131 5083
rect 44131 5049 44140 5083
rect 44088 5040 44140 5049
rect 41052 4972 41104 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 43950 4870 44002 4922
rect 44014 4870 44066 4922
rect 44078 4870 44130 4922
rect 44142 4870 44194 4922
rect 44206 4870 44258 4922
rect 7656 4768 7708 4820
rect 8392 4768 8444 4820
rect 11428 4768 11480 4820
rect 41144 4811 41196 4820
rect 41144 4777 41153 4811
rect 41153 4777 41187 4811
rect 41187 4777 41196 4811
rect 41144 4768 41196 4777
rect 21456 4700 21508 4752
rect 23388 4700 23440 4752
rect 43628 4700 43680 4752
rect 44456 4743 44508 4752
rect 44456 4709 44465 4743
rect 44465 4709 44499 4743
rect 44499 4709 44508 4743
rect 44456 4700 44508 4709
rect 21824 4632 21876 4684
rect 21916 4632 21968 4684
rect 30656 4564 30708 4616
rect 39672 4564 39724 4616
rect 40776 4607 40828 4616
rect 40776 4573 40785 4607
rect 40785 4573 40819 4607
rect 40819 4573 40828 4607
rect 40776 4564 40828 4573
rect 41052 4564 41104 4616
rect 9496 4496 9548 4548
rect 8300 4428 8352 4480
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19616 4428 19668 4437
rect 19984 4471 20036 4480
rect 19984 4437 19993 4471
rect 19993 4437 20027 4471
rect 20027 4437 20036 4471
rect 19984 4428 20036 4437
rect 42800 4496 42852 4548
rect 44088 4471 44140 4480
rect 44088 4437 44097 4471
rect 44097 4437 44131 4471
rect 44131 4437 44140 4471
rect 44088 4428 44140 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 19984 4224 20036 4276
rect 44364 4224 44416 4276
rect 14280 4156 14332 4208
rect 19616 4156 19668 4208
rect 16304 4088 16356 4140
rect 26884 4088 26936 4140
rect 30380 4088 30432 4140
rect 42616 4088 42668 4140
rect 9864 4020 9916 4072
rect 10324 3952 10376 4004
rect 17684 3952 17736 4004
rect 23388 3952 23440 4004
rect 23664 3995 23716 4004
rect 23664 3961 23673 3995
rect 23673 3961 23707 3995
rect 23707 3961 23716 3995
rect 23664 3952 23716 3961
rect 9404 3884 9456 3936
rect 14188 3884 14240 3936
rect 17500 3884 17552 3936
rect 18788 3884 18840 3936
rect 20444 3884 20496 3936
rect 22192 3927 22244 3936
rect 22192 3893 22201 3927
rect 22201 3893 22235 3927
rect 22235 3893 22244 3927
rect 22192 3884 22244 3893
rect 23296 3927 23348 3936
rect 23296 3893 23305 3927
rect 23305 3893 23339 3927
rect 23339 3893 23348 3927
rect 23296 3884 23348 3893
rect 24216 3927 24268 3936
rect 24216 3893 24225 3927
rect 24225 3893 24259 3927
rect 24259 3893 24268 3927
rect 24216 3884 24268 3893
rect 24584 3927 24636 3936
rect 24584 3893 24593 3927
rect 24593 3893 24627 3927
rect 24627 3893 24636 3927
rect 24584 3884 24636 3893
rect 25596 3927 25648 3936
rect 25596 3893 25605 3927
rect 25605 3893 25639 3927
rect 25639 3893 25648 3927
rect 25596 3884 25648 3893
rect 25872 3884 25924 3936
rect 42800 4020 42852 4072
rect 36544 3952 36596 4004
rect 44088 3995 44140 4004
rect 44088 3961 44097 3995
rect 44097 3961 44131 3995
rect 44131 3961 44140 3995
rect 44088 3952 44140 3961
rect 44456 3995 44508 4004
rect 44456 3961 44465 3995
rect 44465 3961 44499 3995
rect 44499 3961 44508 3995
rect 44456 3952 44508 3961
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 43950 3782 44002 3834
rect 44014 3782 44066 3834
rect 44078 3782 44130 3834
rect 44142 3782 44194 3834
rect 44206 3782 44258 3834
rect 8852 3680 8904 3732
rect 11980 3723 12032 3732
rect 11980 3689 11989 3723
rect 11989 3689 12023 3723
rect 12023 3689 12032 3723
rect 11980 3680 12032 3689
rect 12072 3680 12124 3732
rect 14372 3680 14424 3732
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 20904 3680 20956 3732
rect 27620 3680 27672 3732
rect 9956 3612 10008 3664
rect 38568 3612 38620 3664
rect 44456 3655 44508 3664
rect 44456 3621 44465 3655
rect 44465 3621 44499 3655
rect 44499 3621 44508 3655
rect 44456 3612 44508 3621
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 17500 3476 17552 3528
rect 20996 3544 21048 3596
rect 22652 3544 22704 3596
rect 40684 3544 40736 3596
rect 2136 3340 2188 3392
rect 18604 3408 18656 3460
rect 18696 3408 18748 3460
rect 20812 3476 20864 3528
rect 33784 3476 33836 3528
rect 36544 3476 36596 3528
rect 44364 3476 44416 3528
rect 19432 3340 19484 3392
rect 19524 3383 19576 3392
rect 19524 3349 19533 3383
rect 19533 3349 19567 3383
rect 19567 3349 19576 3383
rect 19524 3340 19576 3349
rect 19800 3340 19852 3392
rect 20260 3340 20312 3392
rect 22652 3340 22704 3392
rect 31576 3408 31628 3460
rect 31760 3408 31812 3460
rect 39948 3408 40000 3460
rect 33784 3340 33836 3392
rect 41696 3340 41748 3392
rect 44088 3383 44140 3392
rect 44088 3349 44097 3383
rect 44097 3349 44131 3383
rect 44131 3349 44140 3383
rect 44088 3340 44140 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 9956 3179 10008 3188
rect 9956 3145 9965 3179
rect 9965 3145 9999 3179
rect 9999 3145 10008 3179
rect 9956 3136 10008 3145
rect 9588 3068 9640 3120
rect 16120 3068 16172 3120
rect 1400 3000 1452 3052
rect 7840 3000 7892 3052
rect 10232 3000 10284 3052
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 14464 3000 14516 3052
rect 20904 3068 20956 3120
rect 16304 3000 16356 3052
rect 17684 3000 17736 3052
rect 16580 2932 16632 2984
rect 19708 3000 19760 3052
rect 21364 3179 21416 3188
rect 21364 3145 21373 3179
rect 21373 3145 21407 3179
rect 21407 3145 21416 3179
rect 21364 3136 21416 3145
rect 23940 3136 23992 3188
rect 25044 3068 25096 3120
rect 23480 3000 23532 3052
rect 24216 3043 24268 3052
rect 24216 3009 24225 3043
rect 24225 3009 24259 3043
rect 24259 3009 24268 3043
rect 24216 3000 24268 3009
rect 25504 3043 25556 3052
rect 25504 3009 25513 3043
rect 25513 3009 25547 3043
rect 25547 3009 25556 3043
rect 25504 3000 25556 3009
rect 32680 3068 32732 3120
rect 29276 3000 29328 3052
rect 36176 3043 36228 3052
rect 36176 3009 36185 3043
rect 36185 3009 36219 3043
rect 36219 3009 36228 3043
rect 36176 3000 36228 3009
rect 36084 2932 36136 2984
rect 37280 3136 37332 3188
rect 38292 3179 38344 3188
rect 38292 3145 38301 3179
rect 38301 3145 38335 3179
rect 38335 3145 38344 3179
rect 38292 3136 38344 3145
rect 42892 3136 42944 3188
rect 40040 3068 40092 3120
rect 37280 3043 37332 3052
rect 37280 3009 37289 3043
rect 37289 3009 37323 3043
rect 37323 3009 37332 3043
rect 37280 3000 37332 3009
rect 37372 3000 37424 3052
rect 40132 3000 40184 3052
rect 44456 3179 44508 3188
rect 44456 3145 44465 3179
rect 44465 3145 44499 3179
rect 44499 3145 44508 3179
rect 44456 3136 44508 3145
rect 43076 2932 43128 2984
rect 35716 2864 35768 2916
rect 38384 2864 38436 2916
rect 44088 2907 44140 2916
rect 44088 2873 44097 2907
rect 44097 2873 44131 2907
rect 44131 2873 44140 2907
rect 44088 2864 44140 2873
rect 15752 2839 15804 2848
rect 15752 2805 15761 2839
rect 15761 2805 15795 2839
rect 15795 2805 15804 2839
rect 15752 2796 15804 2805
rect 16120 2839 16172 2848
rect 16120 2805 16129 2839
rect 16129 2805 16163 2839
rect 16163 2805 16172 2839
rect 16120 2796 16172 2805
rect 17684 2839 17736 2848
rect 17684 2805 17693 2839
rect 17693 2805 17727 2839
rect 17727 2805 17736 2839
rect 17684 2796 17736 2805
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 20260 2796 20312 2848
rect 20536 2796 20588 2848
rect 24860 2796 24912 2848
rect 25688 2839 25740 2848
rect 25688 2805 25697 2839
rect 25697 2805 25731 2839
rect 25731 2805 25740 2839
rect 25688 2796 25740 2805
rect 26700 2839 26752 2848
rect 26700 2805 26709 2839
rect 26709 2805 26743 2839
rect 26743 2805 26752 2839
rect 26700 2796 26752 2805
rect 27712 2839 27764 2848
rect 27712 2805 27721 2839
rect 27721 2805 27755 2839
rect 27755 2805 27764 2839
rect 27712 2796 27764 2805
rect 30288 2796 30340 2848
rect 44824 2796 44876 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 43950 2694 44002 2746
rect 44014 2694 44066 2746
rect 44078 2694 44130 2746
rect 44142 2694 44194 2746
rect 44206 2694 44258 2746
rect 19432 2592 19484 2644
rect 43536 2592 43588 2644
rect 19800 2524 19852 2576
rect 36728 2524 36780 2576
rect 37004 2524 37056 2576
rect 18052 2456 18104 2508
rect 16120 2388 16172 2440
rect 36912 2456 36964 2508
rect 42984 2567 43036 2576
rect 42984 2533 42993 2567
rect 42993 2533 43027 2567
rect 43027 2533 43036 2567
rect 42984 2524 43036 2533
rect 44364 2524 44416 2576
rect 44456 2567 44508 2576
rect 44456 2533 44465 2567
rect 44465 2533 44499 2567
rect 44499 2533 44508 2567
rect 44456 2524 44508 2533
rect 12440 2320 12492 2372
rect 26884 2320 26936 2372
rect 37004 2388 37056 2440
rect 43536 2431 43588 2440
rect 43536 2397 43545 2431
rect 43545 2397 43579 2431
rect 43579 2397 43588 2431
rect 43536 2388 43588 2397
rect 5540 2252 5592 2304
rect 25504 2252 25556 2304
rect 30288 2252 30340 2304
rect 43352 2295 43404 2304
rect 43352 2261 43361 2295
rect 43361 2261 43395 2295
rect 43395 2261 43404 2295
rect 43352 2252 43404 2261
rect 44088 2295 44140 2304
rect 44088 2261 44097 2295
rect 44097 2261 44131 2295
rect 44131 2261 44140 2295
rect 44088 2252 44140 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 31392 212 31444 264
rect 40592 212 40644 264
rect 3884 144 3936 196
rect 6000 144 6052 196
rect 37372 144 37424 196
rect 37280 76 37332 128
rect 1860 8 1912 60
rect 36176 8 36228 60
<< metal2 >>
rect 110 11096 166 11152
rect 478 11096 534 11152
rect 846 11096 902 11152
rect 1214 11096 1270 11152
rect 1582 11096 1638 11152
rect 1950 11096 2006 11152
rect 2318 11096 2374 11152
rect 2686 11096 2742 11152
rect 2884 11110 3004 11138
rect 124 8022 152 11096
rect 112 8016 164 8022
rect 112 7958 164 7964
rect 492 7546 520 11096
rect 860 7750 888 11096
rect 1124 9444 1176 9450
rect 1124 9386 1176 9392
rect 1032 9376 1084 9382
rect 1032 9318 1084 9324
rect 848 7744 900 7750
rect 848 7686 900 7692
rect 480 7540 532 7546
rect 480 7482 532 7488
rect 1044 7177 1072 9318
rect 1136 7721 1164 9386
rect 1228 8090 1256 11096
rect 1596 8634 1624 11096
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1780 8265 1808 8978
rect 1964 8634 1992 11096
rect 2332 8634 2360 11096
rect 2504 8900 2556 8906
rect 2504 8842 2556 8848
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2516 8498 2544 8842
rect 2594 8800 2650 8809
rect 2594 8735 2650 8744
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2608 8401 2636 8735
rect 2700 8634 2728 11096
rect 2884 8634 2912 11110
rect 2976 11098 3004 11110
rect 3054 11098 3110 11152
rect 2976 11096 3110 11098
rect 3422 11096 3478 11152
rect 3790 11096 3846 11152
rect 4158 11096 4214 11152
rect 4526 11096 4582 11152
rect 4894 11096 4950 11152
rect 5262 11096 5318 11152
rect 5630 11096 5686 11152
rect 5998 11096 6054 11152
rect 6366 11096 6422 11152
rect 6734 11096 6790 11152
rect 7102 11096 7158 11152
rect 7470 11096 7526 11152
rect 7838 11096 7894 11152
rect 8206 11096 8262 11152
rect 8574 11096 8630 11152
rect 8942 11096 8998 11152
rect 9310 11096 9366 11152
rect 9678 11096 9734 11152
rect 10046 11096 10102 11152
rect 10414 11096 10470 11152
rect 10782 11096 10838 11152
rect 11150 11096 11206 11152
rect 11518 11096 11574 11152
rect 11886 11096 11942 11152
rect 11978 11112 12034 11121
rect 2976 11070 3096 11096
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3436 8634 3464 11096
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3528 8498 3556 8774
rect 3620 8498 3648 9046
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 2594 8392 2650 8401
rect 2594 8327 2650 8336
rect 1766 8256 1822 8265
rect 1766 8191 1822 8200
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 3804 8090 3832 11096
rect 3974 9072 4030 9081
rect 3974 9007 4030 9016
rect 1216 8084 1268 8090
rect 1216 8026 1268 8032
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 1306 7984 1362 7993
rect 1306 7919 1362 7928
rect 1122 7712 1178 7721
rect 1122 7647 1178 7656
rect 1030 7168 1086 7177
rect 1030 7103 1086 7112
rect 1320 4321 1348 7919
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2332 6934 2360 7822
rect 2424 7002 2452 7822
rect 3988 7818 4016 9007
rect 4172 8634 4200 11096
rect 4344 9240 4396 9246
rect 4344 9182 4396 9188
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4356 8498 4384 9182
rect 4540 8634 4568 11096
rect 4908 8634 4936 11096
rect 5276 8634 5304 11096
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 4172 7342 4200 7822
rect 4724 7585 4752 8434
rect 5092 7993 5120 8434
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5078 7984 5134 7993
rect 5078 7919 5134 7928
rect 4710 7576 4766 7585
rect 4710 7511 4766 7520
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 5184 6730 5212 8366
rect 5262 7848 5318 7857
rect 5262 7783 5264 7792
rect 5316 7783 5318 7792
rect 5264 7754 5316 7760
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 5460 6254 5488 8842
rect 5644 8634 5672 11096
rect 6012 8634 6040 11096
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 5538 6352 5594 6361
rect 5538 6287 5594 6296
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2870 4720 2926 4729
rect 2870 4655 2926 4664
rect 2884 4321 2912 4655
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 1306 4312 1362 4321
rect 1306 4247 1362 4256
rect 2870 4312 2926 4321
rect 3010 4315 3318 4324
rect 2870 4247 2926 4256
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2148 3194 2176 3334
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1412 1193 1440 2994
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 5552 2310 5580 6287
rect 5828 5710 5856 8434
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 6196 5030 6224 8434
rect 6380 8090 6408 11096
rect 6748 8634 6776 11096
rect 7116 8634 7144 11096
rect 7484 8634 7512 11096
rect 7852 8634 7880 11096
rect 8220 8634 8248 11096
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6932 6390 6960 8434
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 7300 5574 7328 8434
rect 7668 7313 7696 8434
rect 7654 7304 7710 7313
rect 7654 7239 7710 7248
rect 7852 6361 7880 8434
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 7838 6352 7894 6361
rect 7838 6287 7894 6296
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 7746 4992 7802 5001
rect 7746 4927 7802 4936
rect 7654 4856 7710 4865
rect 7654 4791 7656 4800
rect 7708 4791 7710 4800
rect 7656 4762 7708 4768
rect 7760 4706 7788 4927
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7930 4720 7986 4729
rect 7760 4678 7930 4706
rect 7930 4655 7986 4664
rect 8312 4486 8340 9046
rect 8588 8294 8616 11096
rect 8956 9466 8984 11096
rect 8864 9438 8984 9466
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8864 8090 8892 9438
rect 9324 8888 9352 11096
rect 9324 8860 9444 8888
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 9416 8616 9444 8860
rect 9692 8650 9720 11096
rect 9864 9308 9916 9314
rect 9864 9250 9916 9256
rect 9324 8588 9444 8616
rect 9508 8622 9720 8650
rect 9324 8294 9352 8588
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8574 7576 8630 7585
rect 8574 7511 8630 7520
rect 8588 7041 8616 7511
rect 8574 7032 8630 7041
rect 8574 6967 8630 6976
rect 8390 4856 8446 4865
rect 8390 4791 8392 4800
rect 8444 4791 8446 4800
rect 8392 4762 8444 4768
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 7470 4176 7526 4185
rect 7470 4111 7526 4120
rect 7484 3505 7512 4111
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 8864 3738 8892 7890
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9416 5545 9444 8434
rect 9508 8294 9536 8622
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9402 5536 9458 5545
rect 9010 5468 9318 5477
rect 9402 5471 9458 5480
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 9508 4554 9536 7822
rect 9600 6984 9628 8502
rect 9876 8498 9904 9250
rect 10060 8514 10088 11096
rect 10324 9240 10376 9246
rect 10324 9182 10376 9188
rect 10138 9072 10194 9081
rect 10138 9007 10194 9016
rect 10232 9036 10284 9042
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9968 8486 10088 8514
rect 9692 7970 9720 8434
rect 9968 8294 9996 8486
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 10152 8090 10180 9007
rect 10232 8978 10284 8984
rect 10244 8362 10272 8978
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 9692 7942 9904 7970
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9600 6956 9720 6984
rect 9586 6896 9642 6905
rect 9586 6831 9642 6840
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 9416 3534 9444 3878
rect 9404 3528 9456 3534
rect 7470 3496 7526 3505
rect 9404 3470 9456 3476
rect 7470 3431 7526 3440
rect 8390 3360 8446 3369
rect 8390 3295 8446 3304
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 1398 1184 1454 1193
rect 1398 1119 1454 1128
rect 3884 196 3936 202
rect 3884 138 3936 144
rect 6000 196 6052 202
rect 6000 138 6052 144
rect 1780 66 1900 82
rect 1780 60 1912 66
rect 1780 56 1860 60
rect 1766 54 1860 56
rect 1766 0 1822 54
rect 3896 56 3924 138
rect 6012 56 6040 138
rect 1860 2 1912 8
rect 3882 0 3938 56
rect 5998 0 6054 56
rect 7852 42 7880 2994
rect 8404 2825 8432 3295
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 9600 3126 9628 6831
rect 9692 6458 9720 6956
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9784 5370 9812 7754
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9876 4078 9904 7942
rect 10138 7304 10194 7313
rect 10138 7239 10194 7248
rect 10152 7041 10180 7239
rect 10138 7032 10194 7041
rect 10138 6967 10194 6976
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 10336 4010 10364 9182
rect 10428 8294 10456 11096
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10520 8498 10548 8910
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10520 8090 10548 8298
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10612 6186 10640 8434
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10704 7546 10732 8366
rect 10796 8294 10824 11096
rect 11058 10704 11114 10713
rect 11058 10639 11114 10648
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10888 8090 10916 8978
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10980 7274 11008 8434
rect 11072 7750 11100 10639
rect 11164 8294 11192 11096
rect 11256 8894 11468 8922
rect 11256 8838 11284 8894
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 11256 5846 11284 8570
rect 11348 8498 11376 8774
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11440 4826 11468 8894
rect 11532 8090 11560 11096
rect 11900 8634 11928 11096
rect 12254 11096 12310 11152
rect 12622 11096 12678 11152
rect 12990 11096 13046 11152
rect 13358 11096 13414 11152
rect 13726 11096 13782 11152
rect 14094 11098 14150 11152
rect 14200 11110 14412 11138
rect 14200 11098 14228 11110
rect 14094 11096 14228 11098
rect 11978 11047 12034 11056
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11992 8022 12020 11047
rect 12268 8634 12296 11096
rect 12530 10976 12586 10985
rect 12530 10911 12586 10920
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 12268 7954 12296 8434
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 7410 11928 7686
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 11992 3738 12020 6938
rect 12084 3738 12112 7414
rect 12452 7410 12480 9114
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12544 6866 12572 10911
rect 12636 8634 12664 11096
rect 13004 8634 13032 11096
rect 13174 10840 13230 10849
rect 13174 10775 13230 10784
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12636 7546 12664 7822
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12912 6662 12940 8298
rect 13188 6866 13216 10775
rect 13372 8634 13400 11096
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13280 7818 13308 8434
rect 13556 7818 13584 8774
rect 13740 8634 13768 11096
rect 14108 11070 14228 11096
rect 13818 10568 13874 10577
rect 13818 10503 13874 10512
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13648 8090 13676 8434
rect 13740 8362 13768 8434
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13740 7177 13768 7346
rect 13726 7168 13782 7177
rect 13726 7103 13782 7112
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 13726 6216 13782 6225
rect 13726 6151 13782 6160
rect 13740 5778 13768 6151
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9968 3194 9996 3606
rect 13832 3534 13860 10503
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14292 7206 14320 8910
rect 14384 8090 14412 11110
rect 14462 11096 14518 11152
rect 14830 11096 14886 11152
rect 15198 11098 15254 11152
rect 15304 11110 15424 11138
rect 15304 11098 15332 11110
rect 15198 11096 15332 11098
rect 14476 8634 14504 11096
rect 14844 8634 14872 11096
rect 15212 11070 15332 11096
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15396 8634 15424 11110
rect 15566 11096 15622 11152
rect 15934 11096 15990 11152
rect 16302 11096 16358 11152
rect 16580 11144 16632 11150
rect 15476 10940 15528 10946
rect 15476 10882 15528 10888
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14646 7984 14702 7993
rect 14646 7919 14702 7928
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14280 7200 14332 7206
rect 14384 7177 14412 7346
rect 14280 7142 14332 7148
rect 14370 7168 14426 7177
rect 13950 7100 14258 7109
rect 14370 7103 14426 7112
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14568 7002 14596 7346
rect 14660 7313 14688 7919
rect 14646 7304 14702 7313
rect 14646 7239 14702 7248
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 14292 4706 14320 6870
rect 14200 4678 14320 4706
rect 14200 3942 14228 4678
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14292 3641 14320 4150
rect 14384 3738 14412 6938
rect 14660 6338 14688 7142
rect 14752 6866 14780 8434
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14844 6662 14872 8434
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15396 7546 15424 8434
rect 15488 7750 15516 10882
rect 15580 8634 15608 11096
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15672 7478 15700 8978
rect 15750 8936 15806 8945
rect 15750 8871 15806 8880
rect 15764 7886 15792 8871
rect 15948 8634 15976 11096
rect 16316 8634 16344 11096
rect 16670 11096 16726 11152
rect 17038 11096 17094 11152
rect 17406 11096 17462 11152
rect 17774 11096 17830 11152
rect 18142 11096 18198 11152
rect 18510 11096 18566 11152
rect 18878 11096 18934 11152
rect 19246 11096 19302 11152
rect 19614 11096 19670 11152
rect 19982 11096 20038 11152
rect 20350 11096 20406 11152
rect 20718 11096 20774 11152
rect 20916 11110 21036 11138
rect 16580 11086 16632 11092
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15856 7546 15884 8434
rect 16224 8090 16252 8434
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 16408 6914 16436 10950
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16500 8090 16528 8434
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16592 7954 16620 11086
rect 16684 8634 16712 11096
rect 16948 9240 17000 9246
rect 16948 9182 17000 9188
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16960 8090 16988 9182
rect 17052 8634 17080 11096
rect 17420 8634 17448 11096
rect 17788 8634 17816 11096
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17420 8090 17448 8434
rect 17788 8090 17816 8434
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16316 6886 16436 6914
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14936 6458 14964 6802
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 14660 6310 15056 6338
rect 15028 5846 15056 6310
rect 15016 5840 15068 5846
rect 15016 5782 15068 5788
rect 15290 5672 15346 5681
rect 15290 5607 15292 5616
rect 15344 5607 15346 5616
rect 15292 5578 15344 5584
rect 14554 5536 14610 5545
rect 14554 5471 14610 5480
rect 14568 5137 14596 5471
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 14554 5128 14610 5137
rect 14554 5063 14610 5072
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 16316 4146 16344 6886
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16684 4729 16712 6054
rect 16776 5001 16804 7890
rect 17880 7546 17908 9046
rect 18064 7886 18092 11018
rect 18156 8634 18184 11096
rect 18524 8634 18552 11096
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18156 8294 18184 8434
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 16762 4992 16818 5001
rect 16762 4927 16818 4936
rect 16670 4720 16726 4729
rect 16670 4655 16726 4664
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14278 3632 14334 3641
rect 14278 3567 14334 3576
rect 17512 3534 17540 3878
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 16120 3120 16172 3126
rect 16172 3068 16344 3074
rect 16120 3062 16344 3068
rect 16132 3058 16344 3062
rect 17696 3058 17724 3946
rect 17972 3738 18000 7278
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 18616 3466 18644 9658
rect 18800 3942 18828 10746
rect 18892 8634 18920 11096
rect 19260 9330 19288 11096
rect 19628 9722 19656 11096
rect 19996 10577 20024 11096
rect 20364 10810 20392 11096
rect 20732 11014 20760 11096
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 19982 10568 20038 10577
rect 19982 10503 20038 10512
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19168 9302 19288 9330
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18892 7342 18920 8434
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 19168 6934 19196 9302
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19260 7970 19288 8366
rect 19260 7954 19380 7970
rect 19260 7948 19392 7954
rect 19260 7942 19340 7948
rect 19340 7890 19392 7896
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19156 6928 19208 6934
rect 19156 6870 19208 6876
rect 19156 6384 19208 6390
rect 19156 6326 19208 6332
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 19076 5302 19104 6054
rect 19064 5296 19116 5302
rect 19168 5273 19196 6326
rect 19444 5778 19472 7686
rect 19628 6322 19656 9046
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20350 8256 20406 8265
rect 19950 8188 20258 8197
rect 20350 8191 20406 8200
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19798 8120 19854 8129
rect 19950 8123 20258 8132
rect 20364 8072 20392 8191
rect 19854 8064 20392 8072
rect 19798 8055 20392 8064
rect 19812 8044 20392 8055
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 19706 6760 19762 6769
rect 19706 6695 19762 6704
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 19064 5238 19116 5244
rect 19154 5264 19210 5273
rect 19154 5199 19210 5208
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19628 4214 19656 4422
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 18696 3460 18748 3466
rect 18696 3402 18748 3408
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 14464 3052 14516 3058
rect 16132 3052 16356 3058
rect 16132 3046 16304 3052
rect 14464 2994 14516 3000
rect 16304 2994 16356 3000
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 8390 2816 8446 2825
rect 7950 2748 8258 2757
rect 8390 2751 8446 2760
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 8036 56 8156 82
rect 10244 56 10272 2994
rect 12360 56 12388 2994
rect 12438 2816 12494 2825
rect 12438 2751 12494 2760
rect 12452 2378 12480 2751
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 14476 56 14504 2994
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 15764 1465 15792 2790
rect 16132 2446 16160 2790
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15750 1456 15806 1465
rect 15750 1391 15806 1400
rect 16592 56 16620 2926
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 17696 2417 17724 2790
rect 18064 2514 18092 2790
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 17682 2408 17738 2417
rect 17682 2343 17738 2352
rect 18708 56 18736 3402
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19444 2650 19472 3334
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19536 1737 19564 3334
rect 19720 3058 19748 6695
rect 20640 6254 20668 8434
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20456 5914 20484 6054
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20534 5264 20590 5273
rect 20534 5199 20590 5208
rect 20720 5228 20772 5234
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19996 4282 20024 4422
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 19800 3392 19852 3398
rect 19800 3334 19852 3340
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19812 2582 19840 3334
rect 20272 2854 20300 3334
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 19800 2576 19852 2582
rect 19800 2518 19852 2524
rect 20456 2009 20484 3878
rect 20548 2854 20576 5199
rect 20720 5170 20772 5176
rect 20732 4185 20760 5170
rect 20718 4176 20774 4185
rect 20916 4162 20944 11110
rect 21008 11098 21036 11110
rect 21086 11098 21142 11152
rect 21008 11096 21142 11098
rect 21454 11096 21510 11152
rect 21822 11096 21878 11152
rect 22190 11096 22246 11152
rect 22558 11096 22614 11152
rect 22926 11096 22982 11152
rect 23294 11096 23350 11152
rect 23662 11096 23718 11152
rect 24030 11096 24086 11152
rect 24398 11096 24454 11152
rect 24766 11096 24822 11152
rect 25134 11096 25190 11152
rect 25502 11096 25558 11152
rect 25870 11096 25926 11152
rect 26238 11096 26294 11152
rect 26606 11098 26662 11152
rect 26712 11110 26924 11138
rect 26712 11098 26740 11110
rect 26606 11096 26740 11098
rect 21008 11070 21128 11096
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21376 9178 21404 10950
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21362 7440 21418 7449
rect 21362 7375 21418 7384
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 20916 4134 21036 4162
rect 20718 4111 20774 4120
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20442 2000 20498 2009
rect 20442 1935 20498 1944
rect 19522 1728 19578 1737
rect 19522 1663 19578 1672
rect 20824 56 20852 3470
rect 20916 3126 20944 3674
rect 21008 3602 21036 4134
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21376 3194 21404 7375
rect 21468 4758 21496 11096
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21560 7041 21588 7686
rect 21546 7032 21602 7041
rect 21546 6967 21602 6976
rect 21456 4752 21508 4758
rect 21456 4694 21508 4700
rect 21836 4690 21864 11096
rect 22008 8016 22060 8022
rect 22008 7958 22060 7964
rect 22020 7818 22048 7958
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21928 4690 21956 7686
rect 22204 5710 22232 11096
rect 22374 9208 22430 9217
rect 22374 9143 22430 9152
rect 22388 6662 22416 9143
rect 22572 9110 22600 11096
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22940 6730 22968 11096
rect 23308 7410 23336 11096
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 23400 6662 23428 8298
rect 23676 6798 23704 11096
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22468 6656 22520 6662
rect 22468 6598 22520 6604
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22480 5574 22508 6598
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 23204 5092 23256 5098
rect 23204 5034 23256 5040
rect 22928 5024 22980 5030
rect 23216 4978 23244 5034
rect 22980 4972 23244 4978
rect 22928 4966 23244 4972
rect 22940 4950 23244 4966
rect 23388 4752 23440 4758
rect 23388 4694 23440 4700
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 23400 4010 23428 4694
rect 23662 4040 23718 4049
rect 23388 4004 23440 4010
rect 23662 3975 23664 3984
rect 23388 3946 23440 3952
rect 23716 3975 23718 3984
rect 23664 3946 23716 3952
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 20904 3120 20956 3126
rect 22204 3097 22232 3878
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 22664 3398 22692 3538
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 23308 3233 23336 3878
rect 23294 3224 23350 3233
rect 23952 3194 23980 6326
rect 24044 6322 24072 11096
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 24412 5302 24440 11096
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24688 5817 24716 6258
rect 24674 5808 24730 5817
rect 24674 5743 24730 5752
rect 24400 5296 24452 5302
rect 24400 5238 24452 5244
rect 24780 5234 24808 11096
rect 25148 5710 25176 11096
rect 25226 8256 25282 8265
rect 25226 8191 25282 8200
rect 25240 8090 25268 8191
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 25516 6798 25544 11096
rect 25780 8560 25832 8566
rect 25780 8502 25832 8508
rect 25792 8022 25820 8502
rect 25596 8016 25648 8022
rect 25594 7984 25596 7993
rect 25780 8016 25832 8022
rect 25648 7984 25650 7993
rect 25780 7958 25832 7964
rect 25884 7954 25912 11096
rect 26252 9466 26280 11096
rect 26620 11070 26740 11096
rect 26252 9438 26372 9466
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25594 7919 25650 7928
rect 25872 7948 25924 7954
rect 25872 7890 25924 7896
rect 26344 7886 26372 9438
rect 26514 9344 26570 9353
rect 26514 9279 26570 9288
rect 26528 7954 26556 9279
rect 26896 8514 26924 11110
rect 26974 11096 27030 11152
rect 27342 11096 27398 11152
rect 27710 11096 27766 11152
rect 28078 11096 28134 11152
rect 28446 11096 28502 11152
rect 28814 11096 28870 11152
rect 29182 11096 29238 11152
rect 29550 11096 29606 11152
rect 29918 11096 29974 11152
rect 30286 11096 30342 11152
rect 30654 11096 30710 11152
rect 31022 11098 31078 11152
rect 31128 11110 31340 11138
rect 31128 11098 31156 11110
rect 31022 11096 31156 11098
rect 26988 9081 27016 11096
rect 27356 10713 27384 11096
rect 27724 10946 27752 11096
rect 27712 10940 27764 10946
rect 27712 10882 27764 10888
rect 27342 10704 27398 10713
rect 27342 10639 27398 10648
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 26974 9072 27030 9081
rect 26974 9007 27030 9016
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 26896 8486 27108 8514
rect 26700 8424 26752 8430
rect 26700 8366 26752 8372
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 26332 7880 26384 7886
rect 26332 7822 26384 7828
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25688 6724 25740 6730
rect 25688 6666 25740 6672
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 24584 3936 24636 3942
rect 25596 3936 25648 3942
rect 24584 3878 24636 3884
rect 25594 3904 25596 3913
rect 25648 3904 25650 3913
rect 24228 3505 24256 3878
rect 24596 3641 24624 3878
rect 25594 3839 25650 3848
rect 24582 3632 24638 3641
rect 24582 3567 24638 3576
rect 24214 3496 24270 3505
rect 24214 3431 24270 3440
rect 24858 3496 24914 3505
rect 24858 3431 24914 3440
rect 23294 3159 23350 3168
rect 23940 3188 23992 3194
rect 23940 3130 23992 3136
rect 20904 3062 20956 3068
rect 22190 3088 22246 3097
rect 22190 3023 22246 3032
rect 23480 3052 23532 3058
rect 23480 2994 23532 3000
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 23492 1442 23520 2994
rect 24228 2961 24256 2994
rect 24214 2952 24270 2961
rect 24214 2887 24270 2896
rect 24872 2854 24900 3431
rect 25044 3120 25096 3126
rect 25044 3062 25096 3068
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 23308 1414 23520 1442
rect 22940 56 23060 82
rect 8036 54 8170 56
rect 8036 42 8064 54
rect 7852 14 8064 42
rect 8114 0 8170 54
rect 10230 0 10286 56
rect 12346 0 12402 56
rect 14462 0 14518 56
rect 16578 0 16634 56
rect 18694 0 18750 56
rect 20810 0 20866 56
rect 22926 54 23060 56
rect 22926 0 22982 54
rect 23032 42 23060 54
rect 23308 42 23336 1414
rect 25056 56 25084 3062
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 25516 2310 25544 2994
rect 25700 2854 25728 6666
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26148 5772 26200 5778
rect 26148 5714 26200 5720
rect 26160 5302 26188 5714
rect 26148 5296 26200 5302
rect 26148 5238 26200 5244
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25872 3936 25924 3942
rect 25872 3878 25924 3884
rect 25884 3097 25912 3878
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25870 3088 25926 3097
rect 25870 3023 25926 3032
rect 26712 2854 26740 8366
rect 26792 8016 26844 8022
rect 26976 8016 27028 8022
rect 26844 7976 26976 8004
rect 26792 7958 26844 7964
rect 26976 7958 27028 7964
rect 27080 7886 27108 8486
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 27068 7880 27120 7886
rect 27068 7822 27120 7828
rect 26896 7546 26924 7822
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27252 6112 27304 6118
rect 27252 6054 27304 6060
rect 27264 5778 27292 6054
rect 27526 5808 27582 5817
rect 27252 5772 27304 5778
rect 27526 5743 27582 5752
rect 27252 5714 27304 5720
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 25688 2848 25740 2854
rect 25688 2790 25740 2796
rect 26700 2848 26752 2854
rect 26700 2790 26752 2796
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26896 2378 26924 4082
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 26884 2372 26936 2378
rect 26884 2314 26936 2320
rect 25504 2304 25556 2310
rect 25504 2246 25556 2252
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27172 56 27292 82
rect 23032 14 23336 42
rect 25042 0 25098 56
rect 27158 54 27292 56
rect 27158 0 27214 54
rect 27264 42 27292 54
rect 27540 42 27568 5743
rect 27632 3738 27660 9114
rect 28092 7886 28120 11096
rect 28460 7886 28488 11096
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 28448 7880 28500 7886
rect 28448 7822 28500 7828
rect 28828 7410 28856 11096
rect 28816 7404 28868 7410
rect 28816 7346 28868 7352
rect 29196 6322 29224 11096
rect 29184 6316 29236 6322
rect 29184 6258 29236 6264
rect 29564 5710 29592 11096
rect 29642 8392 29698 8401
rect 29642 8327 29698 8336
rect 29656 5710 29684 8327
rect 29932 8242 29960 11096
rect 30102 8528 30158 8537
rect 30102 8463 30158 8472
rect 29932 8214 30052 8242
rect 29920 6112 29972 6118
rect 29920 6054 29972 6060
rect 29552 5704 29604 5710
rect 29552 5646 29604 5652
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29932 5574 29960 6054
rect 29920 5568 29972 5574
rect 29920 5510 29972 5516
rect 30024 5234 30052 8214
rect 30116 5710 30144 8463
rect 30300 6882 30328 11096
rect 30300 6854 30420 6882
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 30012 5228 30064 5234
rect 30012 5170 30064 5176
rect 30392 4146 30420 6854
rect 30668 4622 30696 11096
rect 31036 11070 31156 11096
rect 31116 9308 31168 9314
rect 31116 9250 31168 9256
rect 31024 5568 31076 5574
rect 31024 5510 31076 5516
rect 31036 5302 31064 5510
rect 31024 5296 31076 5302
rect 31024 5238 31076 5244
rect 31128 5030 31156 9250
rect 31312 5522 31340 11110
rect 31390 11096 31446 11152
rect 31758 11096 31814 11152
rect 32126 11098 32182 11152
rect 32232 11110 32444 11138
rect 32232 11098 32260 11110
rect 32126 11096 32260 11098
rect 31404 5710 31432 11096
rect 31772 6322 31800 11096
rect 32140 11070 32260 11096
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32416 7410 32444 11110
rect 32494 11096 32550 11152
rect 32862 11096 32918 11152
rect 33230 11098 33286 11152
rect 33336 11110 33548 11138
rect 33336 11098 33364 11110
rect 33230 11096 33364 11098
rect 32404 7404 32456 7410
rect 32404 7346 32456 7352
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 32508 6458 32536 11096
rect 32770 9752 32826 9761
rect 32770 9687 32826 9696
rect 32680 9104 32732 9110
rect 32680 9046 32732 9052
rect 32496 6452 32548 6458
rect 32496 6394 32548 6400
rect 31760 6316 31812 6322
rect 31760 6258 31812 6264
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 31392 5704 31444 5710
rect 31392 5646 31444 5652
rect 31312 5494 31616 5522
rect 31220 5370 31432 5386
rect 31208 5364 31432 5370
rect 31260 5358 31432 5364
rect 31208 5306 31260 5312
rect 31404 5166 31432 5358
rect 31588 5302 31616 5494
rect 31576 5296 31628 5302
rect 31576 5238 31628 5244
rect 31392 5160 31444 5166
rect 31392 5102 31444 5108
rect 31116 5024 31168 5030
rect 31116 4966 31168 4972
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 30656 4616 30708 4622
rect 30656 4558 30708 4564
rect 30380 4140 30432 4146
rect 30380 4082 30432 4088
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 31588 3466 31800 3482
rect 31576 3460 31812 3466
rect 31628 3454 31760 3460
rect 31576 3402 31628 3408
rect 31760 3402 31812 3408
rect 32692 3126 32720 9046
rect 32784 7002 32812 9687
rect 32876 7478 32904 11096
rect 33244 11070 33364 11096
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 33520 7886 33548 11110
rect 33598 11096 33654 11152
rect 33966 11098 34022 11152
rect 33888 11096 34022 11098
rect 34334 11096 34390 11152
rect 34612 11144 34664 11150
rect 33612 7954 33640 11096
rect 33888 11082 34008 11096
rect 33876 11076 34008 11082
rect 33928 11070 34008 11076
rect 33876 11018 33928 11024
rect 34348 9246 34376 11096
rect 34702 11098 34758 11152
rect 34664 11096 34758 11098
rect 35070 11096 35126 11152
rect 35438 11096 35494 11152
rect 35806 11096 35862 11152
rect 36174 11096 36230 11152
rect 36542 11096 36598 11152
rect 36910 11096 36966 11152
rect 37278 11096 37334 11152
rect 37646 11112 37702 11152
rect 34664 11092 34744 11096
rect 34612 11086 34744 11092
rect 34624 11070 34744 11086
rect 34336 9240 34388 9246
rect 34336 9182 34388 9188
rect 35084 8945 35112 11096
rect 35452 9042 35480 11096
rect 35820 9761 35848 11096
rect 35806 9752 35862 9761
rect 35806 9687 35862 9696
rect 36188 9217 36216 11096
rect 36556 10849 36584 11096
rect 36924 10985 36952 11096
rect 37292 11014 37320 11096
rect 38014 11096 38070 11152
rect 38382 11096 38438 11152
rect 38750 11096 38806 11152
rect 39118 11098 39174 11152
rect 39224 11110 39436 11138
rect 39224 11098 39252 11110
rect 39118 11096 39252 11098
rect 37646 11047 37702 11056
rect 37280 11008 37332 11014
rect 36910 10976 36966 10985
rect 37280 10950 37332 10956
rect 36910 10911 36966 10920
rect 36542 10840 36598 10849
rect 36542 10775 36598 10784
rect 38028 10062 38056 11096
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 38016 10056 38068 10062
rect 38016 9998 38068 10004
rect 36174 9208 36230 9217
rect 36174 9143 36230 9152
rect 35440 9036 35492 9042
rect 35440 8978 35492 8984
rect 37200 8974 37228 9998
rect 37188 8968 37240 8974
rect 35070 8936 35126 8945
rect 37188 8910 37240 8916
rect 35070 8871 35126 8880
rect 36452 8900 36504 8906
rect 36452 8842 36504 8848
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 33796 8430 33824 8774
rect 33784 8424 33836 8430
rect 33784 8366 33836 8372
rect 35716 8356 35768 8362
rect 35716 8298 35768 8304
rect 33600 7948 33652 7954
rect 33600 7890 33652 7896
rect 33416 7880 33468 7886
rect 33416 7822 33468 7828
rect 33508 7880 33560 7886
rect 33508 7822 33560 7828
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 32864 7472 32916 7478
rect 32864 7414 32916 7420
rect 32772 6996 32824 7002
rect 32772 6938 32824 6944
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32680 3120 32732 3126
rect 32680 3062 32732 3068
rect 29276 3052 29328 3058
rect 29276 2994 29328 3000
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 27724 2553 27752 2790
rect 27710 2544 27766 2553
rect 27710 2479 27766 2488
rect 29288 56 29316 2994
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 30300 2310 30328 2790
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 33428 1329 33456 7822
rect 34334 7304 34390 7313
rect 34334 7239 34336 7248
rect 34388 7239 34390 7248
rect 34336 7210 34388 7216
rect 34152 6860 34204 6866
rect 34152 6802 34204 6808
rect 34164 5846 34192 6802
rect 34520 6248 34572 6254
rect 34980 6248 35032 6254
rect 34520 6190 34572 6196
rect 34978 6216 34980 6225
rect 35032 6216 35034 6225
rect 34428 6180 34480 6186
rect 34428 6122 34480 6128
rect 34244 6112 34296 6118
rect 34440 6066 34468 6122
rect 34532 6118 34560 6190
rect 34978 6151 35034 6160
rect 34296 6060 34468 6066
rect 34244 6054 34468 6060
rect 34520 6112 34572 6118
rect 34520 6054 34572 6060
rect 34256 6038 34468 6054
rect 34152 5840 34204 5846
rect 34152 5782 34204 5788
rect 33508 5568 33560 5574
rect 33508 5510 33560 5516
rect 33600 5568 33652 5574
rect 33600 5510 33652 5516
rect 33520 5370 33548 5510
rect 33508 5364 33560 5370
rect 33508 5306 33560 5312
rect 33506 5128 33562 5137
rect 33506 5063 33508 5072
rect 33560 5063 33562 5072
rect 33508 5034 33560 5040
rect 33612 2774 33640 5510
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 33796 3398 33824 3470
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 35728 2922 35756 8298
rect 36176 8016 36228 8022
rect 36176 7958 36228 7964
rect 35808 7812 35860 7818
rect 35808 7754 35860 7760
rect 35820 5817 35848 7754
rect 36084 6928 36136 6934
rect 36084 6870 36136 6876
rect 35806 5808 35862 5817
rect 35806 5743 35862 5752
rect 36096 2990 36124 6870
rect 36188 5574 36216 7958
rect 36464 7410 36492 8842
rect 38396 8634 38424 11096
rect 38384 8628 38436 8634
rect 38384 8570 38436 8576
rect 38568 8628 38620 8634
rect 38568 8570 38620 8576
rect 38660 8628 38712 8634
rect 38764 8616 38792 11096
rect 39132 11070 39252 11096
rect 39010 8732 39318 8741
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 39408 8634 39436 11110
rect 39486 11096 39542 11152
rect 39854 11096 39910 11152
rect 40222 11096 40278 11152
rect 40590 11098 40646 11152
rect 40696 11110 40908 11138
rect 40696 11098 40724 11110
rect 40590 11096 40724 11098
rect 39500 8634 39528 11096
rect 39672 9376 39724 9382
rect 39672 9318 39724 9324
rect 39580 9172 39632 9178
rect 39580 9114 39632 9120
rect 39028 8628 39080 8634
rect 38764 8588 39028 8616
rect 38660 8570 38712 8576
rect 39028 8570 39080 8576
rect 39396 8628 39448 8634
rect 39396 8570 39448 8576
rect 39488 8628 39540 8634
rect 39488 8570 39540 8576
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36452 7404 36504 7410
rect 36452 7346 36504 7352
rect 36648 7206 36676 8026
rect 36636 7200 36688 7206
rect 36636 7142 36688 7148
rect 36176 5568 36228 5574
rect 36176 5510 36228 5516
rect 36544 4004 36596 4010
rect 36544 3946 36596 3952
rect 36556 3534 36584 3946
rect 36544 3528 36596 3534
rect 36544 3470 36596 3476
rect 37292 3194 37320 8434
rect 38292 8424 38344 8430
rect 38292 8366 38344 8372
rect 37832 8288 37884 8294
rect 37832 8230 37884 8236
rect 37844 8090 37872 8230
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 37832 8084 37884 8090
rect 37832 8026 37884 8032
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 37740 6792 37792 6798
rect 37740 6734 37792 6740
rect 37280 3188 37332 3194
rect 37280 3130 37332 3136
rect 36176 3052 36228 3058
rect 36176 2994 36228 3000
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 36084 2984 36136 2990
rect 36084 2926 36136 2932
rect 35716 2916 35768 2922
rect 35716 2858 35768 2864
rect 33520 2746 33640 2774
rect 33414 1320 33470 1329
rect 33414 1255 33470 1264
rect 31392 264 31444 270
rect 31392 206 31444 212
rect 31404 56 31432 206
rect 33520 56 33548 2746
rect 35622 1320 35678 1329
rect 35622 1255 35678 1264
rect 35636 56 35664 1255
rect 36188 66 36216 2994
rect 36728 2576 36780 2582
rect 37004 2576 37056 2582
rect 36780 2524 36952 2530
rect 36728 2518 36952 2524
rect 37004 2518 37056 2524
rect 36740 2514 36952 2518
rect 36740 2508 36964 2514
rect 36740 2502 36912 2508
rect 36912 2450 36964 2456
rect 37016 2446 37044 2518
rect 37004 2440 37056 2446
rect 37004 2382 37056 2388
rect 37292 134 37320 2994
rect 37384 202 37412 2994
rect 37372 196 37424 202
rect 37372 138 37424 144
rect 37280 128 37332 134
rect 37280 70 37332 76
rect 36176 60 36228 66
rect 27264 14 27568 42
rect 29274 0 29330 56
rect 31390 0 31446 56
rect 33506 0 33562 56
rect 35622 0 35678 56
rect 37752 56 37780 6734
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 38304 3194 38332 8366
rect 38384 8356 38436 8362
rect 38384 8298 38436 8304
rect 38292 3188 38344 3194
rect 38292 3130 38344 3136
rect 38396 2922 38424 8298
rect 38580 3670 38608 8570
rect 38672 8537 38700 8570
rect 38658 8528 38714 8537
rect 39592 8498 39620 9114
rect 39580 8492 39632 8498
rect 38658 8463 38714 8472
rect 38844 8476 38896 8482
rect 39580 8434 39632 8440
rect 38844 8418 38896 8424
rect 38856 8378 38884 8418
rect 38672 8362 38884 8378
rect 38660 8356 38884 8362
rect 38712 8350 38884 8356
rect 38660 8298 38712 8304
rect 39010 7644 39318 7653
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39010 6556 39318 6565
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 39684 4622 39712 9318
rect 39868 8362 39896 11096
rect 40040 8900 40092 8906
rect 40040 8842 40092 8848
rect 39856 8356 39908 8362
rect 39856 8298 39908 8304
rect 39948 8288 40000 8294
rect 39948 8230 40000 8236
rect 39856 7404 39908 7410
rect 39856 7346 39908 7352
rect 39672 4616 39724 4622
rect 39672 4558 39724 4564
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 38568 3664 38620 3670
rect 38568 3606 38620 3612
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 38384 2916 38436 2922
rect 38384 2858 38436 2864
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 39868 56 39896 7346
rect 39960 3466 39988 8230
rect 40052 8090 40080 8842
rect 40236 8634 40264 11096
rect 40604 11070 40724 11096
rect 40776 8968 40828 8974
rect 40776 8910 40828 8916
rect 40224 8628 40276 8634
rect 40224 8570 40276 8576
rect 40222 8528 40278 8537
rect 40222 8463 40224 8472
rect 40276 8463 40278 8472
rect 40224 8434 40276 8440
rect 40684 8424 40736 8430
rect 40684 8366 40736 8372
rect 40040 8084 40092 8090
rect 40040 8026 40092 8032
rect 40592 7880 40644 7886
rect 40592 7822 40644 7828
rect 40038 3496 40094 3505
rect 39948 3460 40000 3466
rect 40038 3431 40094 3440
rect 39948 3402 40000 3408
rect 40052 3126 40080 3431
rect 40040 3120 40092 3126
rect 40040 3062 40092 3068
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 40144 2961 40172 2994
rect 40130 2952 40186 2961
rect 40130 2887 40186 2896
rect 40604 270 40632 7822
rect 40696 3602 40724 8366
rect 40788 8090 40816 8910
rect 40880 8634 40908 11110
rect 40958 11098 41014 11152
rect 41064 11110 41276 11138
rect 41064 11098 41092 11110
rect 40958 11096 41092 11098
rect 40972 11070 41092 11096
rect 40960 9444 41012 9450
rect 40960 9386 41012 9392
rect 40868 8628 40920 8634
rect 40868 8570 40920 8576
rect 40868 8492 40920 8498
rect 40868 8434 40920 8440
rect 40776 8084 40828 8090
rect 40776 8026 40828 8032
rect 40776 7948 40828 7954
rect 40776 7890 40828 7896
rect 40788 7478 40816 7890
rect 40776 7472 40828 7478
rect 40776 7414 40828 7420
rect 40880 6934 40908 8434
rect 40868 6928 40920 6934
rect 40868 6870 40920 6876
rect 40972 6798 41000 9386
rect 41248 8634 41276 11110
rect 41326 11096 41382 11152
rect 41694 11096 41750 11152
rect 42062 11096 42118 11152
rect 42430 11096 42486 11152
rect 42798 11098 42854 11152
rect 42904 11110 43116 11138
rect 42904 11098 42932 11110
rect 42798 11096 42932 11098
rect 41236 8628 41288 8634
rect 41236 8570 41288 8576
rect 41340 8362 41368 11096
rect 41708 8634 41736 11096
rect 41878 9616 41934 9625
rect 41878 9551 41934 9560
rect 41696 8628 41748 8634
rect 41696 8570 41748 8576
rect 41696 8492 41748 8498
rect 41696 8434 41748 8440
rect 41328 8356 41380 8362
rect 41328 8298 41380 8304
rect 41144 8016 41196 8022
rect 41144 7958 41196 7964
rect 40960 6792 41012 6798
rect 40960 6734 41012 6740
rect 41052 5024 41104 5030
rect 41052 4966 41104 4972
rect 41064 4622 41092 4966
rect 41156 4826 41184 7958
rect 41236 7880 41288 7886
rect 41236 7822 41288 7828
rect 41248 7274 41276 7822
rect 41236 7268 41288 7274
rect 41236 7210 41288 7216
rect 41144 4820 41196 4826
rect 41144 4762 41196 4768
rect 40776 4616 40828 4622
rect 40774 4584 40776 4593
rect 41052 4616 41104 4622
rect 40828 4584 40830 4593
rect 41052 4558 41104 4564
rect 40774 4519 40830 4528
rect 40684 3596 40736 3602
rect 40684 3538 40736 3544
rect 41708 3398 41736 8434
rect 41892 7478 41920 9551
rect 42076 8362 42104 11096
rect 42444 8514 42472 11096
rect 42812 11070 42932 11096
rect 42982 9616 43038 9625
rect 42982 9551 43038 9560
rect 42706 9344 42762 9353
rect 42706 9279 42762 9288
rect 42444 8486 42564 8514
rect 42536 8430 42564 8486
rect 42524 8424 42576 8430
rect 42524 8366 42576 8372
rect 42064 8356 42116 8362
rect 42064 8298 42116 8304
rect 42340 8288 42392 8294
rect 42340 8230 42392 8236
rect 42352 8090 42380 8230
rect 42720 8090 42748 9279
rect 42800 9104 42852 9110
rect 42800 9046 42852 9052
rect 42812 8498 42840 9046
rect 42892 8832 42944 8838
rect 42892 8774 42944 8780
rect 42904 8498 42932 8774
rect 42800 8492 42852 8498
rect 42800 8434 42852 8440
rect 42892 8492 42944 8498
rect 42892 8434 42944 8440
rect 42340 8084 42392 8090
rect 42340 8026 42392 8032
rect 42708 8084 42760 8090
rect 42708 8026 42760 8032
rect 42156 7880 42208 7886
rect 42616 7880 42668 7886
rect 42156 7822 42208 7828
rect 42444 7840 42616 7868
rect 42064 7744 42116 7750
rect 42064 7686 42116 7692
rect 41880 7472 41932 7478
rect 41880 7414 41932 7420
rect 41972 7336 42024 7342
rect 41972 7278 42024 7284
rect 41696 3392 41748 3398
rect 41696 3334 41748 3340
rect 40592 264 40644 270
rect 40592 206 40644 212
rect 41984 56 42012 7278
rect 42076 7206 42104 7686
rect 42064 7200 42116 7206
rect 42064 7142 42116 7148
rect 42168 6662 42196 7822
rect 42444 7410 42472 7840
rect 42616 7822 42668 7828
rect 42996 7546 43024 9551
rect 43088 8616 43116 11110
rect 43166 11098 43222 11152
rect 43272 11110 43484 11138
rect 43272 11098 43300 11110
rect 43166 11096 43300 11098
rect 43180 11070 43300 11096
rect 43350 9072 43406 9081
rect 43350 9007 43406 9016
rect 43260 8628 43312 8634
rect 43088 8588 43260 8616
rect 43260 8570 43312 8576
rect 43260 8492 43312 8498
rect 43260 8434 43312 8440
rect 43272 7970 43300 8434
rect 43088 7942 43300 7970
rect 42616 7540 42668 7546
rect 42984 7540 43036 7546
rect 42668 7500 42840 7528
rect 42616 7482 42668 7488
rect 42812 7410 42840 7500
rect 42984 7482 43036 7488
rect 42432 7404 42484 7410
rect 42432 7346 42484 7352
rect 42800 7404 42852 7410
rect 42800 7346 42852 7352
rect 42616 7268 42668 7274
rect 42800 7268 42852 7274
rect 42668 7228 42800 7256
rect 42616 7210 42668 7216
rect 42800 7210 42852 7216
rect 42156 6656 42208 6662
rect 42156 6598 42208 6604
rect 42984 6656 43036 6662
rect 42984 6598 43036 6604
rect 42800 6384 42852 6390
rect 42996 6361 43024 6598
rect 42800 6326 42852 6332
rect 42982 6352 43038 6361
rect 42812 4554 42840 6326
rect 42982 6287 43038 6296
rect 42800 4548 42852 4554
rect 42800 4490 42852 4496
rect 42616 4140 42668 4146
rect 42616 4082 42668 4088
rect 42628 3097 42656 4082
rect 42800 4072 42852 4078
rect 42800 4014 42852 4020
rect 42890 4040 42946 4049
rect 42812 3641 42840 4014
rect 42890 3975 42946 3984
rect 42798 3632 42854 3641
rect 42798 3567 42854 3576
rect 42904 3194 42932 3975
rect 42892 3188 42944 3194
rect 42892 3130 42944 3136
rect 42614 3088 42670 3097
rect 42614 3023 42670 3032
rect 43088 2990 43116 7942
rect 43166 7848 43222 7857
rect 43166 7783 43222 7792
rect 43180 7410 43208 7783
rect 43364 7546 43392 9007
rect 43456 8362 43484 11110
rect 43534 11096 43590 11152
rect 43732 11110 43852 11138
rect 43548 9602 43576 11096
rect 43548 9574 43668 9602
rect 43536 8900 43588 8906
rect 43536 8842 43588 8848
rect 43548 8498 43576 8842
rect 43640 8566 43668 9574
rect 43628 8560 43680 8566
rect 43628 8502 43680 8508
rect 43536 8492 43588 8498
rect 43536 8434 43588 8440
rect 43626 8392 43682 8401
rect 43444 8356 43496 8362
rect 43626 8327 43682 8336
rect 43444 8298 43496 8304
rect 43536 8084 43588 8090
rect 43536 8026 43588 8032
rect 43548 7993 43576 8026
rect 43534 7984 43590 7993
rect 43444 7948 43496 7954
rect 43534 7919 43590 7928
rect 43444 7890 43496 7896
rect 43352 7540 43404 7546
rect 43352 7482 43404 7488
rect 43168 7404 43220 7410
rect 43168 7346 43220 7352
rect 43260 7404 43312 7410
rect 43260 7346 43312 7352
rect 43168 6792 43220 6798
rect 43168 6734 43220 6740
rect 43180 5273 43208 6734
rect 43272 5642 43300 7346
rect 43456 7002 43484 7890
rect 43444 6996 43496 7002
rect 43444 6938 43496 6944
rect 43640 6730 43668 8327
rect 43732 8090 43760 11110
rect 43824 11098 43852 11110
rect 43902 11098 43958 11152
rect 43824 11096 43958 11098
rect 44270 11096 44326 11152
rect 44638 11096 44694 11152
rect 45006 11096 45062 11152
rect 45374 11096 45430 11152
rect 45742 11096 45798 11152
rect 43824 11070 43944 11096
rect 43996 8968 44048 8974
rect 43996 8910 44048 8916
rect 43810 8528 43866 8537
rect 44008 8498 44036 8910
rect 43810 8463 43866 8472
rect 43996 8492 44048 8498
rect 43720 8084 43772 8090
rect 43720 8026 43772 8032
rect 43824 7546 43852 8463
rect 43996 8434 44048 8440
rect 44284 8242 44312 11096
rect 44652 8294 44680 11096
rect 44640 8288 44692 8294
rect 44454 8256 44510 8265
rect 44284 8214 44404 8242
rect 43950 8188 44258 8197
rect 43950 8186 43956 8188
rect 44012 8186 44036 8188
rect 44092 8186 44116 8188
rect 44172 8186 44196 8188
rect 44252 8186 44258 8188
rect 44012 8134 44014 8186
rect 44194 8134 44196 8186
rect 43950 8132 43956 8134
rect 44012 8132 44036 8134
rect 44092 8132 44116 8134
rect 44172 8132 44196 8134
rect 44252 8132 44258 8134
rect 43950 8123 44258 8132
rect 44376 7546 44404 8214
rect 44640 8230 44692 8236
rect 44454 8191 44510 8200
rect 44468 7954 44496 8191
rect 44456 7948 44508 7954
rect 44456 7890 44508 7896
rect 44824 7812 44876 7818
rect 44824 7754 44876 7760
rect 44836 7721 44864 7754
rect 44822 7712 44878 7721
rect 44822 7647 44878 7656
rect 43812 7540 43864 7546
rect 43812 7482 43864 7488
rect 44364 7540 44416 7546
rect 44364 7482 44416 7488
rect 44456 7540 44508 7546
rect 44456 7482 44508 7488
rect 44468 7449 44496 7482
rect 44454 7440 44510 7449
rect 44364 7404 44416 7410
rect 44454 7375 44510 7384
rect 44364 7346 44416 7352
rect 43812 7336 43864 7342
rect 43812 7278 43864 7284
rect 43824 7002 43852 7278
rect 43950 7100 44258 7109
rect 43950 7098 43956 7100
rect 44012 7098 44036 7100
rect 44092 7098 44116 7100
rect 44172 7098 44196 7100
rect 44252 7098 44258 7100
rect 44012 7046 44014 7098
rect 44194 7046 44196 7098
rect 43950 7044 43956 7046
rect 44012 7044 44036 7046
rect 44092 7044 44116 7046
rect 44172 7044 44196 7046
rect 44252 7044 44258 7046
rect 43950 7035 44258 7044
rect 43812 6996 43864 7002
rect 43812 6938 43864 6944
rect 44272 6996 44324 7002
rect 44272 6938 44324 6944
rect 44086 6896 44142 6905
rect 43812 6860 43864 6866
rect 44086 6831 44142 6840
rect 43812 6802 43864 6808
rect 43628 6724 43680 6730
rect 43628 6666 43680 6672
rect 43352 6656 43404 6662
rect 43350 6624 43352 6633
rect 43404 6624 43406 6633
rect 43350 6559 43406 6568
rect 43536 6316 43588 6322
rect 43536 6258 43588 6264
rect 43628 6316 43680 6322
rect 43628 6258 43680 6264
rect 43548 5778 43576 6258
rect 43536 5772 43588 5778
rect 43536 5714 43588 5720
rect 43260 5636 43312 5642
rect 43260 5578 43312 5584
rect 43166 5264 43222 5273
rect 43166 5199 43222 5208
rect 43640 4758 43668 6258
rect 43720 6112 43772 6118
rect 43720 6054 43772 6060
rect 43732 5817 43760 6054
rect 43718 5808 43774 5817
rect 43718 5743 43774 5752
rect 43628 4752 43680 4758
rect 43628 4694 43680 4700
rect 43076 2984 43128 2990
rect 43076 2926 43128 2932
rect 43536 2644 43588 2650
rect 43536 2586 43588 2592
rect 42984 2576 43036 2582
rect 42984 2518 43036 2524
rect 42996 1737 43024 2518
rect 43548 2446 43576 2586
rect 43536 2440 43588 2446
rect 43536 2382 43588 2388
rect 43352 2304 43404 2310
rect 43352 2246 43404 2252
rect 42982 1728 43038 1737
rect 42982 1663 43038 1672
rect 43364 1465 43392 2246
rect 43350 1456 43406 1465
rect 43350 1391 43406 1400
rect 36176 2 36228 8
rect 37738 0 37794 56
rect 39854 0 39910 56
rect 41970 0 42026 56
rect 43824 42 43852 6802
rect 43904 6792 43956 6798
rect 43904 6734 43956 6740
rect 43996 6792 44048 6798
rect 43996 6734 44048 6740
rect 43916 6186 43944 6734
rect 44008 6390 44036 6734
rect 44100 6458 44128 6831
rect 44088 6452 44140 6458
rect 44088 6394 44140 6400
rect 43996 6384 44048 6390
rect 43996 6326 44048 6332
rect 44284 6322 44312 6938
rect 44272 6316 44324 6322
rect 44272 6258 44324 6264
rect 44376 6254 44404 7346
rect 45020 7206 45048 11096
rect 45008 7200 45060 7206
rect 44454 7168 44510 7177
rect 45008 7142 45060 7148
rect 44454 7103 44510 7112
rect 44468 6662 44496 7103
rect 44456 6656 44508 6662
rect 44456 6598 44508 6604
rect 45388 6458 45416 11096
rect 45756 6866 45784 11096
rect 45744 6860 45796 6866
rect 45744 6802 45796 6808
rect 45376 6452 45428 6458
rect 45376 6394 45428 6400
rect 44364 6248 44416 6254
rect 44364 6190 44416 6196
rect 43904 6180 43956 6186
rect 43904 6122 43956 6128
rect 44454 6080 44510 6089
rect 43950 6012 44258 6021
rect 44454 6015 44510 6024
rect 43950 6010 43956 6012
rect 44012 6010 44036 6012
rect 44092 6010 44116 6012
rect 44172 6010 44196 6012
rect 44252 6010 44258 6012
rect 44012 5958 44014 6010
rect 44194 5958 44196 6010
rect 43950 5956 43956 5958
rect 44012 5956 44036 5958
rect 44092 5956 44116 5958
rect 44172 5956 44196 5958
rect 44252 5956 44258 5958
rect 43950 5947 44258 5956
rect 44468 5914 44496 6015
rect 44456 5908 44508 5914
rect 44456 5850 44508 5856
rect 44272 5704 44324 5710
rect 44270 5672 44272 5681
rect 44324 5672 44326 5681
rect 44270 5607 44326 5616
rect 44364 5568 44416 5574
rect 44362 5536 44364 5545
rect 44416 5536 44418 5545
rect 44362 5471 44418 5480
rect 44456 5364 44508 5370
rect 44456 5306 44508 5312
rect 44468 5273 44496 5306
rect 44454 5264 44510 5273
rect 44454 5199 44510 5208
rect 44086 5128 44142 5137
rect 44086 5063 44088 5072
rect 44140 5063 44142 5072
rect 44088 5034 44140 5040
rect 43950 4924 44258 4933
rect 43950 4922 43956 4924
rect 44012 4922 44036 4924
rect 44092 4922 44116 4924
rect 44172 4922 44196 4924
rect 44252 4922 44258 4924
rect 44012 4870 44014 4922
rect 44194 4870 44196 4922
rect 43950 4868 43956 4870
rect 44012 4868 44036 4870
rect 44092 4868 44116 4870
rect 44172 4868 44196 4870
rect 44252 4868 44258 4870
rect 43950 4859 44258 4868
rect 44456 4752 44508 4758
rect 44454 4720 44456 4729
rect 44508 4720 44510 4729
rect 44454 4655 44510 4664
rect 44088 4480 44140 4486
rect 44086 4448 44088 4457
rect 44140 4448 44142 4457
rect 44086 4383 44142 4392
rect 44364 4276 44416 4282
rect 44364 4218 44416 4224
rect 44086 4040 44142 4049
rect 44086 3975 44088 3984
rect 44140 3975 44142 3984
rect 44088 3946 44140 3952
rect 43950 3836 44258 3845
rect 43950 3834 43956 3836
rect 44012 3834 44036 3836
rect 44092 3834 44116 3836
rect 44172 3834 44196 3836
rect 44252 3834 44258 3836
rect 44012 3782 44014 3834
rect 44194 3782 44196 3834
rect 43950 3780 43956 3782
rect 44012 3780 44036 3782
rect 44092 3780 44116 3782
rect 44172 3780 44196 3782
rect 44252 3780 44258 3782
rect 43950 3771 44258 3780
rect 44376 3534 44404 4218
rect 44454 4176 44510 4185
rect 44454 4111 44510 4120
rect 44468 4010 44496 4111
rect 44456 4004 44508 4010
rect 44456 3946 44508 3952
rect 44456 3664 44508 3670
rect 44454 3632 44456 3641
rect 44508 3632 44510 3641
rect 44454 3567 44510 3576
rect 44364 3528 44416 3534
rect 44364 3470 44416 3476
rect 44088 3392 44140 3398
rect 44086 3360 44088 3369
rect 44140 3360 44142 3369
rect 44086 3295 44142 3304
rect 44456 3188 44508 3194
rect 44456 3130 44508 3136
rect 44468 3097 44496 3130
rect 44454 3088 44510 3097
rect 44454 3023 44510 3032
rect 44086 2952 44142 2961
rect 44086 2887 44088 2896
rect 44140 2887 44142 2896
rect 44088 2858 44140 2864
rect 44824 2848 44876 2854
rect 44824 2790 44876 2796
rect 43950 2748 44258 2757
rect 43950 2746 43956 2748
rect 44012 2746 44036 2748
rect 44092 2746 44116 2748
rect 44172 2746 44196 2748
rect 44252 2746 44258 2748
rect 44012 2694 44014 2746
rect 44194 2694 44196 2746
rect 43950 2692 43956 2694
rect 44012 2692 44036 2694
rect 44092 2692 44116 2694
rect 44172 2692 44196 2694
rect 44252 2692 44258 2694
rect 43950 2683 44258 2692
rect 44364 2576 44416 2582
rect 44456 2576 44508 2582
rect 44364 2518 44416 2524
rect 44454 2544 44456 2553
rect 44508 2544 44510 2553
rect 44088 2304 44140 2310
rect 44086 2272 44088 2281
rect 44140 2272 44142 2281
rect 44086 2207 44142 2216
rect 44376 1193 44404 2518
rect 44454 2479 44510 2488
rect 44836 2009 44864 2790
rect 44822 2000 44878 2009
rect 44822 1935 44878 1944
rect 44362 1184 44418 1193
rect 44362 1119 44418 1128
rect 44008 56 44128 82
rect 44008 54 44142 56
rect 44008 42 44036 54
rect 43824 14 44036 42
rect 44086 0 44142 54
<< via2 >>
rect 2594 8744 2650 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 2594 8336 2650 8392
rect 1766 8200 1822 8256
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 3974 9016 4030 9072
rect 1306 7928 1362 7984
rect 1122 7656 1178 7712
rect 1030 7112 1086 7168
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 5078 7928 5134 7984
rect 4710 7520 4766 7576
rect 5262 7812 5318 7848
rect 5262 7792 5264 7812
rect 5264 7792 5316 7812
rect 5316 7792 5318 7812
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 5538 6296 5594 6352
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2870 4664 2926 4720
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 1306 4256 1362 4312
rect 2870 4256 2926 4312
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 7654 7248 7710 7304
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 7838 6296 7894 6352
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 7746 4936 7802 4992
rect 7654 4820 7710 4856
rect 7654 4800 7656 4820
rect 7656 4800 7708 4820
rect 7708 4800 7710 4820
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7930 4664 7986 4720
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 8574 7520 8630 7576
rect 8574 6976 8630 7032
rect 8390 4820 8446 4856
rect 8390 4800 8392 4820
rect 8392 4800 8444 4820
rect 8444 4800 8446 4820
rect 7470 4120 7526 4176
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9402 5480 9458 5536
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 10138 9016 10194 9072
rect 9586 6840 9642 6896
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 7470 3440 7526 3496
rect 8390 3304 8446 3360
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 1398 1128 1454 1184
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 10138 7248 10194 7304
rect 10138 6976 10194 7032
rect 11058 10648 11114 10704
rect 11978 11056 12034 11112
rect 12530 10920 12586 10976
rect 13174 10784 13230 10840
rect 13818 10512 13874 10568
rect 13726 7112 13782 7168
rect 13726 6160 13782 6216
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 14646 7928 14702 7984
rect 14370 7112 14426 7168
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 14646 7248 14702 7304
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15750 8880 15806 8936
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 15290 5636 15346 5672
rect 15290 5616 15292 5636
rect 15292 5616 15344 5636
rect 15344 5616 15346 5636
rect 14554 5480 14610 5536
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 14554 5072 14610 5128
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 16762 4936 16818 4992
rect 16670 4664 16726 4720
rect 14278 3576 14334 3632
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 19982 10512 20038 10568
rect 20350 8200 20406 8256
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19798 8064 19854 8120
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19706 6704 19762 6760
rect 19154 5208 19210 5264
rect 8390 2760 8446 2816
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 12438 2760 12494 2816
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 15750 1400 15806 1456
rect 17682 2352 17738 2408
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 20534 5208 20590 5264
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 20718 4120 20774 4176
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21362 7384 21418 7440
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 20442 1944 20498 2000
rect 19522 1672 19578 1728
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21546 6976 21602 7032
rect 22374 9152 22430 9208
rect 23662 4004 23718 4040
rect 23662 3984 23664 4004
rect 23664 3984 23716 4004
rect 23716 3984 23718 4004
rect 23294 3168 23350 3224
rect 24674 5752 24730 5808
rect 25226 8200 25282 8256
rect 25594 7964 25596 7984
rect 25596 7964 25648 7984
rect 25648 7964 25650 7984
rect 25594 7928 25650 7964
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 26514 9288 26570 9344
rect 27342 10648 27398 10704
rect 26974 9016 27030 9072
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25594 3884 25596 3904
rect 25596 3884 25648 3904
rect 25648 3884 25650 3904
rect 25594 3848 25650 3884
rect 24582 3576 24638 3632
rect 24214 3440 24270 3496
rect 24858 3440 24914 3496
rect 22190 3032 22246 3088
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 24214 2896 24270 2952
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25870 3032 25926 3088
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27526 5752 27582 5808
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 29642 8336 29698 8392
rect 30102 8472 30158 8528
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 32770 9696 32826 9752
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 35806 9696 35862 9752
rect 37646 11056 37702 11112
rect 36910 10920 36966 10976
rect 36542 10784 36598 10840
rect 36174 9152 36230 9208
rect 35070 8880 35126 8936
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 27710 2488 27766 2544
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 34334 7268 34390 7304
rect 34334 7248 34336 7268
rect 34336 7248 34388 7268
rect 34388 7248 34390 7268
rect 34978 6196 34980 6216
rect 34980 6196 35032 6216
rect 35032 6196 35034 6216
rect 34978 6160 35034 6196
rect 33506 5092 33562 5128
rect 33506 5072 33508 5092
rect 33508 5072 33560 5092
rect 33560 5072 33562 5092
rect 35806 5752 35862 5808
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 33414 1264 33470 1320
rect 35622 1264 35678 1320
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 38658 8472 38714 8528
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 40222 8492 40278 8528
rect 40222 8472 40224 8492
rect 40224 8472 40276 8492
rect 40276 8472 40278 8492
rect 40038 3440 40094 3496
rect 40130 2896 40186 2952
rect 41878 9560 41934 9616
rect 40774 4564 40776 4584
rect 40776 4564 40828 4584
rect 40828 4564 40830 4584
rect 40774 4528 40830 4564
rect 42982 9560 43038 9616
rect 42706 9288 42762 9344
rect 43350 9016 43406 9072
rect 42982 6296 43038 6352
rect 42890 3984 42946 4040
rect 42798 3576 42854 3632
rect 42614 3032 42670 3088
rect 43166 7792 43222 7848
rect 43626 8336 43682 8392
rect 43534 7928 43590 7984
rect 43810 8472 43866 8528
rect 43956 8186 44012 8188
rect 44036 8186 44092 8188
rect 44116 8186 44172 8188
rect 44196 8186 44252 8188
rect 43956 8134 44002 8186
rect 44002 8134 44012 8186
rect 44036 8134 44066 8186
rect 44066 8134 44078 8186
rect 44078 8134 44092 8186
rect 44116 8134 44130 8186
rect 44130 8134 44142 8186
rect 44142 8134 44172 8186
rect 44196 8134 44206 8186
rect 44206 8134 44252 8186
rect 43956 8132 44012 8134
rect 44036 8132 44092 8134
rect 44116 8132 44172 8134
rect 44196 8132 44252 8134
rect 44454 8200 44510 8256
rect 44822 7656 44878 7712
rect 44454 7384 44510 7440
rect 43956 7098 44012 7100
rect 44036 7098 44092 7100
rect 44116 7098 44172 7100
rect 44196 7098 44252 7100
rect 43956 7046 44002 7098
rect 44002 7046 44012 7098
rect 44036 7046 44066 7098
rect 44066 7046 44078 7098
rect 44078 7046 44092 7098
rect 44116 7046 44130 7098
rect 44130 7046 44142 7098
rect 44142 7046 44172 7098
rect 44196 7046 44206 7098
rect 44206 7046 44252 7098
rect 43956 7044 44012 7046
rect 44036 7044 44092 7046
rect 44116 7044 44172 7046
rect 44196 7044 44252 7046
rect 44086 6840 44142 6896
rect 43350 6604 43352 6624
rect 43352 6604 43404 6624
rect 43404 6604 43406 6624
rect 43350 6568 43406 6604
rect 43166 5208 43222 5264
rect 43718 5752 43774 5808
rect 42982 1672 43038 1728
rect 43350 1400 43406 1456
rect 44454 7112 44510 7168
rect 44454 6024 44510 6080
rect 43956 6010 44012 6012
rect 44036 6010 44092 6012
rect 44116 6010 44172 6012
rect 44196 6010 44252 6012
rect 43956 5958 44002 6010
rect 44002 5958 44012 6010
rect 44036 5958 44066 6010
rect 44066 5958 44078 6010
rect 44078 5958 44092 6010
rect 44116 5958 44130 6010
rect 44130 5958 44142 6010
rect 44142 5958 44172 6010
rect 44196 5958 44206 6010
rect 44206 5958 44252 6010
rect 43956 5956 44012 5958
rect 44036 5956 44092 5958
rect 44116 5956 44172 5958
rect 44196 5956 44252 5958
rect 44270 5652 44272 5672
rect 44272 5652 44324 5672
rect 44324 5652 44326 5672
rect 44270 5616 44326 5652
rect 44362 5516 44364 5536
rect 44364 5516 44416 5536
rect 44416 5516 44418 5536
rect 44362 5480 44418 5516
rect 44454 5208 44510 5264
rect 44086 5092 44142 5128
rect 44086 5072 44088 5092
rect 44088 5072 44140 5092
rect 44140 5072 44142 5092
rect 43956 4922 44012 4924
rect 44036 4922 44092 4924
rect 44116 4922 44172 4924
rect 44196 4922 44252 4924
rect 43956 4870 44002 4922
rect 44002 4870 44012 4922
rect 44036 4870 44066 4922
rect 44066 4870 44078 4922
rect 44078 4870 44092 4922
rect 44116 4870 44130 4922
rect 44130 4870 44142 4922
rect 44142 4870 44172 4922
rect 44196 4870 44206 4922
rect 44206 4870 44252 4922
rect 43956 4868 44012 4870
rect 44036 4868 44092 4870
rect 44116 4868 44172 4870
rect 44196 4868 44252 4870
rect 44454 4700 44456 4720
rect 44456 4700 44508 4720
rect 44508 4700 44510 4720
rect 44454 4664 44510 4700
rect 44086 4428 44088 4448
rect 44088 4428 44140 4448
rect 44140 4428 44142 4448
rect 44086 4392 44142 4428
rect 44086 4004 44142 4040
rect 44086 3984 44088 4004
rect 44088 3984 44140 4004
rect 44140 3984 44142 4004
rect 43956 3834 44012 3836
rect 44036 3834 44092 3836
rect 44116 3834 44172 3836
rect 44196 3834 44252 3836
rect 43956 3782 44002 3834
rect 44002 3782 44012 3834
rect 44036 3782 44066 3834
rect 44066 3782 44078 3834
rect 44078 3782 44092 3834
rect 44116 3782 44130 3834
rect 44130 3782 44142 3834
rect 44142 3782 44172 3834
rect 44196 3782 44206 3834
rect 44206 3782 44252 3834
rect 43956 3780 44012 3782
rect 44036 3780 44092 3782
rect 44116 3780 44172 3782
rect 44196 3780 44252 3782
rect 44454 4120 44510 4176
rect 44454 3612 44456 3632
rect 44456 3612 44508 3632
rect 44508 3612 44510 3632
rect 44454 3576 44510 3612
rect 44086 3340 44088 3360
rect 44088 3340 44140 3360
rect 44140 3340 44142 3360
rect 44086 3304 44142 3340
rect 44454 3032 44510 3088
rect 44086 2916 44142 2952
rect 44086 2896 44088 2916
rect 44088 2896 44140 2916
rect 44140 2896 44142 2916
rect 43956 2746 44012 2748
rect 44036 2746 44092 2748
rect 44116 2746 44172 2748
rect 44196 2746 44252 2748
rect 43956 2694 44002 2746
rect 44002 2694 44012 2746
rect 44036 2694 44066 2746
rect 44066 2694 44078 2746
rect 44078 2694 44092 2746
rect 44116 2694 44130 2746
rect 44130 2694 44142 2746
rect 44142 2694 44172 2746
rect 44196 2694 44206 2746
rect 44206 2694 44252 2746
rect 43956 2692 44012 2694
rect 44036 2692 44092 2694
rect 44116 2692 44172 2694
rect 44196 2692 44252 2694
rect 44454 2524 44456 2544
rect 44456 2524 44508 2544
rect 44508 2524 44510 2544
rect 44086 2252 44088 2272
rect 44088 2252 44140 2272
rect 44140 2252 44142 2272
rect 44086 2216 44142 2252
rect 44454 2488 44510 2524
rect 44822 1944 44878 2000
rect 44362 1128 44418 1184
<< metal3 >>
rect 11973 11114 12039 11117
rect 37641 11114 37707 11117
rect 11973 11112 37707 11114
rect 11973 11056 11978 11112
rect 12034 11056 37646 11112
rect 37702 11056 37707 11112
rect 11973 11054 37707 11056
rect 11973 11051 12039 11054
rect 37641 11051 37707 11054
rect 12525 10978 12591 10981
rect 36905 10978 36971 10981
rect 12525 10976 36971 10978
rect 12525 10920 12530 10976
rect 12586 10920 36910 10976
rect 36966 10920 36971 10976
rect 12525 10918 36971 10920
rect 12525 10915 12591 10918
rect 36905 10915 36971 10918
rect 13169 10842 13235 10845
rect 36537 10842 36603 10845
rect 13169 10840 36603 10842
rect 13169 10784 13174 10840
rect 13230 10784 36542 10840
rect 36598 10784 36603 10840
rect 13169 10782 36603 10784
rect 13169 10779 13235 10782
rect 36537 10779 36603 10782
rect 11053 10706 11119 10709
rect 27337 10706 27403 10709
rect 11053 10704 27403 10706
rect 11053 10648 11058 10704
rect 11114 10648 27342 10704
rect 27398 10648 27403 10704
rect 11053 10646 27403 10648
rect 11053 10643 11119 10646
rect 27337 10643 27403 10646
rect 13813 10570 13879 10573
rect 19977 10570 20043 10573
rect 13813 10568 20043 10570
rect 13813 10512 13818 10568
rect 13874 10512 19982 10568
rect 20038 10512 20043 10568
rect 13813 10510 20043 10512
rect 13813 10507 13879 10510
rect 19977 10507 20043 10510
rect 32765 9754 32831 9757
rect 35801 9754 35867 9757
rect 32765 9752 35867 9754
rect 32765 9696 32770 9752
rect 32826 9696 35806 9752
rect 35862 9696 35867 9752
rect 32765 9694 35867 9696
rect 32765 9691 32831 9694
rect 35801 9691 35867 9694
rect 0 9618 120 9648
rect 41873 9618 41939 9621
rect 0 9616 41939 9618
rect 0 9560 41878 9616
rect 41934 9560 41939 9616
rect 0 9558 41939 9560
rect 0 9528 120 9558
rect 41873 9555 41939 9558
rect 42977 9618 43043 9621
rect 45880 9618 46000 9648
rect 42977 9616 46000 9618
rect 42977 9560 42982 9616
rect 43038 9560 46000 9616
rect 42977 9558 46000 9560
rect 42977 9555 43043 9558
rect 45880 9528 46000 9558
rect 0 9346 120 9376
rect 26509 9346 26575 9349
rect 0 9344 26575 9346
rect 0 9288 26514 9344
rect 26570 9288 26575 9344
rect 0 9286 26575 9288
rect 0 9256 120 9286
rect 26509 9283 26575 9286
rect 42701 9346 42767 9349
rect 45880 9346 46000 9376
rect 42701 9344 46000 9346
rect 42701 9288 42706 9344
rect 42762 9288 46000 9344
rect 42701 9286 46000 9288
rect 42701 9283 42767 9286
rect 45880 9256 46000 9286
rect 22369 9210 22435 9213
rect 36169 9210 36235 9213
rect 22369 9208 36235 9210
rect 22369 9152 22374 9208
rect 22430 9152 36174 9208
rect 36230 9152 36235 9208
rect 22369 9150 36235 9152
rect 22369 9147 22435 9150
rect 36169 9147 36235 9150
rect 0 9074 120 9104
rect 3969 9074 4035 9077
rect 0 9072 4035 9074
rect 0 9016 3974 9072
rect 4030 9016 4035 9072
rect 0 9014 4035 9016
rect 0 8984 120 9014
rect 3969 9011 4035 9014
rect 10133 9074 10199 9077
rect 26969 9074 27035 9077
rect 10133 9072 27035 9074
rect 10133 9016 10138 9072
rect 10194 9016 26974 9072
rect 27030 9016 27035 9072
rect 10133 9014 27035 9016
rect 10133 9011 10199 9014
rect 26969 9011 27035 9014
rect 43345 9074 43411 9077
rect 45880 9074 46000 9104
rect 43345 9072 46000 9074
rect 43345 9016 43350 9072
rect 43406 9016 46000 9072
rect 43345 9014 46000 9016
rect 43345 9011 43411 9014
rect 45880 8984 46000 9014
rect 15745 8938 15811 8941
rect 35065 8938 35131 8941
rect 15745 8936 35131 8938
rect 15745 8880 15750 8936
rect 15806 8880 35070 8936
rect 35126 8880 35131 8936
rect 15745 8878 35131 8880
rect 15745 8875 15811 8878
rect 35065 8875 35131 8878
rect 0 8802 120 8832
rect 2589 8802 2655 8805
rect 45880 8802 46000 8832
rect 0 8800 2655 8802
rect 0 8744 2594 8800
rect 2650 8744 2655 8800
rect 0 8742 2655 8744
rect 0 8712 120 8742
rect 2589 8739 2655 8742
rect 43670 8742 46000 8802
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 39006 8671 39322 8672
rect 0 8530 120 8560
rect 30097 8530 30163 8533
rect 0 8528 30163 8530
rect 0 8472 30102 8528
rect 30158 8472 30163 8528
rect 0 8470 30163 8472
rect 0 8440 120 8470
rect 30097 8467 30163 8470
rect 38653 8530 38719 8533
rect 40217 8530 40283 8533
rect 38653 8528 40283 8530
rect 38653 8472 38658 8528
rect 38714 8472 40222 8528
rect 40278 8472 40283 8528
rect 38653 8470 40283 8472
rect 38653 8467 38719 8470
rect 40217 8467 40283 8470
rect 43670 8397 43730 8742
rect 45880 8712 46000 8742
rect 43805 8530 43871 8533
rect 45880 8530 46000 8560
rect 43805 8528 46000 8530
rect 43805 8472 43810 8528
rect 43866 8472 46000 8528
rect 43805 8470 46000 8472
rect 43805 8467 43871 8470
rect 45880 8440 46000 8470
rect 2589 8394 2655 8397
rect 29637 8394 29703 8397
rect 2589 8392 29703 8394
rect 2589 8336 2594 8392
rect 2650 8336 29642 8392
rect 29698 8336 29703 8392
rect 2589 8334 29703 8336
rect 2589 8331 2655 8334
rect 29637 8331 29703 8334
rect 43621 8392 43730 8397
rect 43621 8336 43626 8392
rect 43682 8336 43730 8392
rect 43621 8334 43730 8336
rect 43621 8331 43687 8334
rect 0 8258 120 8288
rect 1761 8258 1827 8261
rect 0 8256 1827 8258
rect 0 8200 1766 8256
rect 1822 8200 1827 8256
rect 0 8198 1827 8200
rect 0 8168 120 8198
rect 1761 8195 1827 8198
rect 20345 8258 20411 8261
rect 25221 8258 25287 8261
rect 20345 8256 25287 8258
rect 20345 8200 20350 8256
rect 20406 8200 25226 8256
rect 25282 8200 25287 8256
rect 20345 8198 25287 8200
rect 20345 8195 20411 8198
rect 25221 8195 25287 8198
rect 44449 8258 44515 8261
rect 45880 8258 46000 8288
rect 44449 8256 46000 8258
rect 44449 8200 44454 8256
rect 44510 8200 46000 8256
rect 44449 8198 46000 8200
rect 44449 8195 44515 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 37946 8127 38262 8128
rect 43946 8192 44262 8193
rect 43946 8128 43952 8192
rect 44016 8128 44032 8192
rect 44096 8128 44112 8192
rect 44176 8128 44192 8192
rect 44256 8128 44262 8192
rect 45880 8168 46000 8198
rect 43946 8127 44262 8128
rect 19793 8122 19859 8125
rect 14414 8120 19859 8122
rect 14414 8064 19798 8120
rect 19854 8064 19859 8120
rect 14414 8062 19859 8064
rect 0 7986 120 8016
rect 1301 7986 1367 7989
rect 0 7984 1367 7986
rect 0 7928 1306 7984
rect 1362 7928 1367 7984
rect 0 7926 1367 7928
rect 0 7896 120 7926
rect 1301 7923 1367 7926
rect 5073 7986 5139 7989
rect 14414 7986 14474 8062
rect 19793 8059 19859 8062
rect 5073 7984 14474 7986
rect 5073 7928 5078 7984
rect 5134 7928 14474 7984
rect 5073 7926 14474 7928
rect 14641 7986 14707 7989
rect 25589 7986 25655 7989
rect 14641 7984 25655 7986
rect 14641 7928 14646 7984
rect 14702 7928 25594 7984
rect 25650 7928 25655 7984
rect 14641 7926 25655 7928
rect 5073 7923 5139 7926
rect 14641 7923 14707 7926
rect 25589 7923 25655 7926
rect 43529 7986 43595 7989
rect 45880 7986 46000 8016
rect 43529 7984 46000 7986
rect 43529 7928 43534 7984
rect 43590 7928 46000 7984
rect 43529 7926 46000 7928
rect 43529 7923 43595 7926
rect 45880 7896 46000 7926
rect 5257 7850 5323 7853
rect 43161 7850 43227 7853
rect 5257 7848 43227 7850
rect 5257 7792 5262 7848
rect 5318 7792 43166 7848
rect 43222 7792 43227 7848
rect 5257 7790 43227 7792
rect 5257 7787 5323 7790
rect 43161 7787 43227 7790
rect 0 7714 120 7744
rect 1117 7714 1183 7717
rect 0 7712 1183 7714
rect 0 7656 1122 7712
rect 1178 7656 1183 7712
rect 0 7654 1183 7656
rect 0 7624 120 7654
rect 1117 7651 1183 7654
rect 44817 7714 44883 7717
rect 45880 7714 46000 7744
rect 44817 7712 46000 7714
rect 44817 7656 44822 7712
rect 44878 7656 46000 7712
rect 44817 7654 46000 7656
rect 44817 7651 44883 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 45880 7624 46000 7654
rect 39006 7583 39322 7584
rect 4705 7578 4771 7581
rect 8569 7578 8635 7581
rect 4705 7576 8635 7578
rect 4705 7520 4710 7576
rect 4766 7520 8574 7576
rect 8630 7520 8635 7576
rect 4705 7518 8635 7520
rect 4705 7515 4771 7518
rect 8569 7515 8635 7518
rect 0 7442 120 7472
rect 21357 7442 21423 7445
rect 0 7440 21423 7442
rect 0 7384 21362 7440
rect 21418 7384 21423 7440
rect 0 7382 21423 7384
rect 0 7352 120 7382
rect 21357 7379 21423 7382
rect 44449 7442 44515 7445
rect 45880 7442 46000 7472
rect 44449 7440 46000 7442
rect 44449 7384 44454 7440
rect 44510 7384 46000 7440
rect 44449 7382 46000 7384
rect 44449 7379 44515 7382
rect 45880 7352 46000 7382
rect 7649 7306 7715 7309
rect 10133 7306 10199 7309
rect 14641 7306 14707 7309
rect 34329 7306 34395 7309
rect 7649 7304 10058 7306
rect 7649 7248 7654 7304
rect 7710 7248 10058 7304
rect 7649 7246 10058 7248
rect 7649 7243 7715 7246
rect 0 7170 120 7200
rect 1025 7170 1091 7173
rect 0 7168 1091 7170
rect 0 7112 1030 7168
rect 1086 7112 1091 7168
rect 0 7110 1091 7112
rect 9998 7170 10058 7246
rect 10133 7304 14707 7306
rect 10133 7248 10138 7304
rect 10194 7248 14646 7304
rect 14702 7248 14707 7304
rect 10133 7246 14707 7248
rect 10133 7243 10199 7246
rect 14641 7243 14707 7246
rect 16530 7304 34395 7306
rect 16530 7248 34334 7304
rect 34390 7248 34395 7304
rect 16530 7246 34395 7248
rect 13721 7170 13787 7173
rect 9998 7168 13787 7170
rect 9998 7112 13726 7168
rect 13782 7112 13787 7168
rect 9998 7110 13787 7112
rect 0 7080 120 7110
rect 1025 7107 1091 7110
rect 13721 7107 13787 7110
rect 14365 7170 14431 7173
rect 16530 7170 16590 7246
rect 34329 7243 34395 7246
rect 14365 7168 16590 7170
rect 14365 7112 14370 7168
rect 14426 7112 16590 7168
rect 14365 7110 16590 7112
rect 44449 7170 44515 7173
rect 45880 7170 46000 7200
rect 44449 7168 46000 7170
rect 44449 7112 44454 7168
rect 44510 7112 46000 7168
rect 44449 7110 46000 7112
rect 14365 7107 14431 7110
rect 44449 7107 44515 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 37946 7039 38262 7040
rect 43946 7104 44262 7105
rect 43946 7040 43952 7104
rect 44016 7040 44032 7104
rect 44096 7040 44112 7104
rect 44176 7040 44192 7104
rect 44256 7040 44262 7104
rect 45880 7080 46000 7110
rect 43946 7039 44262 7040
rect 8569 7034 8635 7037
rect 10133 7034 10199 7037
rect 8569 7032 10199 7034
rect 8569 6976 8574 7032
rect 8630 6976 10138 7032
rect 10194 6976 10199 7032
rect 8569 6974 10199 6976
rect 8569 6971 8635 6974
rect 10133 6971 10199 6974
rect 11094 6972 11100 7036
rect 11164 7034 11170 7036
rect 21541 7034 21607 7037
rect 11164 6974 13738 7034
rect 11164 6972 11170 6974
rect 0 6898 120 6928
rect 9581 6898 9647 6901
rect 0 6896 9647 6898
rect 0 6840 9586 6896
rect 9642 6840 9647 6896
rect 0 6838 9647 6840
rect 13678 6898 13738 6974
rect 14414 6974 19810 7034
rect 14414 6898 14474 6974
rect 13678 6838 14474 6898
rect 19750 6930 19810 6974
rect 20486 7032 21607 7034
rect 20486 6976 21546 7032
rect 21602 6976 21607 7032
rect 20486 6974 21607 6976
rect 20486 6930 20546 6974
rect 21541 6971 21607 6974
rect 19750 6870 20546 6930
rect 44081 6898 44147 6901
rect 45880 6898 46000 6928
rect 44081 6896 46000 6898
rect 44081 6840 44086 6896
rect 44142 6840 46000 6896
rect 44081 6838 46000 6840
rect 0 6808 120 6838
rect 9581 6835 9647 6838
rect 44081 6835 44147 6838
rect 45880 6808 46000 6838
rect 19701 6762 19767 6765
rect 2730 6760 19767 6762
rect 2730 6704 19706 6760
rect 19762 6704 19767 6760
rect 2730 6702 19767 6704
rect 0 6626 120 6656
rect 2730 6626 2790 6702
rect 19701 6699 19767 6702
rect 0 6566 2790 6626
rect 43345 6626 43411 6629
rect 45880 6626 46000 6656
rect 43345 6624 46000 6626
rect 43345 6568 43350 6624
rect 43406 6568 46000 6624
rect 43345 6566 46000 6568
rect 0 6536 120 6566
rect 43345 6563 43411 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 45880 6536 46000 6566
rect 39006 6495 39322 6496
rect 0 6354 120 6384
rect 5533 6354 5599 6357
rect 0 6352 5599 6354
rect 0 6296 5538 6352
rect 5594 6296 5599 6352
rect 0 6294 5599 6296
rect 0 6264 120 6294
rect 5533 6291 5599 6294
rect 7833 6354 7899 6357
rect 42977 6354 43043 6357
rect 45880 6354 46000 6384
rect 7833 6352 16590 6354
rect 7833 6296 7838 6352
rect 7894 6296 16590 6352
rect 7833 6294 16590 6296
rect 7833 6291 7899 6294
rect 13721 6218 13787 6221
rect 1718 6216 13787 6218
rect 1718 6160 13726 6216
rect 13782 6160 13787 6216
rect 1718 6158 13787 6160
rect 16530 6218 16590 6294
rect 42977 6352 46000 6354
rect 42977 6296 42982 6352
rect 43038 6296 46000 6352
rect 42977 6294 46000 6296
rect 42977 6291 43043 6294
rect 45880 6264 46000 6294
rect 34973 6218 35039 6221
rect 16530 6216 35039 6218
rect 16530 6160 34978 6216
rect 35034 6160 35039 6216
rect 16530 6158 35039 6160
rect 0 6082 120 6112
rect 1718 6082 1778 6158
rect 13721 6155 13787 6158
rect 34973 6155 35039 6158
rect 0 6022 1778 6082
rect 44449 6082 44515 6085
rect 45880 6082 46000 6112
rect 44449 6080 46000 6082
rect 44449 6024 44454 6080
rect 44510 6024 46000 6080
rect 44449 6022 46000 6024
rect 0 5992 120 6022
rect 44449 6019 44515 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 37946 5951 38262 5952
rect 43946 6016 44262 6017
rect 43946 5952 43952 6016
rect 44016 5952 44032 6016
rect 44096 5952 44112 6016
rect 44176 5952 44192 6016
rect 44256 5952 44262 6016
rect 45880 5992 46000 6022
rect 43946 5951 44262 5952
rect 0 5810 120 5840
rect 24669 5810 24735 5813
rect 0 5808 24735 5810
rect 0 5752 24674 5808
rect 24730 5752 24735 5808
rect 0 5750 24735 5752
rect 0 5720 120 5750
rect 24669 5747 24735 5750
rect 27521 5810 27587 5813
rect 35801 5810 35867 5813
rect 27521 5808 35867 5810
rect 27521 5752 27526 5808
rect 27582 5752 35806 5808
rect 35862 5752 35867 5808
rect 27521 5750 35867 5752
rect 27521 5747 27587 5750
rect 35801 5747 35867 5750
rect 43713 5810 43779 5813
rect 45880 5810 46000 5840
rect 43713 5808 46000 5810
rect 43713 5752 43718 5808
rect 43774 5752 46000 5808
rect 43713 5750 46000 5752
rect 43713 5747 43779 5750
rect 45880 5720 46000 5750
rect 15285 5674 15351 5677
rect 44265 5674 44331 5677
rect 2822 5614 3618 5674
rect 0 5538 120 5568
rect 2822 5538 2882 5614
rect 0 5478 2882 5538
rect 3558 5538 3618 5614
rect 15285 5672 44331 5674
rect 15285 5616 15290 5672
rect 15346 5616 44270 5672
rect 44326 5616 44331 5672
rect 15285 5614 44331 5616
rect 15285 5611 15351 5614
rect 44265 5611 44331 5614
rect 9397 5538 9463 5541
rect 14549 5538 14615 5541
rect 3558 5478 7850 5538
rect 0 5448 120 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 0 5266 120 5296
rect 7790 5266 7850 5478
rect 9397 5536 14615 5538
rect 9397 5480 9402 5536
rect 9458 5480 14554 5536
rect 14610 5480 14615 5536
rect 9397 5478 14615 5480
rect 9397 5475 9463 5478
rect 14549 5475 14615 5478
rect 44357 5538 44423 5541
rect 45880 5538 46000 5568
rect 44357 5536 46000 5538
rect 44357 5480 44362 5536
rect 44418 5480 46000 5536
rect 44357 5478 46000 5480
rect 44357 5475 44423 5478
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 45880 5448 46000 5478
rect 39006 5407 39322 5408
rect 19149 5266 19215 5269
rect 0 5206 7666 5266
rect 7790 5264 19215 5266
rect 7790 5208 19154 5264
rect 19210 5208 19215 5264
rect 7790 5206 19215 5208
rect 0 5176 120 5206
rect 7606 5130 7666 5206
rect 19149 5203 19215 5206
rect 20529 5266 20595 5269
rect 43161 5266 43227 5269
rect 20529 5264 43227 5266
rect 20529 5208 20534 5264
rect 20590 5208 43166 5264
rect 43222 5208 43227 5264
rect 20529 5206 43227 5208
rect 20529 5203 20595 5206
rect 43161 5203 43227 5206
rect 44449 5266 44515 5269
rect 45880 5266 46000 5296
rect 44449 5264 46000 5266
rect 44449 5208 44454 5264
rect 44510 5208 46000 5264
rect 44449 5206 46000 5208
rect 44449 5203 44515 5206
rect 45880 5176 46000 5206
rect 14549 5130 14615 5133
rect 33501 5130 33567 5133
rect 1718 5070 2790 5130
rect 7606 5070 14474 5130
rect 0 4994 120 5024
rect 1718 4994 1778 5070
rect 0 4934 1778 4994
rect 2730 4994 2790 5070
rect 7741 4994 7807 4997
rect 2730 4992 7807 4994
rect 2730 4936 7746 4992
rect 7802 4936 7807 4992
rect 2730 4934 7807 4936
rect 14414 4994 14474 5070
rect 14549 5128 33567 5130
rect 14549 5072 14554 5128
rect 14610 5072 33506 5128
rect 33562 5072 33567 5128
rect 14549 5070 33567 5072
rect 14549 5067 14615 5070
rect 33501 5067 33567 5070
rect 44081 5130 44147 5133
rect 44081 5128 45018 5130
rect 44081 5072 44086 5128
rect 44142 5072 45018 5128
rect 44081 5070 45018 5072
rect 44081 5067 44147 5070
rect 16757 4994 16823 4997
rect 14414 4992 16823 4994
rect 14414 4936 16762 4992
rect 16818 4936 16823 4992
rect 14414 4934 16823 4936
rect 44958 4994 45018 5070
rect 45880 4994 46000 5024
rect 44958 4934 46000 4994
rect 0 4904 120 4934
rect 7741 4931 7807 4934
rect 16757 4931 16823 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 37946 4863 38262 4864
rect 43946 4928 44262 4929
rect 43946 4864 43952 4928
rect 44016 4864 44032 4928
rect 44096 4864 44112 4928
rect 44176 4864 44192 4928
rect 44256 4864 44262 4928
rect 45880 4904 46000 4934
rect 43946 4863 44262 4864
rect 7649 4858 7715 4861
rect 2730 4856 7715 4858
rect 2730 4800 7654 4856
rect 7710 4800 7715 4856
rect 2730 4798 7715 4800
rect 0 4722 120 4752
rect 2730 4722 2790 4798
rect 7649 4795 7715 4798
rect 8385 4858 8451 4861
rect 11094 4858 11100 4860
rect 8385 4856 11100 4858
rect 8385 4800 8390 4856
rect 8446 4800 11100 4856
rect 8385 4798 11100 4800
rect 8385 4795 8451 4798
rect 11094 4796 11100 4798
rect 11164 4796 11170 4860
rect 0 4662 2790 4722
rect 2865 4722 2931 4725
rect 7925 4722 7991 4725
rect 16665 4722 16731 4725
rect 2865 4720 7850 4722
rect 2865 4664 2870 4720
rect 2926 4664 7850 4720
rect 2865 4662 7850 4664
rect 0 4632 120 4662
rect 2865 4659 2931 4662
rect 7790 4586 7850 4662
rect 7925 4720 16731 4722
rect 7925 4664 7930 4720
rect 7986 4664 16670 4720
rect 16726 4664 16731 4720
rect 7925 4662 16731 4664
rect 7925 4659 7991 4662
rect 16665 4659 16731 4662
rect 44449 4722 44515 4725
rect 45880 4722 46000 4752
rect 44449 4720 46000 4722
rect 44449 4664 44454 4720
rect 44510 4664 46000 4720
rect 44449 4662 46000 4664
rect 44449 4659 44515 4662
rect 45880 4632 46000 4662
rect 40769 4586 40835 4589
rect 2730 4526 7666 4586
rect 7790 4584 40835 4586
rect 7790 4528 40774 4584
rect 40830 4528 40835 4584
rect 7790 4526 40835 4528
rect 0 4450 120 4480
rect 2730 4450 2790 4526
rect 0 4390 2790 4450
rect 0 4360 120 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 1301 4314 1367 4317
rect 2865 4314 2931 4317
rect 1301 4312 2931 4314
rect 1301 4256 1306 4312
rect 1362 4256 2870 4312
rect 2926 4256 2931 4312
rect 1301 4254 2931 4256
rect 1301 4251 1367 4254
rect 2865 4251 2931 4254
rect 0 4178 120 4208
rect 7465 4178 7531 4181
rect 0 4176 7531 4178
rect 0 4120 7470 4176
rect 7526 4120 7531 4176
rect 0 4118 7531 4120
rect 7606 4178 7666 4526
rect 40769 4523 40835 4526
rect 44081 4450 44147 4453
rect 45880 4450 46000 4480
rect 44081 4448 46000 4450
rect 44081 4392 44086 4448
rect 44142 4392 46000 4448
rect 44081 4390 46000 4392
rect 44081 4387 44147 4390
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 45880 4360 46000 4390
rect 39006 4319 39322 4320
rect 20713 4178 20779 4181
rect 7606 4118 14658 4178
rect 0 4088 120 4118
rect 7465 4115 7531 4118
rect 14598 4042 14658 4118
rect 19566 4176 20779 4178
rect 19566 4120 20718 4176
rect 20774 4120 20779 4176
rect 19566 4118 20779 4120
rect 19566 4042 19626 4118
rect 20713 4115 20779 4118
rect 44449 4178 44515 4181
rect 45880 4178 46000 4208
rect 44449 4176 46000 4178
rect 44449 4120 44454 4176
rect 44510 4120 46000 4176
rect 44449 4118 46000 4120
rect 44449 4115 44515 4118
rect 45880 4088 46000 4118
rect 23657 4042 23723 4045
rect 42885 4042 42951 4045
rect 1718 3982 14474 4042
rect 14598 3982 19626 4042
rect 19750 3982 22110 4042
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 0 3846 1778 3906
rect 14414 3906 14474 3982
rect 19750 3906 19810 3982
rect 14414 3846 19810 3906
rect 22050 3906 22110 3982
rect 23657 4040 42951 4042
rect 23657 3984 23662 4040
rect 23718 3984 42890 4040
rect 42946 3984 42951 4040
rect 23657 3982 42951 3984
rect 23657 3979 23723 3982
rect 42885 3979 42951 3982
rect 44081 4042 44147 4045
rect 44081 4040 45018 4042
rect 44081 3984 44086 4040
rect 44142 3984 45018 4040
rect 44081 3982 45018 3984
rect 44081 3979 44147 3982
rect 25589 3906 25655 3909
rect 22050 3904 25655 3906
rect 22050 3848 25594 3904
rect 25650 3848 25655 3904
rect 22050 3846 25655 3848
rect 44958 3906 45018 3982
rect 45880 3906 46000 3936
rect 44958 3846 46000 3906
rect 0 3816 120 3846
rect 25589 3843 25655 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 37946 3775 38262 3776
rect 43946 3840 44262 3841
rect 43946 3776 43952 3840
rect 44016 3776 44032 3840
rect 44096 3776 44112 3840
rect 44176 3776 44192 3840
rect 44256 3776 44262 3840
rect 45880 3816 46000 3846
rect 43946 3775 44262 3776
rect 0 3634 120 3664
rect 14273 3634 14339 3637
rect 0 3632 14339 3634
rect 0 3576 14278 3632
rect 14334 3576 14339 3632
rect 0 3574 14339 3576
rect 0 3544 120 3574
rect 14273 3571 14339 3574
rect 24577 3634 24643 3637
rect 42793 3634 42859 3637
rect 24577 3632 42859 3634
rect 24577 3576 24582 3632
rect 24638 3576 42798 3632
rect 42854 3576 42859 3632
rect 24577 3574 42859 3576
rect 24577 3571 24643 3574
rect 42793 3571 42859 3574
rect 44449 3634 44515 3637
rect 45880 3634 46000 3664
rect 44449 3632 46000 3634
rect 44449 3576 44454 3632
rect 44510 3576 46000 3632
rect 44449 3574 46000 3576
rect 44449 3571 44515 3574
rect 45880 3544 46000 3574
rect 7465 3498 7531 3501
rect 24209 3498 24275 3501
rect 2730 3438 3618 3498
rect 0 3362 120 3392
rect 2730 3362 2790 3438
rect 0 3302 2790 3362
rect 3558 3362 3618 3438
rect 7465 3496 24275 3498
rect 7465 3440 7470 3496
rect 7526 3440 24214 3496
rect 24270 3440 24275 3496
rect 7465 3438 24275 3440
rect 7465 3435 7531 3438
rect 24209 3435 24275 3438
rect 24853 3498 24919 3501
rect 40033 3498 40099 3501
rect 24853 3496 40099 3498
rect 24853 3440 24858 3496
rect 24914 3440 40038 3496
rect 40094 3440 40099 3496
rect 24853 3438 40099 3440
rect 24853 3435 24919 3438
rect 40033 3435 40099 3438
rect 8385 3362 8451 3365
rect 3558 3360 8451 3362
rect 3558 3304 8390 3360
rect 8446 3304 8451 3360
rect 3558 3302 8451 3304
rect 0 3272 120 3302
rect 8385 3299 8451 3302
rect 44081 3362 44147 3365
rect 45880 3362 46000 3392
rect 44081 3360 46000 3362
rect 44081 3304 44086 3360
rect 44142 3304 46000 3360
rect 44081 3302 46000 3304
rect 44081 3299 44147 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 45880 3272 46000 3302
rect 39006 3231 39322 3232
rect 23289 3226 23355 3229
rect 21958 3224 23355 3226
rect 21958 3168 23294 3224
rect 23350 3168 23355 3224
rect 21958 3166 23355 3168
rect 0 3090 120 3120
rect 21958 3090 22018 3166
rect 23289 3163 23355 3166
rect 0 3030 22018 3090
rect 22185 3090 22251 3093
rect 25865 3090 25931 3093
rect 42609 3090 42675 3093
rect 22185 3088 25698 3090
rect 22185 3032 22190 3088
rect 22246 3032 25698 3088
rect 22185 3030 25698 3032
rect 0 3000 120 3030
rect 22185 3027 22251 3030
rect 24209 2954 24275 2957
rect 1718 2952 24275 2954
rect 1718 2896 24214 2952
rect 24270 2896 24275 2952
rect 1718 2894 24275 2896
rect 25638 2954 25698 3030
rect 25865 3088 42675 3090
rect 25865 3032 25870 3088
rect 25926 3032 42614 3088
rect 42670 3032 42675 3088
rect 25865 3030 42675 3032
rect 25865 3027 25931 3030
rect 42609 3027 42675 3030
rect 44449 3090 44515 3093
rect 45880 3090 46000 3120
rect 44449 3088 46000 3090
rect 44449 3032 44454 3088
rect 44510 3032 46000 3088
rect 44449 3030 46000 3032
rect 44449 3027 44515 3030
rect 45880 3000 46000 3030
rect 40125 2954 40191 2957
rect 25638 2952 40191 2954
rect 25638 2896 40130 2952
rect 40186 2896 40191 2952
rect 25638 2894 40191 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 24209 2891 24275 2894
rect 40125 2891 40191 2894
rect 44081 2954 44147 2957
rect 44081 2952 45018 2954
rect 44081 2896 44086 2952
rect 44142 2896 45018 2952
rect 44081 2894 45018 2896
rect 44081 2891 44147 2894
rect 0 2758 1778 2818
rect 8385 2818 8451 2821
rect 12433 2818 12499 2821
rect 8385 2816 12499 2818
rect 8385 2760 8390 2816
rect 8446 2760 12438 2816
rect 12494 2760 12499 2816
rect 8385 2758 12499 2760
rect 44958 2818 45018 2894
rect 45880 2818 46000 2848
rect 44958 2758 46000 2818
rect 0 2728 120 2758
rect 8385 2755 8451 2758
rect 12433 2755 12499 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 37946 2687 38262 2688
rect 43946 2752 44262 2753
rect 43946 2688 43952 2752
rect 44016 2688 44032 2752
rect 44096 2688 44112 2752
rect 44176 2688 44192 2752
rect 44256 2688 44262 2752
rect 45880 2728 46000 2758
rect 43946 2687 44262 2688
rect 0 2546 120 2576
rect 27705 2546 27771 2549
rect 0 2544 27771 2546
rect 0 2488 27710 2544
rect 27766 2488 27771 2544
rect 0 2486 27771 2488
rect 0 2456 120 2486
rect 27705 2483 27771 2486
rect 44449 2546 44515 2549
rect 45880 2546 46000 2576
rect 44449 2544 46000 2546
rect 44449 2488 44454 2544
rect 44510 2488 46000 2544
rect 44449 2486 46000 2488
rect 44449 2483 44515 2486
rect 45880 2456 46000 2486
rect 17677 2410 17743 2413
rect 2822 2408 17743 2410
rect 2822 2352 17682 2408
rect 17738 2352 17743 2408
rect 2822 2350 17743 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 17677 2347 17743 2350
rect 0 2214 2882 2274
rect 44081 2274 44147 2277
rect 45880 2274 46000 2304
rect 44081 2272 46000 2274
rect 44081 2216 44086 2272
rect 44142 2216 46000 2272
rect 44081 2214 46000 2216
rect 0 2184 120 2214
rect 44081 2211 44147 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 45880 2184 46000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 20437 2002 20503 2005
rect 0 2000 20503 2002
rect 0 1944 20442 2000
rect 20498 1944 20503 2000
rect 0 1942 20503 1944
rect 0 1912 120 1942
rect 20437 1939 20503 1942
rect 44817 2002 44883 2005
rect 45880 2002 46000 2032
rect 44817 2000 46000 2002
rect 44817 1944 44822 2000
rect 44878 1944 46000 2000
rect 44817 1942 46000 1944
rect 44817 1939 44883 1942
rect 45880 1912 46000 1942
rect 0 1730 120 1760
rect 19517 1730 19583 1733
rect 0 1728 19583 1730
rect 0 1672 19522 1728
rect 19578 1672 19583 1728
rect 0 1670 19583 1672
rect 0 1640 120 1670
rect 19517 1667 19583 1670
rect 42977 1730 43043 1733
rect 45880 1730 46000 1760
rect 42977 1728 46000 1730
rect 42977 1672 42982 1728
rect 43038 1672 46000 1728
rect 42977 1670 46000 1672
rect 42977 1667 43043 1670
rect 45880 1640 46000 1670
rect 0 1458 120 1488
rect 15745 1458 15811 1461
rect 0 1456 15811 1458
rect 0 1400 15750 1456
rect 15806 1400 15811 1456
rect 0 1398 15811 1400
rect 0 1368 120 1398
rect 15745 1395 15811 1398
rect 43345 1458 43411 1461
rect 45880 1458 46000 1488
rect 43345 1456 46000 1458
rect 43345 1400 43350 1456
rect 43406 1400 46000 1456
rect 43345 1398 46000 1400
rect 43345 1395 43411 1398
rect 45880 1368 46000 1398
rect 33409 1322 33475 1325
rect 35617 1322 35683 1325
rect 33409 1320 35683 1322
rect 33409 1264 33414 1320
rect 33470 1264 35622 1320
rect 35678 1264 35683 1320
rect 33409 1262 35683 1264
rect 33409 1259 33475 1262
rect 35617 1259 35683 1262
rect 0 1186 120 1216
rect 1393 1186 1459 1189
rect 0 1184 1459 1186
rect 0 1128 1398 1184
rect 1454 1128 1459 1184
rect 0 1126 1459 1128
rect 0 1096 120 1126
rect 1393 1123 1459 1126
rect 44357 1186 44423 1189
rect 45880 1186 46000 1216
rect 44357 1184 46000 1186
rect 44357 1128 44362 1184
rect 44418 1128 46000 1184
rect 44357 1126 46000 1128
rect 44357 1123 44423 1126
rect 45880 1096 46000 1126
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 43952 8188 44016 8192
rect 43952 8132 43956 8188
rect 43956 8132 44012 8188
rect 44012 8132 44016 8188
rect 43952 8128 44016 8132
rect 44032 8188 44096 8192
rect 44032 8132 44036 8188
rect 44036 8132 44092 8188
rect 44092 8132 44096 8188
rect 44032 8128 44096 8132
rect 44112 8188 44176 8192
rect 44112 8132 44116 8188
rect 44116 8132 44172 8188
rect 44172 8132 44176 8188
rect 44112 8128 44176 8132
rect 44192 8188 44256 8192
rect 44192 8132 44196 8188
rect 44196 8132 44252 8188
rect 44252 8132 44256 8188
rect 44192 8128 44256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 43952 7100 44016 7104
rect 43952 7044 43956 7100
rect 43956 7044 44012 7100
rect 44012 7044 44016 7100
rect 43952 7040 44016 7044
rect 44032 7100 44096 7104
rect 44032 7044 44036 7100
rect 44036 7044 44092 7100
rect 44092 7044 44096 7100
rect 44032 7040 44096 7044
rect 44112 7100 44176 7104
rect 44112 7044 44116 7100
rect 44116 7044 44172 7100
rect 44172 7044 44176 7100
rect 44112 7040 44176 7044
rect 44192 7100 44256 7104
rect 44192 7044 44196 7100
rect 44196 7044 44252 7100
rect 44252 7044 44256 7100
rect 44192 7040 44256 7044
rect 11100 6972 11164 7036
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 43952 6012 44016 6016
rect 43952 5956 43956 6012
rect 43956 5956 44012 6012
rect 44012 5956 44016 6012
rect 43952 5952 44016 5956
rect 44032 6012 44096 6016
rect 44032 5956 44036 6012
rect 44036 5956 44092 6012
rect 44092 5956 44096 6012
rect 44032 5952 44096 5956
rect 44112 6012 44176 6016
rect 44112 5956 44116 6012
rect 44116 5956 44172 6012
rect 44172 5956 44176 6012
rect 44112 5952 44176 5956
rect 44192 6012 44256 6016
rect 44192 5956 44196 6012
rect 44196 5956 44252 6012
rect 44252 5956 44256 6012
rect 44192 5952 44256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 43952 4924 44016 4928
rect 43952 4868 43956 4924
rect 43956 4868 44012 4924
rect 44012 4868 44016 4924
rect 43952 4864 44016 4868
rect 44032 4924 44096 4928
rect 44032 4868 44036 4924
rect 44036 4868 44092 4924
rect 44092 4868 44096 4924
rect 44032 4864 44096 4868
rect 44112 4924 44176 4928
rect 44112 4868 44116 4924
rect 44116 4868 44172 4924
rect 44172 4868 44176 4924
rect 44112 4864 44176 4868
rect 44192 4924 44256 4928
rect 44192 4868 44196 4924
rect 44196 4868 44252 4924
rect 44252 4868 44256 4924
rect 44192 4864 44256 4868
rect 11100 4796 11164 4860
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 43952 3836 44016 3840
rect 43952 3780 43956 3836
rect 43956 3780 44012 3836
rect 44012 3780 44016 3836
rect 43952 3776 44016 3780
rect 44032 3836 44096 3840
rect 44032 3780 44036 3836
rect 44036 3780 44092 3836
rect 44092 3780 44096 3836
rect 44032 3776 44096 3780
rect 44112 3836 44176 3840
rect 44112 3780 44116 3836
rect 44116 3780 44172 3836
rect 44172 3780 44176 3836
rect 44112 3776 44176 3780
rect 44192 3836 44256 3840
rect 44192 3780 44196 3836
rect 44196 3780 44252 3836
rect 44252 3780 44256 3836
rect 44192 3776 44256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 43952 2748 44016 2752
rect 43952 2692 43956 2748
rect 43956 2692 44012 2748
rect 44012 2692 44016 2748
rect 43952 2688 44016 2692
rect 44032 2748 44096 2752
rect 44032 2692 44036 2748
rect 44036 2692 44092 2748
rect 44092 2692 44096 2748
rect 44032 2688 44096 2692
rect 44112 2748 44176 2752
rect 44112 2692 44116 2748
rect 44116 2692 44172 2748
rect 44172 2692 44176 2748
rect 44112 2688 44176 2692
rect 44192 2748 44256 2752
rect 44192 2692 44196 2748
rect 44196 2692 44252 2748
rect 44252 2692 44256 2748
rect 44192 2688 44256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
<< metal4 >>
rect 1944 8192 2264 11152
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11152
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11152
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11152
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 13944 8192 14264 11152
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 11099 7036 11165 7037
rect 11099 6972 11100 7036
rect 11164 6972 11165 7036
rect 11099 6971 11165 6972
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 11102 4861 11162 6971
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 11099 4860 11165 4861
rect 11099 4796 11100 4860
rect 11164 4796 11165 4860
rect 11099 4795 11165 4796
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11152
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11152
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11152
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11152
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11152
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11152
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11152
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11152
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11152
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
rect 43944 8192 44264 11152
rect 43944 8128 43952 8192
rect 44016 8128 44032 8192
rect 44096 8128 44112 8192
rect 44176 8128 44192 8192
rect 44256 8128 44264 8192
rect 43944 7104 44264 8128
rect 43944 7040 43952 7104
rect 44016 7040 44032 7104
rect 44096 7040 44112 7104
rect 44176 7040 44192 7104
rect 44256 7040 44264 7104
rect 43944 6016 44264 7040
rect 43944 5952 43952 6016
rect 44016 5952 44032 6016
rect 44096 5952 44112 6016
rect 44176 5952 44192 6016
rect 44256 5952 44264 6016
rect 43944 4928 44264 5952
rect 43944 4864 43952 4928
rect 44016 4864 44032 4928
rect 44096 4864 44112 4928
rect 44176 4864 44192 4928
rect 44256 4864 44264 4928
rect 43944 3840 44264 4864
rect 43944 3776 43952 3840
rect 44016 3776 44032 3840
rect 44096 3776 44112 3840
rect 44176 3776 44192 3840
rect 44256 3776 44264 3840
rect 43944 2752 44264 3776
rect 43944 2688 43952 2752
rect 44016 2688 44032 2752
rect 44096 2688 44112 2752
rect 44176 2688 44192 2752
rect 44256 2688 44264 2752
rect 43944 0 44264 2688
use sky130_fd_sc_hd__clkbuf_2  _000_
timestamp -3599
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform 1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _003_
timestamp -3599
transform -1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _004_
timestamp -3599
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _005_
timestamp -3599
transform 1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform 1 0 24380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _009_
timestamp -3599
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 25760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 24380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _014_
timestamp -3599
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _015_
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 20240 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 27048 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _018_
timestamp -3599
transform 1 0 14996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 25484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _021_
timestamp -3599
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _022_
timestamp -3599
transform -1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _023_
timestamp -3599
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _024_
timestamp -3599
transform -1 0 41216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _025_
timestamp -3599
transform -1 0 41216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _026_
timestamp -3599
transform -1 0 36708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 30268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 29716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _029_
timestamp -3599
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 26680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp -3599
transform -1 0 42320 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp -3599
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp -3599
transform -1 0 38364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _034_
timestamp -3599
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _035_
timestamp -3599
transform 1 0 9752 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _036_
timestamp -3599
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _037_
timestamp -3599
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _038_
timestamp -3599
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _039_
timestamp -3599
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform -1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _041_
timestamp -3599
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _042_
timestamp -3599
transform 1 0 26496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform -1 0 40112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _044_
timestamp -3599
transform 1 0 30636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform -1 0 40848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform -1 0 41400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _047_
timestamp -3599
transform 1 0 29900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform -1 0 37812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform -1 0 41308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 42780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 42780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp -3599
transform -1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp -3599
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp -3599
transform -1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp -3599
transform -1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp -3599
transform -1 0 21620 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _057_
timestamp -3599
transform -1 0 20424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp -3599
transform -1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp -3599
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp -3599
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp -3599
transform -1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp -3599
transform -1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _063_
timestamp -3599
transform -1 0 16468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp -3599
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _065_
timestamp -3599
transform -1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp -3599
transform -1 0 25484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _067_
timestamp -3599
transform -1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp -3599
transform -1 0 24288 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _069_
timestamp -3599
transform -1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _070_
timestamp -3599
transform -1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _071_
timestamp -3599
transform -1 0 22724 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _072_
timestamp -3599
transform -1 0 34592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp -3599
transform -1 0 35328 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _074_
timestamp -3599
transform -1 0 34408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _075_
timestamp -3599
transform -1 0 33764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _076_
timestamp -3599
transform -1 0 33304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _077_
timestamp -3599
transform -1 0 32384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _078_
timestamp -3599
transform -1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _079_
timestamp -3599
transform -1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _080_
timestamp -3599
transform -1 0 28428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _081_
timestamp -3599
transform -1 0 28520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _082_
timestamp -3599
transform -1 0 28704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _083_
timestamp -3599
transform -1 0 27876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform -1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform -1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform -1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp -3599
transform -1 0 27232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform -1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform -1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform -1 0 12696 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp -3599
transform -1 0 12972 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp -3599
transform -1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp -3599
transform -1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp -3599
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp -3599
transform -1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp -3599
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp -3599
transform -1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform -1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp -3599
transform 1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _100_
timestamp -3599
transform -1 0 38272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _101_
timestamp -3599
transform -1 0 36248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp -3599
transform -1 0 36432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _103_
timestamp -3599
transform -1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform 1 0 36156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 25576 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 24380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 21712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform 1 0 20056 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 27508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform 1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 15732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 20240 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 10948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform 1 0 40756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform 1 0 30084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 19688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform 1 0 26496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform -1 0 42044 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform 1 0 17664 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform 1 0 27692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform 1 0 24196 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform 1 0 23276 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 27416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 19780 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 10212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 13340 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform -1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform -1 0 17848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform -1 0 17020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp -3599
transform -1 0 15272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp -3599
transform -1 0 10948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6
timestamp -3599
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp -3599
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12
timestamp -3599
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18
timestamp -3599
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21
timestamp -3599
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp -3599
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35
timestamp -3599
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp -3599
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp -3599
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47
timestamp -3599
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50
timestamp -3599
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60
timestamp -3599
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp -3599
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp -3599
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp -3599
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78
timestamp -3599
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_88
timestamp -3599
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91
timestamp -3599
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp -3599
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp -3599
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100
timestamp -3599
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103
timestamp -3599
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106
timestamp -3599
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_116
timestamp -3599
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp -3599
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_122
timestamp -3599
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp -3599
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_128
timestamp -3599
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_131
timestamp -3599
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_134
timestamp -3599
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_144
timestamp -3599
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_147
timestamp -3599
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_150
timestamp -3599
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_153
timestamp -3599
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp -3599
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_159
timestamp -3599
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_162
timestamp -3599
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_172
timestamp -3599
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_175
timestamp -3599
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_178
timestamp -3599
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp -3599
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_184
timestamp -3599
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp -3599
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_190
timestamp -3599
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_200
timestamp -3599
transform 1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_203
timestamp -3599
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_206
timestamp -3599
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_209
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_212
timestamp -3599
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_215
timestamp -3599
transform 1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp -3599
transform 1 0 21160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_228
timestamp -3599
transform 1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_231
timestamp -3599
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_234
timestamp -3599
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_237
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_240
timestamp -3599
transform 1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_243
timestamp -3599
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_246
timestamp -3599
transform 1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_256
timestamp -3599
transform 1 0 24656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_259
timestamp -3599
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_262
timestamp -3599
transform 1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_265
timestamp -3599
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_268
timestamp -3599
transform 1 0 25760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_271
timestamp -3599
transform 1 0 26036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_274
timestamp -3599
transform 1 0 26312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_281
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_284
timestamp -3599
transform 1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_287
timestamp -3599
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_290
timestamp -3599
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_293
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp -3599
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_299
timestamp -3599
transform 1 0 28612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_302
timestamp -3599
transform 1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_312
timestamp -3599
transform 1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_315
timestamp -3599
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_318
timestamp -3599
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_321
timestamp -3599
transform 1 0 30636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_324
timestamp -3599
transform 1 0 30912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_327
timestamp -3599
transform 1 0 31188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_330
timestamp -3599
transform 1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_337
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_340
timestamp -3599
transform 1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_343
timestamp -3599
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_346
timestamp -3599
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_349
timestamp -3599
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_352
timestamp -3599
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_355
timestamp -3599
transform 1 0 33764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_358
timestamp -3599
transform 1 0 34040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_365
timestamp -3599
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_368
timestamp -3599
transform 1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_371
timestamp -3599
transform 1 0 35236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_374
timestamp -3599
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp -3599
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_380
timestamp -3599
transform 1 0 36064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_383
timestamp -3599
transform 1 0 36340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_386
timestamp -3599
transform 1 0 36616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_396
timestamp -3599
transform 1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_399
timestamp -3599
transform 1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_402
timestamp -3599
transform 1 0 38088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_405
timestamp -3599
transform 1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_408
timestamp -3599
transform 1 0 38640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_411
timestamp -3599
transform 1 0 38916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_414
timestamp -3599
transform 1 0 39192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp -3599
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_421
timestamp -3599
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_424
timestamp -3599
transform 1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_427
timestamp -3599
transform 1 0 40388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_430
timestamp -3599
transform 1 0 40664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_433
timestamp -3599
transform 1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_436
timestamp -3599
transform 1 0 41216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_439
timestamp -3599
transform 1 0 41492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_442
timestamp -3599
transform 1 0 41768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp -3599
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_449
timestamp -3599
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_452
timestamp -3599
transform 1 0 42688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6
timestamp -3599
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_13
timestamp -3599
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_16
timestamp -3599
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_19
timestamp -3599
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_22
timestamp -3599
transform 1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_25
timestamp -3599
transform 1 0 3404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_28
timestamp -3599
transform 1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_31
timestamp -3599
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_34
timestamp -3599
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_37
timestamp -3599
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_40
timestamp -3599
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_43
timestamp -3599
transform 1 0 5060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_46
timestamp -3599
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_49
timestamp -3599
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_52
timestamp -3599
transform 1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_60
timestamp -3599
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_63
timestamp -3599
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_66
timestamp -3599
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp -3599
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp -3599
transform 1 0 7728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp -3599
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp -3599
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_84
timestamp -3599
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_87
timestamp -3599
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_90
timestamp -3599
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_93
timestamp -3599
transform 1 0 9660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_98
timestamp -3599
transform 1 0 10120 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_101
timestamp -3599
transform 1 0 10396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_104
timestamp -3599
transform 1 0 10672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_116
timestamp -3599
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_119
timestamp -3599
transform 1 0 12052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp -3599
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_128
timestamp -3599
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_131
timestamp -3599
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_134
timestamp -3599
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_137
timestamp -3599
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_140
timestamp -3599
transform 1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp -3599
transform 1 0 14260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_146
timestamp -3599
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_153
timestamp -3599
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_156
timestamp -3599
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_164
timestamp -3599
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_172
timestamp -3599
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_175
timestamp -3599
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp -3599
transform 1 0 17480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_188
timestamp -3599
transform 1 0 18400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_191
timestamp -3599
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_194
timestamp -3599
transform 1 0 18952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_197
timestamp -3599
transform 1 0 19228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_200
timestamp -3599
transform 1 0 19504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_203
timestamp -3599
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_211
timestamp -3599
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_214
timestamp -3599
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_217
timestamp -3599
transform 1 0 21068 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_228
timestamp -3599
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_231
timestamp -3599
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_234
timestamp -3599
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_237
timestamp -3599
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_240
timestamp -3599
transform 1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_243
timestamp -3599
transform 1 0 23460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_246
timestamp -3599
transform 1 0 23736 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_250
timestamp -3599
transform 1 0 24104 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_256
timestamp -3599
transform 1 0 24656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_259
timestamp -3599
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_262
timestamp -3599
transform 1 0 25208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_268
timestamp -3599
transform 1 0 25760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_271
timestamp -3599
transform 1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_274
timestamp -3599
transform 1 0 26312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_284
timestamp -3599
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_287
timestamp -3599
transform 1 0 27508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_294
timestamp -3599
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_297
timestamp -3599
transform 1 0 28428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_300
timestamp -3599
transform 1 0 28704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_303
timestamp -3599
transform 1 0 28980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_306
timestamp -3599
transform 1 0 29256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_309
timestamp -3599
transform 1 0 29532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_312
timestamp -3599
transform 1 0 29808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_315
timestamp -3599
transform 1 0 30084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_318
timestamp -3599
transform 1 0 30360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_324
timestamp -3599
transform 1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_327
timestamp -3599
transform 1 0 31188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_330
timestamp -3599
transform 1 0 31464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp -3599
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_340
timestamp -3599
transform 1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_343
timestamp -3599
transform 1 0 32660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_346
timestamp -3599
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_349
timestamp -3599
transform 1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_352
timestamp -3599
transform 1 0 33488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_355
timestamp -3599
transform 1 0 33764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_358
timestamp -3599
transform 1 0 34040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_361
timestamp -3599
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_364
timestamp -3599
transform 1 0 34592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_367
timestamp -3599
transform 1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_370
timestamp -3599
transform 1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_373
timestamp -3599
transform 1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_376
timestamp -3599
transform 1 0 35696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_379
timestamp -3599
transform 1 0 35972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_385
timestamp -3599
transform 1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_388
timestamp -3599
transform 1 0 36800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_396
timestamp -3599
transform 1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_399
timestamp -3599
transform 1 0 37812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_405
timestamp -3599
transform 1 0 38364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_408
timestamp -3599
transform 1 0 38640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_411
timestamp -3599
transform 1 0 38916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_414
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_417
timestamp -3599
transform 1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_420
timestamp -3599
transform 1 0 39744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_423
timestamp -3599
transform 1 0 40020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_426
timestamp -3599
transform 1 0 40296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_429
timestamp -3599
transform 1 0 40572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_432
timestamp -3599
transform 1 0 40848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_435
timestamp -3599
transform 1 0 41124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_438
timestamp -3599
transform 1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_441
timestamp -3599
transform 1 0 41676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_444
timestamp -3599
transform 1 0 41952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp -3599
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_449
timestamp -3599
transform 1 0 42412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_452
timestamp -3599
transform 1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_455
timestamp -3599
transform 1 0 42964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_458
timestamp -3599
transform 1 0 43240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_6
timestamp -3599
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_9
timestamp -3599
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_12
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_18
timestamp -3599
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_21
timestamp -3599
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_24
timestamp -3599
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp -3599
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_35
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_38
timestamp -3599
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp -3599
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_44
timestamp -3599
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_47
timestamp -3599
transform 1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp -3599
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp -3599
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp -3599
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_59
timestamp -3599
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_62
timestamp -3599
transform 1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_65
timestamp -3599
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp -3599
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_71
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_74
timestamp -3599
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_80
timestamp -3599
transform 1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_91
timestamp -3599
transform 1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_94
timestamp -3599
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp -3599
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_100
timestamp -3599
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_103
timestamp -3599
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_106
timestamp -3599
transform 1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp -3599
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_112
timestamp -3599
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_115
timestamp -3599
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_121
timestamp -3599
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_124
timestamp -3599
transform 1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_127
timestamp -3599
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_130
timestamp -3599
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_144
timestamp -3599
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_147
timestamp -3599
transform 1 0 14628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_152
timestamp -3599
transform 1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_155
timestamp -3599
transform 1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_158
timestamp -3599
transform 1 0 15640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_161
timestamp -3599
transform 1 0 15916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_164
timestamp -3599
transform 1 0 16192 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_167
timestamp -3599
transform 1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_170
timestamp -3599
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_173
timestamp -3599
transform 1 0 17020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_176
timestamp -3599
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_179
timestamp -3599
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_182
timestamp -3599
transform 1 0 17848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_186
timestamp -3599
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_189
timestamp -3599
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_192
timestamp -3599
transform 1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -3599
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_208
timestamp -3599
transform 1 0 20240 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp -3599
transform 1 0 20516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_214
timestamp -3599
transform 1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_217
timestamp -3599
transform 1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_220
timestamp -3599
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_223
timestamp -3599
transform 1 0 21620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_226
timestamp -3599
transform 1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_229
timestamp -3599
transform 1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_232
timestamp -3599
transform 1 0 22448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_238
timestamp -3599
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_241
timestamp -3599
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_244
timestamp -3599
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_247
timestamp -3599
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp -3599
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_256
timestamp -3599
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_259
timestamp -3599
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_262
timestamp -3599
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_265
timestamp -3599
transform 1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_268
timestamp -3599
transform 1 0 25760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_271
timestamp -3599
transform 1 0 26036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_274
timestamp -3599
transform 1 0 26312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_277
timestamp -3599
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_280
timestamp -3599
transform 1 0 26864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_283
timestamp -3599
transform 1 0 27140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_286
timestamp -3599
transform 1 0 27416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_289
timestamp -3599
transform 1 0 27692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_292
timestamp -3599
transform 1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_295
timestamp -3599
transform 1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_298
timestamp -3599
transform 1 0 28520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_301
timestamp -3599
transform 1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_304
timestamp -3599
transform 1 0 29072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp -3599
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_312
timestamp -3599
transform 1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_315
timestamp -3599
transform 1 0 30084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_318
timestamp -3599
transform 1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_321
timestamp -3599
transform 1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_324
timestamp -3599
transform 1 0 30912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_327
timestamp -3599
transform 1 0 31188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_330
timestamp -3599
transform 1 0 31464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_333
timestamp -3599
transform 1 0 31740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_336
timestamp -3599
transform 1 0 32016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_339
timestamp -3599
transform 1 0 32292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_342
timestamp -3599
transform 1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_345
timestamp -3599
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_348
timestamp -3599
transform 1 0 33120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_351
timestamp -3599
transform 1 0 33396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_354
timestamp -3599
transform 1 0 33672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_357
timestamp -3599
transform 1 0 33948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_360
timestamp -3599
transform 1 0 34224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp -3599
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_365
timestamp -3599
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_368
timestamp -3599
transform 1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_371
timestamp -3599
transform 1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_374
timestamp -3599
transform 1 0 35512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_377
timestamp -3599
transform 1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_380
timestamp -3599
transform 1 0 36064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_383
timestamp -3599
transform 1 0 36340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_386
timestamp -3599
transform 1 0 36616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_389
timestamp -3599
transform 1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_392
timestamp -3599
transform 1 0 37168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_395
timestamp -3599
transform 1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_398
timestamp -3599
transform 1 0 37720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_401
timestamp -3599
transform 1 0 37996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_404
timestamp -3599
transform 1 0 38272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_407
timestamp -3599
transform 1 0 38548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_410
timestamp -3599
transform 1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_413
timestamp -3599
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_416
timestamp -3599
transform 1 0 39376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp -3599
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_421
timestamp -3599
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_424
timestamp -3599
transform 1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_427
timestamp -3599
transform 1 0 40388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_430
timestamp -3599
transform 1 0 40664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_433
timestamp -3599
transform 1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_436
timestamp -3599
transform 1 0 41216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_439
timestamp -3599
transform 1 0 41492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_442
timestamp -3599
transform 1 0 41768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_445
timestamp -3599
transform 1 0 42044 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_448
timestamp -3599
transform 1 0 42320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_451
timestamp -3599
transform 1 0 42596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_454
timestamp -3599
transform 1 0 42872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_457
timestamp -3599
transform 1 0 43148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_460
timestamp -3599
transform 1 0 43424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_463
timestamp -3599
transform 1 0 43700 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_6
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_9
timestamp -3599
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_12
timestamp -3599
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_18
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_21
timestamp -3599
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_24
timestamp -3599
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp -3599
transform 1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_30
timestamp -3599
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_33
timestamp -3599
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_36
timestamp -3599
transform 1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_39
timestamp -3599
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_42
timestamp -3599
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_45
timestamp -3599
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_48
timestamp -3599
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp -3599
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_60
timestamp -3599
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_63
timestamp -3599
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_66
timestamp -3599
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_69
timestamp -3599
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_72
timestamp -3599
transform 1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_75
timestamp -3599
transform 1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_78
timestamp -3599
transform 1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_81
timestamp -3599
transform 1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_84
timestamp -3599
transform 1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_87
timestamp -3599
transform 1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_90
timestamp -3599
transform 1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_93
timestamp -3599
transform 1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_96
timestamp -3599
transform 1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_99
timestamp -3599
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_102
timestamp -3599
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_108
timestamp -3599
transform 1 0 11040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_116
timestamp -3599
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp -3599
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_122
timestamp -3599
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_125
timestamp -3599
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_128
timestamp -3599
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_131
timestamp -3599
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_134
timestamp -3599
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_137
timestamp -3599
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_140
timestamp -3599
transform 1 0 13984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_143
timestamp -3599
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_146
timestamp -3599
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_149
timestamp -3599
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_152
timestamp -3599
transform 1 0 15088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_155
timestamp -3599
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_158
timestamp -3599
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_172
timestamp -3599
transform 1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_175
timestamp -3599
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_178
timestamp -3599
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp -3599
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp -3599
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_187
timestamp -3599
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_190
timestamp -3599
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_193
timestamp -3599
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_196
timestamp -3599
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_199
timestamp -3599
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_202
timestamp -3599
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_205
timestamp -3599
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_208
timestamp -3599
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_211
timestamp -3599
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_214
timestamp -3599
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp -3599
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp -3599
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_230
timestamp -3599
transform 1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_233
timestamp -3599
transform 1 0 22540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_236
timestamp -3599
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_239
timestamp -3599
transform 1 0 23092 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_246
timestamp -3599
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp -3599
transform 1 0 24012 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_256
timestamp -3599
transform 1 0 24656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_259
timestamp -3599
transform 1 0 24932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_262
timestamp -3599
transform 1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_265
timestamp -3599
transform 1 0 25484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_271
timestamp -3599
transform 1 0 26036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_274
timestamp -3599
transform 1 0 26312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp -3599
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_286
timestamp -3599
transform 1 0 27416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_289
timestamp -3599
transform 1 0 27692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_292
timestamp -3599
transform 1 0 27968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_295
timestamp -3599
transform 1 0 28244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_298
timestamp -3599
transform 1 0 28520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_301
timestamp -3599
transform 1 0 28796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_304
timestamp -3599
transform 1 0 29072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_307
timestamp -3599
transform 1 0 29348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_310
timestamp -3599
transform 1 0 29624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_313
timestamp -3599
transform 1 0 29900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_316
timestamp -3599
transform 1 0 30176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_319
timestamp -3599
transform 1 0 30452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_322
timestamp -3599
transform 1 0 30728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_325
timestamp -3599
transform 1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_328
timestamp -3599
transform 1 0 31280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_331
timestamp -3599
transform 1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp -3599
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_340
timestamp -3599
transform 1 0 32384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_343
timestamp -3599
transform 1 0 32660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_346
timestamp -3599
transform 1 0 32936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_349
timestamp -3599
transform 1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_352
timestamp -3599
transform 1 0 33488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_355
timestamp -3599
transform 1 0 33764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_358
timestamp -3599
transform 1 0 34040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_361
timestamp -3599
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_364
timestamp -3599
transform 1 0 34592 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_367
timestamp -3599
transform 1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_370
timestamp -3599
transform 1 0 35144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_373
timestamp -3599
transform 1 0 35420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_376
timestamp -3599
transform 1 0 35696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_379
timestamp -3599
transform 1 0 35972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_382
timestamp -3599
transform 1 0 36248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_388
timestamp -3599
transform 1 0 36800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_393
timestamp -3599
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_396
timestamp -3599
transform 1 0 37536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_399
timestamp -3599
transform 1 0 37812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_402
timestamp -3599
transform 1 0 38088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_405
timestamp -3599
transform 1 0 38364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_408
timestamp -3599
transform 1 0 38640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_411
timestamp -3599
transform 1 0 38916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_414
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_417
timestamp -3599
transform 1 0 39468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_420
timestamp -3599
transform 1 0 39744 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_423
timestamp -3599
transform 1 0 40020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_426
timestamp -3599
transform 1 0 40296 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_429
timestamp -3599
transform 1 0 40572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_432
timestamp -3599
transform 1 0 40848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_435
timestamp -3599
transform 1 0 41124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_438
timestamp -3599
transform 1 0 41400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_441
timestamp -3599
transform 1 0 41676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_444
timestamp -3599
transform 1 0 41952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp -3599
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_449
timestamp -3599
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_452
timestamp -3599
transform 1 0 42688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_455
timestamp -3599
transform 1 0 42964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_458
timestamp -3599
transform 1 0 43240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_461
timestamp -3599
transform 1 0 43516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_464
timestamp -3599
transform 1 0 43792 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_6
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp -3599
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_12
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_18
timestamp -3599
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_21
timestamp -3599
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_24
timestamp -3599
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp -3599
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_35
timestamp -3599
transform 1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp -3599
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_44
timestamp -3599
transform 1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_47
timestamp -3599
transform 1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_50
timestamp -3599
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp -3599
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_56
timestamp -3599
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_59
timestamp -3599
transform 1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_62
timestamp -3599
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp -3599
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_68
timestamp -3599
transform 1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_71
timestamp -3599
transform 1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_74
timestamp -3599
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_80
timestamp -3599
transform 1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_88
timestamp -3599
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_91
timestamp -3599
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_94
timestamp -3599
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_100
timestamp -3599
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_103
timestamp -3599
transform 1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_106
timestamp -3599
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp -3599
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_112
timestamp -3599
transform 1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_115
timestamp -3599
transform 1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_118
timestamp -3599
transform 1 0 11960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_121
timestamp -3599
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_124
timestamp -3599
transform 1 0 12512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_127
timestamp -3599
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_130
timestamp -3599
transform 1 0 13064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_133
timestamp -3599
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_136
timestamp -3599
transform 1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_144
timestamp -3599
transform 1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_147
timestamp -3599
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp -3599
transform 1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_153
timestamp -3599
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp -3599
transform 1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_159
timestamp -3599
transform 1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_162
timestamp -3599
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp -3599
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_168
timestamp -3599
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_171
timestamp -3599
transform 1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_174
timestamp -3599
transform 1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_177
timestamp -3599
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_180
timestamp -3599
transform 1 0 17664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_183
timestamp -3599
transform 1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp -3599
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp -3599
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_200
timestamp -3599
transform 1 0 19504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_206
timestamp -3599
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp -3599
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_212
timestamp -3599
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_215
timestamp -3599
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_218
timestamp -3599
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp -3599
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_224
timestamp -3599
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_227
timestamp -3599
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_230
timestamp -3599
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_233
timestamp -3599
transform 1 0 22540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_236
timestamp -3599
transform 1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_239
timestamp -3599
transform 1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_242
timestamp -3599
transform 1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_245
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_248
timestamp -3599
transform 1 0 23920 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_256
timestamp -3599
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_259
timestamp -3599
transform 1 0 24932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_262
timestamp -3599
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_265
timestamp -3599
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_268
timestamp -3599
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_271
timestamp -3599
transform 1 0 26036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_274
timestamp -3599
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_277
timestamp -3599
transform 1 0 26588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_280
timestamp -3599
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_283
timestamp -3599
transform 1 0 27140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_286
timestamp -3599
transform 1 0 27416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_289
timestamp -3599
transform 1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_292
timestamp -3599
transform 1 0 27968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_295
timestamp -3599
transform 1 0 28244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_298
timestamp -3599
transform 1 0 28520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_301
timestamp -3599
transform 1 0 28796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_304
timestamp -3599
transform 1 0 29072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_312
timestamp -3599
transform 1 0 29808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_315
timestamp -3599
transform 1 0 30084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_318
timestamp -3599
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_324
timestamp -3599
transform 1 0 30912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_327
timestamp -3599
transform 1 0 31188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_330
timestamp -3599
transform 1 0 31464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp -3599
transform 1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_336
timestamp -3599
transform 1 0 32016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_339
timestamp -3599
transform 1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_342
timestamp -3599
transform 1 0 32568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_345
timestamp -3599
transform 1 0 32844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_350
timestamp -3599
transform 1 0 33304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_353
timestamp -3599
transform 1 0 33580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_356
timestamp -3599
transform 1 0 33856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_359
timestamp -3599
transform 1 0 34132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp -3599
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_365
timestamp -3599
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_368
timestamp -3599
transform 1 0 34960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_371
timestamp -3599
transform 1 0 35236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_374
timestamp -3599
transform 1 0 35512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_377
timestamp -3599
transform 1 0 35788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_380
timestamp -3599
transform 1 0 36064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_383
timestamp -3599
transform 1 0 36340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_386
timestamp -3599
transform 1 0 36616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_389
timestamp -3599
transform 1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_392
timestamp -3599
transform 1 0 37168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_395
timestamp -3599
transform 1 0 37444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_398
timestamp -3599
transform 1 0 37720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_401
timestamp -3599
transform 1 0 37996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_404
timestamp -3599
transform 1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_407
timestamp -3599
transform 1 0 38548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_410
timestamp -3599
transform 1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_413
timestamp -3599
transform 1 0 39100 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_417
timestamp -3599
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_421
timestamp -3599
transform 1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_424
timestamp -3599
transform 1 0 40112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_427
timestamp -3599
transform 1 0 40388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_430
timestamp -3599
transform 1 0 40664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_436
timestamp -3599
transform 1 0 41216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_439
timestamp -3599
transform 1 0 41492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_442
timestamp -3599
transform 1 0 41768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_445
timestamp -3599
transform 1 0 42044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_448
timestamp -3599
transform 1 0 42320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_451
timestamp -3599
transform 1 0 42596 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_454
timestamp -3599
transform 1 0 42872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_457
timestamp -3599
transform 1 0 43148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_460
timestamp -3599
transform 1 0 43424 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_463
timestamp -3599
transform 1 0 43700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_6
timestamp -3599
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_9
timestamp -3599
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp -3599
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_18
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_21
timestamp -3599
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp -3599
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_33
timestamp -3599
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_36
timestamp -3599
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_42
timestamp -3599
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_45
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_48
timestamp -3599
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_60
timestamp -3599
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_63
timestamp -3599
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_66
timestamp -3599
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_72
timestamp -3599
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp -3599
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_84
timestamp -3599
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_87
timestamp -3599
transform 1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_90
timestamp -3599
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp -3599
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_96
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_99
timestamp -3599
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_102
timestamp -3599
transform 1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_108
timestamp -3599
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_116
timestamp -3599
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp -3599
transform 1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_122
timestamp -3599
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp -3599
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_128
timestamp -3599
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_131
timestamp -3599
transform 1 0 13156 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_134
timestamp -3599
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_137
timestamp -3599
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_140
timestamp -3599
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp -3599
transform 1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_146
timestamp -3599
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp -3599
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_152
timestamp -3599
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_155
timestamp -3599
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_158
timestamp -3599
transform 1 0 15640 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_164
timestamp -3599
transform 1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_172
timestamp -3599
transform 1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_175
timestamp -3599
transform 1 0 17204 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_178
timestamp -3599
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_181
timestamp -3599
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp -3599
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_187
timestamp -3599
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_190
timestamp -3599
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_193
timestamp -3599
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_196
timestamp -3599
transform 1 0 19136 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_199
timestamp -3599
transform 1 0 19412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_202
timestamp -3599
transform 1 0 19688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_205
timestamp -3599
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_208
timestamp -3599
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_211
timestamp -3599
transform 1 0 20516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_214
timestamp -3599
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp -3599
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_228
timestamp -3599
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_231
timestamp -3599
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_234
timestamp -3599
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_243
timestamp -3599
transform 1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_246
timestamp -3599
transform 1 0 23736 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_252
timestamp -3599
transform 1 0 24288 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_255
timestamp -3599
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_258
timestamp -3599
transform 1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_261
timestamp -3599
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_264
timestamp -3599
transform 1 0 25392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_267
timestamp -3599
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_270
timestamp -3599
transform 1 0 25944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_276
timestamp -3599
transform 1 0 26496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_284
timestamp -3599
transform 1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_287
timestamp -3599
transform 1 0 27508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_290
timestamp -3599
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_293
timestamp -3599
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_296
timestamp -3599
transform 1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_299
timestamp -3599
transform 1 0 28612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_302
timestamp -3599
transform 1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_305
timestamp -3599
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_308
timestamp -3599
transform 1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_311
timestamp -3599
transform 1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_314
timestamp -3599
transform 1 0 29992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_317
timestamp -3599
transform 1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_320
timestamp -3599
transform 1 0 30544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_323
timestamp -3599
transform 1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_329
timestamp -3599
transform 1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_332
timestamp -3599
transform 1 0 31648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp -3599
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_337
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_340
timestamp -3599
transform 1 0 32384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_343
timestamp -3599
transform 1 0 32660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_346
timestamp -3599
transform 1 0 32936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_349
timestamp -3599
transform 1 0 33212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_355
timestamp -3599
transform 1 0 33764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_358
timestamp -3599
transform 1 0 34040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_361
timestamp -3599
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_364
timestamp -3599
transform 1 0 34592 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_367
timestamp -3599
transform 1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_370
timestamp -3599
transform 1 0 35144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_373
timestamp -3599
transform 1 0 35420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_376
timestamp -3599
transform 1 0 35696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_379
timestamp -3599
transform 1 0 35972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_382
timestamp -3599
transform 1 0 36248 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_388
timestamp -3599
transform 1 0 36800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_393
timestamp -3599
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_396
timestamp -3599
transform 1 0 37536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_399
timestamp -3599
transform 1 0 37812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_402
timestamp -3599
transform 1 0 38088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_405
timestamp -3599
transform 1 0 38364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_408
timestamp -3599
transform 1 0 38640 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_411
timestamp -3599
transform 1 0 38916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_414
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_417
timestamp -3599
transform 1 0 39468 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_420
timestamp -3599
transform 1 0 39744 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_423
timestamp -3599
transform 1 0 40020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_426
timestamp -3599
transform 1 0 40296 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_429
timestamp -3599
transform 1 0 40572 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_432
timestamp -3599
transform 1 0 40848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_435
timestamp -3599
transform 1 0 41124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_438
timestamp -3599
transform 1 0 41400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_441
timestamp -3599
transform 1 0 41676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_444
timestamp -3599
transform 1 0 41952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp -3599
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_449
timestamp -3599
transform 1 0 42412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_452
timestamp -3599
transform 1 0 42688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_455
timestamp -3599
transform 1 0 42964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_458
timestamp -3599
transform 1 0 43240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_461
timestamp -3599
transform 1 0 43516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_464
timestamp -3599
transform 1 0 43792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_6
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_9
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_12
timestamp -3599
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_15
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_18
timestamp -3599
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_21
timestamp -3599
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_24
timestamp -3599
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_38
timestamp -3599
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_44
timestamp -3599
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_47
timestamp -3599
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_50
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp -3599
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp -3599
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_59
timestamp -3599
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_62
timestamp -3599
transform 1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_65
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_68
timestamp -3599
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_71
timestamp -3599
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_74
timestamp -3599
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_77
timestamp -3599
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_80
timestamp -3599
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_88
timestamp -3599
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_91
timestamp -3599
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_94
timestamp -3599
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_97
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_100
timestamp -3599
transform 1 0 10304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_103
timestamp -3599
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_106
timestamp -3599
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_109
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_112
timestamp -3599
transform 1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_115
timestamp -3599
transform 1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_118
timestamp -3599
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp -3599
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_124
timestamp -3599
transform 1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_127
timestamp -3599
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_130
timestamp -3599
transform 1 0 13064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_136
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_144
timestamp -3599
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_147
timestamp -3599
transform 1 0 14628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_155
timestamp -3599
transform 1 0 15364 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_158
timestamp -3599
transform 1 0 15640 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_161
timestamp -3599
transform 1 0 15916 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_164
timestamp -3599
transform 1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_167
timestamp -3599
transform 1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_170
timestamp -3599
transform 1 0 16744 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_173
timestamp -3599
transform 1 0 17020 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_176
timestamp -3599
transform 1 0 17296 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_179
timestamp -3599
transform 1 0 17572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_182
timestamp -3599
transform 1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_185
timestamp -3599
transform 1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_188
timestamp -3599
transform 1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp -3599
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_200
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_203
timestamp -3599
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_206
timestamp -3599
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_212
timestamp -3599
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp -3599
transform 1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_218
timestamp -3599
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_221
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_224
timestamp -3599
transform 1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_227
timestamp -3599
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_230
timestamp -3599
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_233
timestamp -3599
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_236
timestamp -3599
transform 1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_239
timestamp -3599
transform 1 0 23092 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_242
timestamp -3599
transform 1 0 23368 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_245
timestamp -3599
transform 1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_248
timestamp -3599
transform 1 0 23920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -3599
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_256
timestamp -3599
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_259
timestamp -3599
transform 1 0 24932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_268
timestamp -3599
transform 1 0 25760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_271
timestamp -3599
transform 1 0 26036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_274
timestamp -3599
transform 1 0 26312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_277
timestamp -3599
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_280
timestamp -3599
transform 1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_283
timestamp -3599
transform 1 0 27140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_286
timestamp -3599
transform 1 0 27416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_289
timestamp -3599
transform 1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_292
timestamp -3599
transform 1 0 27968 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_295
timestamp -3599
transform 1 0 28244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_298
timestamp -3599
transform 1 0 28520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_301
timestamp -3599
transform 1 0 28796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_304
timestamp -3599
transform 1 0 29072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_314
timestamp -3599
transform 1 0 29992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_323
timestamp -3599
transform 1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_326
timestamp -3599
transform 1 0 31096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_329
timestamp -3599
transform 1 0 31372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_332
timestamp -3599
transform 1 0 31648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_335
timestamp -3599
transform 1 0 31924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_338
timestamp -3599
transform 1 0 32200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_341
timestamp -3599
transform 1 0 32476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_344
timestamp -3599
transform 1 0 32752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_347
timestamp -3599
transform 1 0 33028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_350
timestamp -3599
transform 1 0 33304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_353
timestamp -3599
transform 1 0 33580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_356
timestamp -3599
transform 1 0 33856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp -3599
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_365
timestamp -3599
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_368
timestamp -3599
transform 1 0 34960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_371
timestamp -3599
transform 1 0 35236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_374
timestamp -3599
transform 1 0 35512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_377
timestamp -3599
transform 1 0 35788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_380
timestamp -3599
transform 1 0 36064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_383
timestamp -3599
transform 1 0 36340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_386
timestamp -3599
transform 1 0 36616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_389
timestamp -3599
transform 1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_392
timestamp -3599
transform 1 0 37168 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_395
timestamp -3599
transform 1 0 37444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_398
timestamp -3599
transform 1 0 37720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_401
timestamp -3599
transform 1 0 37996 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_404
timestamp -3599
transform 1 0 38272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_407
timestamp -3599
transform 1 0 38548 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_410
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_413
timestamp -3599
transform 1 0 39100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_416
timestamp -3599
transform 1 0 39376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp -3599
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_421
timestamp -3599
transform 1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_424
timestamp -3599
transform 1 0 40112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_427
timestamp -3599
transform 1 0 40388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_430
timestamp -3599
transform 1 0 40664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_433
timestamp -3599
transform 1 0 40940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_436
timestamp -3599
transform 1 0 41216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_439
timestamp -3599
transform 1 0 41492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_442
timestamp -3599
transform 1 0 41768 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_445
timestamp -3599
transform 1 0 42044 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_448
timestamp -3599
transform 1 0 42320 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_451
timestamp -3599
transform 1 0 42596 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_454
timestamp -3599
transform 1 0 42872 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_457
timestamp -3599
transform 1 0 43148 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_460
timestamp -3599
transform 1 0 43424 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_463
timestamp -3599
transform 1 0 43700 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_6
timestamp -3599
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_9
timestamp -3599
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_12
timestamp -3599
transform 1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_18
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_21
timestamp -3599
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_30
timestamp -3599
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_33
timestamp -3599
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_36
timestamp -3599
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_39
timestamp -3599
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_42
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_45
timestamp -3599
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_48
timestamp -3599
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp -3599
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_60
timestamp -3599
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_63
timestamp -3599
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_66
timestamp -3599
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp -3599
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_75
timestamp -3599
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_78
timestamp -3599
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_81
timestamp -3599
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_84
timestamp -3599
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_87
timestamp -3599
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_90
timestamp -3599
transform 1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_93
timestamp -3599
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_96
timestamp -3599
transform 1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_99
timestamp -3599
transform 1 0 10212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_102
timestamp -3599
transform 1 0 10488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_105
timestamp -3599
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_108
timestamp -3599
transform 1 0 11040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_116
timestamp -3599
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp -3599
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp -3599
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_125
timestamp -3599
transform 1 0 12604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_128
timestamp -3599
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_131
timestamp -3599
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_134
timestamp -3599
transform 1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_137
timestamp -3599
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_140
timestamp -3599
transform 1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_143
timestamp -3599
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_146
timestamp -3599
transform 1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_149
timestamp -3599
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_152
timestamp -3599
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_155
timestamp -3599
transform 1 0 15364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_158
timestamp -3599
transform 1 0 15640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_164
timestamp -3599
transform 1 0 16192 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_174
timestamp -3599
transform 1 0 17112 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_177
timestamp -3599
transform 1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_180
timestamp -3599
transform 1 0 17664 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_183
timestamp -3599
transform 1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_186
timestamp -3599
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_189
timestamp -3599
transform 1 0 18492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_192
timestamp -3599
transform 1 0 18768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_195
timestamp -3599
transform 1 0 19044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_201
timestamp -3599
transform 1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp -3599
transform 1 0 19872 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_211
timestamp -3599
transform 1 0 20516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_214
timestamp -3599
transform 1 0 20792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp -3599
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_220
timestamp -3599
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_228
timestamp -3599
transform 1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_231
timestamp -3599
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_234
timestamp -3599
transform 1 0 22632 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_240
timestamp -3599
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_243
timestamp -3599
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_246
timestamp -3599
transform 1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_249
timestamp -3599
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_252
timestamp -3599
transform 1 0 24288 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_255
timestamp -3599
transform 1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_258
timestamp -3599
transform 1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_261
timestamp -3599
transform 1 0 25116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_264
timestamp -3599
transform 1 0 25392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_267
timestamp -3599
transform 1 0 25668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_270
timestamp -3599
transform 1 0 25944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_273
timestamp -3599
transform 1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_276
timestamp -3599
transform 1 0 26496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -3599
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_281
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_287
timestamp -3599
transform 1 0 27508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_290
timestamp -3599
transform 1 0 27784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_297
timestamp -3599
transform 1 0 28428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_300
timestamp -3599
transform 1 0 28704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_303
timestamp -3599
transform 1 0 28980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_306
timestamp -3599
transform 1 0 29256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_309
timestamp -3599
transform 1 0 29532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_312
timestamp -3599
transform 1 0 29808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_315
timestamp -3599
transform 1 0 30084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_318
timestamp -3599
transform 1 0 30360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_321
timestamp -3599
transform 1 0 30636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_324
timestamp -3599
transform 1 0 30912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_327
timestamp -3599
transform 1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_330
timestamp -3599
transform 1 0 31464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp -3599
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_340
timestamp -3599
transform 1 0 32384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_343
timestamp -3599
transform 1 0 32660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_346
timestamp -3599
transform 1 0 32936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_349
timestamp -3599
transform 1 0 33212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_352
timestamp -3599
transform 1 0 33488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_355
timestamp -3599
transform 1 0 33764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_358
timestamp -3599
transform 1 0 34040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_361
timestamp -3599
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_364
timestamp -3599
transform 1 0 34592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_367
timestamp -3599
transform 1 0 34868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_372
timestamp -3599
transform 1 0 35328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_375
timestamp -3599
transform 1 0 35604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_378
timestamp -3599
transform 1 0 35880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_381
timestamp -3599
transform 1 0 36156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_384
timestamp -3599
transform 1 0 36432 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_388
timestamp -3599
transform 1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_393
timestamp -3599
transform 1 0 37260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_396
timestamp -3599
transform 1 0 37536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_399
timestamp -3599
transform 1 0 37812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_402
timestamp -3599
transform 1 0 38088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_405
timestamp -3599
transform 1 0 38364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_408
timestamp -3599
transform 1 0 38640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_411
timestamp -3599
transform 1 0 38916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_414
timestamp -3599
transform 1 0 39192 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_417
timestamp -3599
transform 1 0 39468 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_420
timestamp -3599
transform 1 0 39744 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_423
timestamp -3599
transform 1 0 40020 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_426
timestamp -3599
transform 1 0 40296 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_429
timestamp -3599
transform 1 0 40572 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_432
timestamp -3599
transform 1 0 40848 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_435
timestamp -3599
transform 1 0 41124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_438
timestamp -3599
transform 1 0 41400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_441
timestamp -3599
transform 1 0 41676 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_444
timestamp -3599
transform 1 0 41952 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp -3599
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_449
timestamp -3599
transform 1 0 42412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_452
timestamp -3599
transform 1 0 42688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_455
timestamp -3599
transform 1 0 42964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_458
timestamp -3599
transform 1 0 43240 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_6
timestamp -3599
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_9
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_12
timestamp -3599
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp -3599
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_18
timestamp -3599
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_21
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp -3599
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_35
timestamp -3599
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp -3599
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp -3599
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_47
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_50
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp -3599
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_56
timestamp -3599
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_59
timestamp -3599
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_68
timestamp -3599
transform 1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_71
timestamp -3599
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_74
timestamp -3599
transform 1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_77
timestamp -3599
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_80
timestamp -3599
transform 1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_88
timestamp -3599
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_91
timestamp -3599
transform 1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_94
timestamp -3599
transform 1 0 9752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp -3599
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_100
timestamp -3599
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_103
timestamp -3599
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_106
timestamp -3599
transform 1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_109
timestamp -3599
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_112
timestamp -3599
transform 1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_115
timestamp -3599
transform 1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_118
timestamp -3599
transform 1 0 11960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_121
timestamp -3599
transform 1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp -3599
transform 1 0 12972 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_136
timestamp -3599
transform 1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_144
timestamp -3599
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_147
timestamp -3599
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp -3599
transform 1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp -3599
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_159
timestamp -3599
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_162
timestamp -3599
transform 1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp -3599
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp -3599
transform 1 0 16560 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_171
timestamp -3599
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_174
timestamp -3599
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_180
timestamp -3599
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_183
timestamp -3599
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_186
timestamp -3599
transform 1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_192
timestamp -3599
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_200
timestamp -3599
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_203
timestamp -3599
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_206
timestamp -3599
transform 1 0 20056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_210
timestamp -3599
transform 1 0 20424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_213
timestamp -3599
transform 1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_216
timestamp -3599
transform 1 0 20976 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_219
timestamp -3599
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_222
timestamp -3599
transform 1 0 21528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_225
timestamp -3599
transform 1 0 21804 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_228
timestamp -3599
transform 1 0 22080 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_231
timestamp -3599
transform 1 0 22356 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_235
timestamp -3599
transform 1 0 22724 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_238
timestamp -3599
transform 1 0 23000 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_241
timestamp -3599
transform 1 0 23276 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_244
timestamp -3599
transform 1 0 23552 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_247
timestamp -3599
transform 1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp -3599
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_256
timestamp -3599
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_259
timestamp -3599
transform 1 0 24932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_265
timestamp -3599
transform 1 0 25484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_268
timestamp -3599
transform 1 0 25760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_271
timestamp -3599
transform 1 0 26036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_274
timestamp -3599
transform 1 0 26312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_277
timestamp -3599
transform 1 0 26588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_280
timestamp -3599
transform 1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_283
timestamp -3599
transform 1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_286
timestamp -3599
transform 1 0 27416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_289
timestamp -3599
transform 1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_292
timestamp -3599
transform 1 0 27968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_295
timestamp -3599
transform 1 0 28244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_298
timestamp -3599
transform 1 0 28520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_301
timestamp -3599
transform 1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_304
timestamp -3599
transform 1 0 29072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_312
timestamp -3599
transform 1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_315
timestamp -3599
transform 1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_318
timestamp -3599
transform 1 0 30360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_321
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_324
timestamp -3599
transform 1 0 30912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_327
timestamp -3599
transform 1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_330
timestamp -3599
transform 1 0 31464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_333
timestamp -3599
transform 1 0 31740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_336
timestamp -3599
transform 1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_339
timestamp -3599
transform 1 0 32292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_342
timestamp -3599
transform 1 0 32568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_345
timestamp -3599
transform 1 0 32844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_348
timestamp -3599
transform 1 0 33120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_351
timestamp -3599
transform 1 0 33396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_354
timestamp -3599
transform 1 0 33672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_357
timestamp -3599
transform 1 0 33948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_360
timestamp -3599
transform 1 0 34224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp -3599
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_365
timestamp -3599
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_368
timestamp -3599
transform 1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_371
timestamp -3599
transform 1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_374
timestamp -3599
transform 1 0 35512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_377
timestamp -3599
transform 1 0 35788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_380
timestamp -3599
transform 1 0 36064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_383
timestamp -3599
transform 1 0 36340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_386
timestamp -3599
transform 1 0 36616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_389
timestamp -3599
transform 1 0 36892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_392
timestamp -3599
transform 1 0 37168 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_395
timestamp -3599
transform 1 0 37444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_399
timestamp -3599
transform 1 0 37812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_402
timestamp -3599
transform 1 0 38088 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_405
timestamp -3599
transform 1 0 38364 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_408
timestamp -3599
transform 1 0 38640 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_411
timestamp -3599
transform 1 0 38916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_414
timestamp -3599
transform 1 0 39192 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_417
timestamp -3599
transform 1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_421
timestamp -3599
transform 1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_424
timestamp -3599
transform 1 0 40112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_427
timestamp -3599
transform 1 0 40388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_430
timestamp -3599
transform 1 0 40664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_436
timestamp -3599
transform 1 0 41216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_439
timestamp -3599
transform 1 0 41492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_442
timestamp -3599
transform 1 0 41768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_445
timestamp -3599
transform 1 0 42044 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_448
timestamp -3599
transform 1 0 42320 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7
timestamp -3599
transform 1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_10
timestamp -3599
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_13
timestamp -3599
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_16
timestamp -3599
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_19
timestamp -3599
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_22
timestamp -3599
transform 1 0 3128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_25
timestamp -3599
transform 1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_28
timestamp -3599
transform 1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_31
timestamp -3599
transform 1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_34
timestamp -3599
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_37
timestamp -3599
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_40
timestamp -3599
transform 1 0 4784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_43
timestamp -3599
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_46
timestamp -3599
transform 1 0 5336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_49
timestamp -3599
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_52
timestamp -3599
transform 1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_60
timestamp -3599
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_63
timestamp -3599
transform 1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_66
timestamp -3599
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_72
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_75
timestamp -3599
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_78
timestamp -3599
transform 1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp -3599
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_84
timestamp -3599
transform 1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_87
timestamp -3599
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_93
timestamp -3599
transform 1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_96
timestamp -3599
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_99
timestamp -3599
transform 1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_102
timestamp -3599
transform 1 0 10488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_108
timestamp -3599
transform 1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_116
timestamp -3599
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp -3599
transform 1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_122
timestamp -3599
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_126
timestamp -3599
transform 1 0 12696 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_129
timestamp -3599
transform 1 0 12972 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_132
timestamp -3599
transform 1 0 13248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_135
timestamp -3599
transform 1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_138
timestamp -3599
transform 1 0 13800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_141
timestamp -3599
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_144
timestamp -3599
transform 1 0 14352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_149
timestamp -3599
transform 1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_157
timestamp -3599
transform 1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_160
timestamp -3599
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_163
timestamp -3599
transform 1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp -3599
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_172
timestamp -3599
transform 1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_175
timestamp -3599
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_178
timestamp -3599
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_181
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_184
timestamp -3599
transform 1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_187
timestamp -3599
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_190
timestamp -3599
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp -3599
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_196
timestamp -3599
transform 1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_199
timestamp -3599
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_202
timestamp -3599
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_205
timestamp -3599
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_208
timestamp -3599
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_211
timestamp -3599
transform 1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_214
timestamp -3599
transform 1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_217
timestamp -3599
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_228
timestamp -3599
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_231
timestamp -3599
transform 1 0 22356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_234
timestamp -3599
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_237
timestamp -3599
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_240
timestamp -3599
transform 1 0 23184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_243
timestamp -3599
transform 1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_246
timestamp -3599
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_249
timestamp -3599
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_252
timestamp -3599
transform 1 0 24288 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_255
timestamp -3599
transform 1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_258
timestamp -3599
transform 1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_261
timestamp -3599
transform 1 0 25116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_264
timestamp -3599
transform 1 0 25392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_267
timestamp -3599
transform 1 0 25668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_270
timestamp -3599
transform 1 0 25944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_273
timestamp -3599
transform 1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_276
timestamp -3599
transform 1 0 26496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -3599
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_284
timestamp -3599
transform 1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_287
timestamp -3599
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_290
timestamp -3599
transform 1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_293
timestamp -3599
transform 1 0 28060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_298
timestamp -3599
transform 1 0 28520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_301
timestamp -3599
transform 1 0 28796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_304
timestamp -3599
transform 1 0 29072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_307
timestamp -3599
transform 1 0 29348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_310
timestamp -3599
transform 1 0 29624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_313
timestamp -3599
transform 1 0 29900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_316
timestamp -3599
transform 1 0 30176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_319
timestamp -3599
transform 1 0 30452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_322
timestamp -3599
transform 1 0 30728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_325
timestamp -3599
transform 1 0 31004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_328
timestamp -3599
transform 1 0 31280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_331
timestamp -3599
transform 1 0 31556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp -3599
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_340
timestamp -3599
transform 1 0 32384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_343
timestamp -3599
transform 1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_346
timestamp -3599
transform 1 0 32936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_349
timestamp -3599
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_352
timestamp -3599
transform 1 0 33488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_355
timestamp -3599
transform 1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_358
timestamp -3599
transform 1 0 34040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_364
timestamp -3599
transform 1 0 34592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_367
timestamp -3599
transform 1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_370
timestamp -3599
transform 1 0 35144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_373
timestamp -3599
transform 1 0 35420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_376
timestamp -3599
transform 1 0 35696 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_379
timestamp -3599
transform 1 0 35972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_387
timestamp -3599
transform 1 0 36708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp -3599
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_396
timestamp -3599
transform 1 0 37536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_399
timestamp -3599
transform 1 0 37812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_402
timestamp -3599
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_405
timestamp -3599
transform 1 0 38364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_408
timestamp -3599
transform 1 0 38640 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_411
timestamp -3599
transform 1 0 38916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_414
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_417
timestamp -3599
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_420
timestamp -3599
transform 1 0 39744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_423
timestamp -3599
transform 1 0 40020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_426
timestamp -3599
transform 1 0 40296 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_429
timestamp -3599
transform 1 0 40572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_432
timestamp -3599
transform 1 0 40848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_437
timestamp -3599
transform 1 0 41308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_440
timestamp -3599
transform 1 0 41584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_449
timestamp -3599
transform 1 0 42412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_18
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_24
timestamp -3599
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_34
timestamp -3599
transform 1 0 4232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_37
timestamp -3599
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp -3599
transform 1 0 4784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_46
timestamp -3599
transform 1 0 5336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_49
timestamp -3599
transform 1 0 5612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_52
timestamp -3599
transform 1 0 5888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_55
timestamp -3599
transform 1 0 6164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_62
timestamp -3599
transform 1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_65
timestamp -3599
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_68
timestamp -3599
transform 1 0 7360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_71
timestamp -3599
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_74
timestamp -3599
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_77
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_80
timestamp -3599
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_90
timestamp -3599
transform 1 0 9384 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_96
timestamp -3599
transform 1 0 9936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_102
timestamp -3599
transform 1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_110
timestamp -3599
transform 1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_113
timestamp -3599
transform 1 0 11500 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_125
timestamp -3599
transform 1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_128
timestamp -3599
transform 1 0 12880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_131
timestamp -3599
transform 1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_134
timestamp -3599
transform 1 0 13432 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp -3599
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_146
timestamp -3599
transform 1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_149
timestamp -3599
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_152
timestamp -3599
transform 1 0 15088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_155
timestamp -3599
transform 1 0 15364 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp -3599
transform 1 0 15640 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_162
timestamp -3599
transform 1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_168
timestamp -3599
transform 1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_176
timestamp -3599
transform 1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_179
timestamp -3599
transform 1 0 17572 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_185
timestamp -3599
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_188
timestamp -3599
transform 1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_191
timestamp -3599
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp -3599
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_202
timestamp -3599
transform 1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_205
timestamp -3599
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_208
timestamp -3599
transform 1 0 20240 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp -3599
transform 1 0 20516 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_214
timestamp -3599
transform 1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_217
timestamp -3599
transform 1 0 21068 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_220
timestamp -3599
transform 1 0 21344 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_227
timestamp -3599
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp -3599
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_233
timestamp -3599
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_236
timestamp -3599
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_239
timestamp -3599
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_242
timestamp -3599
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_248
timestamp -3599
transform 1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_256
timestamp -3599
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_259
timestamp -3599
transform 1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp -3599
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_269
timestamp -3599
transform 1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_272
timestamp -3599
transform 1 0 26128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_275
timestamp -3599
transform 1 0 26404 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_284
timestamp -3599
transform 1 0 27232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_287
timestamp -3599
transform 1 0 27508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_291
timestamp -3599
transform 1 0 27876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_294
timestamp -3599
transform 1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_300
timestamp -3599
transform 1 0 28704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_303
timestamp -3599
transform 1 0 28980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp -3599
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_312
timestamp -3599
transform 1 0 29808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_316
timestamp -3599
transform 1 0 30176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_319
timestamp -3599
transform 1 0 30452 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_322
timestamp -3599
transform 1 0 30728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_325
timestamp -3599
transform 1 0 31004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_328
timestamp -3599
transform 1 0 31280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_331
timestamp -3599
transform 1 0 31556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_334
timestamp -3599
transform 1 0 31832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_337
timestamp -3599
transform 1 0 32108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_340
timestamp -3599
transform 1 0 32384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_343
timestamp -3599
transform 1 0 32660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_346
timestamp -3599
transform 1 0 32936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_349
timestamp -3599
transform 1 0 33212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_352
timestamp -3599
transform 1 0 33488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_355
timestamp -3599
transform 1 0 33764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_358
timestamp -3599
transform 1 0 34040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp -3599
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_365
timestamp -3599
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_368
timestamp -3599
transform 1 0 34960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_371
timestamp -3599
transform 1 0 35236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_374
timestamp -3599
transform 1 0 35512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_377
timestamp -3599
transform 1 0 35788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_382
timestamp -3599
transform 1 0 36248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_385
timestamp -3599
transform 1 0 36524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_388
timestamp -3599
transform 1 0 36800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_391
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_394
timestamp -3599
transform 1 0 37352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_397
timestamp -3599
transform 1 0 37628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_400
timestamp -3599
transform 1 0 37904 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_404
timestamp -3599
transform 1 0 38272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_407
timestamp -3599
transform 1 0 38548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_410
timestamp -3599
transform 1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_413
timestamp -3599
transform 1 0 39100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_416
timestamp -3599
transform 1 0 39376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp -3599
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_424
timestamp -3599
transform 1 0 40112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_427
timestamp -3599
transform 1 0 40388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_432
timestamp -3599
transform 1 0 40848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_438
timestamp -3599
transform 1 0 41400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_441
timestamp -3599
transform 1 0 41676 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_470
timestamp -3599
transform 1 0 44344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp -3599
transform 1 0 18952 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_201
timestamp -3599
transform 1 0 19596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_204
timestamp -3599
transform 1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_207
timestamp -3599
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_210
timestamp -3599
transform 1 0 20424 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_213
timestamp -3599
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_216
timestamp -3599
transform 1 0 20976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_219
timestamp -3599
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_228
timestamp -3599
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_231
timestamp -3599
transform 1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_234
timestamp -3599
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_237
timestamp -3599
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_240
timestamp -3599
transform 1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_243
timestamp -3599
transform 1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_246
timestamp -3599
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_249
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_253
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_256
timestamp -3599
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_259
timestamp -3599
transform 1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_262
timestamp -3599
transform 1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_265
timestamp -3599
transform 1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_268
timestamp -3599
transform 1 0 25760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_271
timestamp -3599
transform 1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_274
timestamp -3599
transform 1 0 26312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp -3599
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_284
timestamp -3599
transform 1 0 27232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_287
timestamp -3599
transform 1 0 27508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_290
timestamp -3599
transform 1 0 27784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_293
timestamp -3599
transform 1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_296
timestamp -3599
transform 1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_299
timestamp -3599
transform 1 0 28612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_302
timestamp -3599
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp -3599
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_309
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_312
timestamp -3599
transform 1 0 29808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_315
timestamp -3599
transform 1 0 30084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_318
timestamp -3599
transform 1 0 30360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_321
timestamp -3599
transform 1 0 30636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_324
timestamp -3599
transform 1 0 30912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_327
timestamp -3599
transform 1 0 31188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_330
timestamp -3599
transform 1 0 31464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp -3599
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_340
timestamp -3599
transform 1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_343
timestamp -3599
transform 1 0 32660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_346
timestamp -3599
transform 1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_349
timestamp -3599
transform 1 0 33212 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_352
timestamp -3599
transform 1 0 33488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_355
timestamp -3599
transform 1 0 33764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_358
timestamp -3599
transform 1 0 34040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_361
timestamp -3599
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_365
timestamp -3599
transform 1 0 34684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_368
timestamp -3599
transform 1 0 34960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_371
timestamp -3599
transform 1 0 35236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_374
timestamp -3599
transform 1 0 35512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_377
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_380
timestamp -3599
transform 1 0 36064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_383
timestamp -3599
transform 1 0 36340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_386
timestamp -3599
transform 1 0 36616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_393
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_396
timestamp -3599
transform 1 0 37536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_399
timestamp -3599
transform 1 0 37812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_402
timestamp -3599
transform 1 0 38088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_405
timestamp -3599
transform 1 0 38364 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_409
timestamp -3599
transform 1 0 38732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_418
timestamp -3599
transform 1 0 39560 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp -3599
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 43884 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 44252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 43884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 43884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 44252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 43884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 43516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 44252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 42780 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 43148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 43884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 44252 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 44252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 43608 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 43240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 42872 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 43516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 43884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 43148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 42504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 42780 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 43884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 44252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 43884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 43884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 44252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform 1 0 38824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform 1 0 43148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform 1 0 43516 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform 1 0 43884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform 1 0 44252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 43976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 43884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 42136 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 41768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 44252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 43516 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform 1 0 39192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 39836 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 40204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 40572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 40940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform 1 0 41308 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform 1 0 41676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform 1 0 42412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform 1 0 42780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform -1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform -1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform -1 0 1840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform -1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform -1 0 2576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform -1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform -1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform -1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform -1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform -1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform -1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform -1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform -1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform -1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform -1 0 9384 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform -1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 18584 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform -1 0 18952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform -1 0 19596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform 1 0 14168 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform 1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform 1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 16744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 38732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 44896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 44896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 44896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 44896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp -3599
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp -3599
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_46
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_47
timestamp -3599
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_54
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_55
timestamp -3599
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_59
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_62
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_63
timestamp -3599
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_67
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp -3599
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_73
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_77
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp -3599
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_82
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_86
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_87
timestamp -3599
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_89
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_90
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_91
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_92
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_93
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_94
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_95
timestamp -3599
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_96
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_97
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_98
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_103
timestamp -3599
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_106
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_107
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_108
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_109
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_110
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_111
timestamp -3599
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_112
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_114
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_115
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_116
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_118
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_119
timestamp -3599
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_122
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_123
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_124
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_125
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_127
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_128
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_129
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_130
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_131
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp -3599
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp -3599
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1096 120 1216 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 45880 1096 46000 1216 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 45880 3816 46000 3936 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 45880 4088 46000 4208 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 45880 4360 46000 4480 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 45880 4632 46000 4752 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 45880 4904 46000 5024 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 45880 5176 46000 5296 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 45880 5448 46000 5568 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 45880 5720 46000 5840 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 45880 5992 46000 6112 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 45880 6264 46000 6384 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 45880 1368 46000 1488 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 45880 6536 46000 6656 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 45880 6808 46000 6928 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 45880 7080 46000 7200 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 45880 7352 46000 7472 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 45880 7624 46000 7744 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 45880 7896 46000 8016 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 45880 8168 46000 8288 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 45880 8440 46000 8560 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 45880 8712 46000 8832 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 45880 8984 46000 9104 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 45880 1640 46000 1760 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 45880 9256 46000 9376 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 45880 9528 46000 9648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 45880 1912 46000 2032 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 45880 2184 46000 2304 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 45880 2456 46000 2576 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 45880 2728 46000 2848 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 45880 3000 46000 3120 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 45880 3272 46000 3392 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 45880 3544 46000 3664 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 3882 0 3938 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 25042 0 25098 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 27158 0 27214 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 29274 0 29330 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 31390 0 31446 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 33506 0 33562 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 35622 0 35678 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 37738 0 37794 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 39854 0 39910 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 41970 0 42026 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 44086 0 44142 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 5998 0 6054 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 8114 0 8170 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 10230 0 10286 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 12346 0 12402 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 14462 0 14518 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 16578 0 16634 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 18694 0 18750 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 20810 0 20866 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 22926 0 22982 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 38750 11096 38806 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 42430 11096 42486 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 42798 11096 42854 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 43166 11096 43222 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 43534 11096 43590 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 43902 11096 43958 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 44270 11096 44326 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 44638 11096 44694 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 45006 11096 45062 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 45374 11096 45430 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 45742 11096 45798 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 39118 11096 39174 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 39486 11096 39542 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 39854 11096 39910 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 40222 11096 40278 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 40590 11096 40646 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 40958 11096 41014 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 41326 11096 41382 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 41694 11096 41750 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 42062 11096 42118 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 110 11096 166 11152 0 FreeSans 224 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 478 11096 534 11152 0 FreeSans 224 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 846 11096 902 11152 0 FreeSans 224 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 1214 11096 1270 11152 0 FreeSans 224 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 1582 11096 1638 11152 0 FreeSans 224 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 1950 11096 2006 11152 0 FreeSans 224 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 2318 11096 2374 11152 0 FreeSans 224 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 2686 11096 2742 11152 0 FreeSans 224 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 3054 11096 3110 11152 0 FreeSans 224 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 3422 11096 3478 11152 0 FreeSans 224 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 3790 11096 3846 11152 0 FreeSans 224 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 4158 11096 4214 11152 0 FreeSans 224 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 4526 11096 4582 11152 0 FreeSans 224 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 4894 11096 4950 11152 0 FreeSans 224 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 5262 11096 5318 11152 0 FreeSans 224 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 5630 11096 5686 11152 0 FreeSans 224 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 5998 11096 6054 11152 0 FreeSans 224 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 6366 11096 6422 11152 0 FreeSans 224 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 6734 11096 6790 11152 0 FreeSans 224 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 7102 11096 7158 11152 0 FreeSans 224 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 7470 11096 7526 11152 0 FreeSans 224 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 11150 11096 11206 11152 0 FreeSans 224 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 11518 11096 11574 11152 0 FreeSans 224 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 11886 11096 11942 11152 0 FreeSans 224 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 12254 11096 12310 11152 0 FreeSans 224 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 12622 11096 12678 11152 0 FreeSans 224 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 12990 11096 13046 11152 0 FreeSans 224 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 7838 11096 7894 11152 0 FreeSans 224 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 8206 11096 8262 11152 0 FreeSans 224 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 8574 11096 8630 11152 0 FreeSans 224 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 8942 11096 8998 11152 0 FreeSans 224 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 9310 11096 9366 11152 0 FreeSans 224 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 9678 11096 9734 11152 0 FreeSans 224 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 10046 11096 10102 11152 0 FreeSans 224 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 10414 11096 10470 11152 0 FreeSans 224 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 10782 11096 10838 11152 0 FreeSans 224 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 13358 11096 13414 11152 0 FreeSans 224 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal2 s 17038 11096 17094 11152 0 FreeSans 224 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal2 s 17406 11096 17462 11152 0 FreeSans 224 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal2 s 17774 11096 17830 11152 0 FreeSans 224 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal2 s 18142 11096 18198 11152 0 FreeSans 224 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal2 s 18510 11096 18566 11152 0 FreeSans 224 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal2 s 18878 11096 18934 11152 0 FreeSans 224 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal2 s 13726 11096 13782 11152 0 FreeSans 224 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal2 s 14094 11096 14150 11152 0 FreeSans 224 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal2 s 14462 11096 14518 11152 0 FreeSans 224 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal2 s 14830 11096 14886 11152 0 FreeSans 224 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal2 s 15198 11096 15254 11152 0 FreeSans 224 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal2 s 15566 11096 15622 11152 0 FreeSans 224 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal2 s 15934 11096 15990 11152 0 FreeSans 224 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal2 s 16302 11096 16358 11152 0 FreeSans 224 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal2 s 16670 11096 16726 11152 0 FreeSans 224 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal2 s 19246 11096 19302 11152 0 FreeSans 224 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal2 s 19614 11096 19670 11152 0 FreeSans 224 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal2 s 19982 11096 20038 11152 0 FreeSans 224 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal2 s 20350 11096 20406 11152 0 FreeSans 224 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal2 s 23662 11096 23718 11152 0 FreeSans 224 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal2 s 24030 11096 24086 11152 0 FreeSans 224 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal2 s 24398 11096 24454 11152 0 FreeSans 224 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal2 s 24766 11096 24822 11152 0 FreeSans 224 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal2 s 25134 11096 25190 11152 0 FreeSans 224 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal2 s 25502 11096 25558 11152 0 FreeSans 224 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal2 s 25870 11096 25926 11152 0 FreeSans 224 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal2 s 26238 11096 26294 11152 0 FreeSans 224 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal2 s 20718 11096 20774 11152 0 FreeSans 224 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal2 s 21086 11096 21142 11152 0 FreeSans 224 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal2 s 21454 11096 21510 11152 0 FreeSans 224 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal2 s 21822 11096 21878 11152 0 FreeSans 224 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal2 s 22190 11096 22246 11152 0 FreeSans 224 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal2 s 22558 11096 22614 11152 0 FreeSans 224 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal2 s 22926 11096 22982 11152 0 FreeSans 224 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal2 s 23294 11096 23350 11152 0 FreeSans 224 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal2 s 26606 11096 26662 11152 0 FreeSans 224 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal2 s 30286 11096 30342 11152 0 FreeSans 224 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal2 s 30654 11096 30710 11152 0 FreeSans 224 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal2 s 31022 11096 31078 11152 0 FreeSans 224 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal2 s 31390 11096 31446 11152 0 FreeSans 224 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal2 s 31758 11096 31814 11152 0 FreeSans 224 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal2 s 32126 11096 32182 11152 0 FreeSans 224 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal2 s 26974 11096 27030 11152 0 FreeSans 224 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal2 s 27342 11096 27398 11152 0 FreeSans 224 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal2 s 27710 11096 27766 11152 0 FreeSans 224 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal2 s 28078 11096 28134 11152 0 FreeSans 224 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal2 s 28446 11096 28502 11152 0 FreeSans 224 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal2 s 28814 11096 28870 11152 0 FreeSans 224 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal2 s 29182 11096 29238 11152 0 FreeSans 224 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal2 s 29550 11096 29606 11152 0 FreeSans 224 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal2 s 29918 11096 29974 11152 0 FreeSans 224 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal2 s 32494 11096 32550 11152 0 FreeSans 224 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal2 s 36174 11096 36230 11152 0 FreeSans 224 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal2 s 36542 11096 36598 11152 0 FreeSans 224 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal2 s 36910 11096 36966 11152 0 FreeSans 224 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal2 s 37278 11096 37334 11152 0 FreeSans 224 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal2 s 37646 11096 37702 11152 0 FreeSans 224 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal2 s 38014 11096 38070 11152 0 FreeSans 224 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal2 s 32862 11096 32918 11152 0 FreeSans 224 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal2 s 33230 11096 33286 11152 0 FreeSans 224 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal2 s 33598 11096 33654 11152 0 FreeSans 224 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal2 s 33966 11096 34022 11152 0 FreeSans 224 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal2 s 34334 11096 34390 11152 0 FreeSans 224 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal2 s 34702 11096 34758 11152 0 FreeSans 224 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal2 s 35070 11096 35126 11152 0 FreeSans 224 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal2 s 35438 11096 35494 11152 0 FreeSans 224 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal2 s 35806 11096 35862 11152 0 FreeSans 224 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal2 s 1766 0 1822 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 38382 11096 38438 11152 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3004 0 3324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 11092 3324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 11092 9324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 11092 15324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 11092 21324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 11092 27324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 11092 33324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 11092 39324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 11092 2264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 11092 8264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 11092 14264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 11092 20264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 11092 26264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 11092 32264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 11092 38264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 0 44264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 0 44264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 11092 44264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 23000 8704 23000 8704 0 VGND
rlabel metal1 23000 8160 23000 8160 0 VPWR
rlabel metal3 758 1156 758 1156 0 FrameData[0]
rlabel metal3 919 3876 919 3876 0 FrameData[10]
rlabel metal2 7498 3808 7498 3808 0 FrameData[11]
rlabel metal3 19596 4080 19596 4080 0 FrameData[12]
rlabel metal2 21574 7361 21574 7361 0 FrameData[13]
rlabel metal3 919 4964 919 4964 0 FrameData[14]
rlabel metal1 19274 7888 19274 7888 0 FrameData[15]
rlabel metal1 19642 6358 19642 6358 0 FrameData[16]
rlabel metal1 25898 6290 25898 6290 0 FrameData[17]
rlabel metal3 919 6052 919 6052 0 FrameData[18]
rlabel metal1 15548 2278 15548 2278 0 FrameData[19]
rlabel metal2 15778 2125 15778 2125 0 FrameData[1]
rlabel metal1 19918 3026 19918 3026 0 FrameData[20]
rlabel metal1 10212 3094 10212 3094 0 FrameData[21]
rlabel metal3 574 7140 574 7140 0 FrameData[22]
rlabel metal1 21436 3026 21436 3026 0 FrameData[23]
rlabel metal3 620 7684 620 7684 0 FrameData[24]
rlabel metal3 712 7956 712 7956 0 FrameData[25]
rlabel metal3 942 8228 942 8228 0 FrameData[26]
rlabel metal2 30130 7089 30130 7089 0 FrameData[27]
rlabel metal3 1356 8772 1356 8772 0 FrameData[28]
rlabel metal2 4002 8415 4002 8415 0 FrameData[29]
rlabel metal2 19550 2533 19550 2533 0 FrameData[2]
rlabel metal2 26542 8619 26542 8619 0 FrameData[30]
rlabel metal2 41906 8517 41906 8517 0 FrameData[31]
rlabel metal1 21160 3910 21160 3910 0 FrameData[3]
rlabel metal3 1471 2244 1471 2244 0 FrameData[4]
rlabel metal3 13914 2516 13914 2516 0 FrameData[5]
rlabel metal3 919 2788 919 2788 0 FrameData[6]
rlabel metal3 21988 3128 21988 3128 0 FrameData[7]
rlabel metal2 12466 2567 12466 2567 0 FrameData[8]
rlabel metal2 19642 4318 19642 4318 0 FrameData[9]
rlabel metal3 45150 1156 45150 1156 0 FrameData_O[0]
rlabel metal3 45449 3876 45449 3876 0 FrameData_O[10]
rlabel metal3 45196 4148 45196 4148 0 FrameData_O[11]
rlabel metal3 45012 4420 45012 4420 0 FrameData_O[12]
rlabel metal3 45196 4692 45196 4692 0 FrameData_O[13]
rlabel metal3 45449 4964 45449 4964 0 FrameData_O[14]
rlabel metal3 45196 5236 45196 5236 0 FrameData_O[15]
rlabel metal3 45150 5508 45150 5508 0 FrameData_O[16]
rlabel metal3 44828 5780 44828 5780 0 FrameData_O[17]
rlabel metal2 44482 5967 44482 5967 0 FrameData_O[18]
rlabel metal3 44460 6324 44460 6324 0 FrameData_O[19]
rlabel metal3 44644 1428 44644 1428 0 FrameData_O[1]
rlabel metal3 44644 6596 44644 6596 0 FrameData_O[20]
rlabel metal2 44114 6647 44114 6647 0 FrameData_O[21]
rlabel metal2 44482 6885 44482 6885 0 FrameData_O[22]
rlabel metal3 45196 7412 45196 7412 0 FrameData_O[23]
rlabel metal3 45380 7684 45380 7684 0 FrameData_O[24]
rlabel metal3 44736 7956 44736 7956 0 FrameData_O[25]
rlabel metal1 43470 7990 43470 7990 0 FrameData_O[26]
rlabel metal1 43792 7514 43792 7514 0 FrameData_O[27]
rlabel metal1 44114 6664 44114 6664 0 FrameData_O[28]
rlabel metal2 43378 8279 43378 8279 0 FrameData_O[29]
rlabel metal3 44460 1700 44460 1700 0 FrameData_O[2]
rlabel metal2 42734 8687 42734 8687 0 FrameData_O[30]
rlabel metal2 43010 8551 43010 8551 0 FrameData_O[31]
rlabel metal3 45380 1972 45380 1972 0 FrameData_O[3]
rlabel metal3 45012 2244 45012 2244 0 FrameData_O[4]
rlabel metal3 45196 2516 45196 2516 0 FrameData_O[5]
rlabel metal3 45449 2788 45449 2788 0 FrameData_O[6]
rlabel metal3 45196 3060 45196 3060 0 FrameData_O[7]
rlabel metal3 45012 3332 45012 3332 0 FrameData_O[8]
rlabel metal3 45196 3604 45196 3604 0 FrameData_O[9]
rlabel metal2 3910 106 3910 106 0 FrameStrobe[0]
rlabel metal1 25806 3094 25806 3094 0 FrameStrobe[10]
rlabel metal2 27186 55 27186 55 0 FrameStrobe[11]
rlabel metal1 29992 3026 29992 3026 0 FrameStrobe[12]
rlabel metal2 31418 140 31418 140 0 FrameStrobe[13]
rlabel metal2 33534 1401 33534 1401 0 FrameStrobe[14]
rlabel metal2 35650 667 35650 667 0 FrameStrobe[15]
rlabel metal1 37674 6766 37674 6766 0 FrameStrobe[16]
rlabel metal1 40480 7378 40480 7378 0 FrameStrobe[17]
rlabel metal1 42274 7310 42274 7310 0 FrameStrobe[18]
rlabel metal2 44114 55 44114 55 0 FrameStrobe[19]
rlabel metal2 6026 106 6026 106 0 FrameStrobe[1]
rlabel metal2 8142 55 8142 55 0 FrameStrobe[2]
rlabel metal1 10074 3026 10074 3026 0 FrameStrobe[3]
rlabel metal2 12374 1534 12374 1534 0 FrameStrobe[4]
rlabel metal2 14490 1534 14490 1534 0 FrameStrobe[5]
rlabel metal2 16606 1500 16606 1500 0 FrameStrobe[6]
rlabel metal2 18722 1738 18722 1738 0 FrameStrobe[7]
rlabel metal2 20838 1772 20838 1772 0 FrameStrobe[8]
rlabel metal2 22954 55 22954 55 0 FrameStrobe[9]
rlabel metal2 38916 8602 38916 8602 0 FrameStrobe_O[0]
rlabel metal1 43378 8364 43378 8364 0 FrameStrobe_O[10]
rlabel metal1 43516 8602 43516 8602 0 FrameStrobe_O[11]
rlabel metal1 43792 8330 43792 8330 0 FrameStrobe_O[12]
rlabel metal1 44482 8568 44482 8568 0 FrameStrobe_O[13]
rlabel metal1 43976 8058 43976 8058 0 FrameStrobe_O[14]
rlabel metal1 44252 7514 44252 7514 0 FrameStrobe_O[15]
rlabel metal2 42366 8160 42366 8160 0 FrameStrobe_O[16]
rlabel metal1 42044 7718 42044 7718 0 FrameStrobe_O[17]
rlabel metal1 44942 6426 44942 6426 0 FrameStrobe_O[18]
rlabel metal1 43838 6902 43838 6902 0 FrameStrobe_O[19]
rlabel metal2 39422 9863 39422 9863 0 FrameStrobe_O[1]
rlabel metal1 39790 8602 39790 8602 0 FrameStrobe_O[2]
rlabel metal1 40158 8330 40158 8330 0 FrameStrobe_O[3]
rlabel metal1 40526 8602 40526 8602 0 FrameStrobe_O[4]
rlabel metal1 41032 8602 41032 8602 0 FrameStrobe_O[5]
rlabel metal2 40986 11097 40986 11097 0 FrameStrobe_O[6]
rlabel metal2 41354 9720 41354 9720 0 FrameStrobe_O[7]
rlabel metal1 42182 8602 42182 8602 0 FrameStrobe_O[8]
rlabel metal1 42550 8330 42550 8330 0 FrameStrobe_O[9]
rlabel metal1 1012 7990 1012 7990 0 N1BEG[0]
rlabel metal1 1012 7514 1012 7514 0 N1BEG[1]
rlabel metal1 1564 7718 1564 7718 0 N1BEG[2]
rlabel metal1 1380 8058 1380 8058 0 N1BEG[3]
rlabel metal2 1610 9856 1610 9856 0 N2BEG[0]
rlabel metal2 1978 9856 1978 9856 0 N2BEG[1]
rlabel metal2 2346 9856 2346 9856 0 N2BEG[2]
rlabel metal2 2714 9856 2714 9856 0 N2BEG[3]
rlabel metal1 2990 8602 2990 8602 0 N2BEG[4]
rlabel metal2 3450 9856 3450 9856 0 N2BEG[5]
rlabel metal1 3910 8058 3910 8058 0 N2BEG[6]
rlabel metal2 4186 9856 4186 9856 0 N2BEG[7]
rlabel metal2 4554 9856 4554 9856 0 N2BEGb[0]
rlabel metal2 4922 9856 4922 9856 0 N2BEGb[1]
rlabel metal2 5290 9856 5290 9856 0 N2BEGb[2]
rlabel metal2 5658 9856 5658 9856 0 N2BEGb[3]
rlabel metal2 6026 9856 6026 9856 0 N2BEGb[4]
rlabel metal1 6486 8058 6486 8058 0 N2BEGb[5]
rlabel metal2 6762 9856 6762 9856 0 N2BEGb[6]
rlabel metal2 7130 9856 7130 9856 0 N2BEGb[7]
rlabel metal2 7498 9856 7498 9856 0 N4BEG[0]
rlabel metal2 11178 9686 11178 9686 0 N4BEG[10]
rlabel metal1 11960 8058 11960 8058 0 N4BEG[11]
rlabel metal1 11960 8602 11960 8602 0 N4BEG[12]
rlabel metal1 12328 8602 12328 8602 0 N4BEG[13]
rlabel metal1 12696 8602 12696 8602 0 N4BEG[14]
rlabel metal2 13018 9856 13018 9856 0 N4BEG[15]
rlabel metal2 7866 9856 7866 9856 0 N4BEG[1]
rlabel metal2 8234 9856 8234 9856 0 N4BEG[2]
rlabel metal2 8602 9686 8602 9686 0 N4BEG[3]
rlabel metal1 9016 8058 9016 8058 0 N4BEG[4]
rlabel metal2 9338 8432 9338 8432 0 N4BEG[5]
rlabel metal1 9614 8262 9614 8262 0 N4BEG[6]
rlabel metal1 10028 8262 10028 8262 0 N4BEG[7]
rlabel metal2 10442 9686 10442 9686 0 N4BEG[8]
rlabel metal2 10810 9686 10810 9686 0 N4BEG[9]
rlabel metal1 13432 8602 13432 8602 0 NN4BEG[0]
rlabel metal1 17158 8602 17158 8602 0 NN4BEG[10]
rlabel metal1 17526 8602 17526 8602 0 NN4BEG[11]
rlabel metal1 17894 8602 17894 8602 0 NN4BEG[12]
rlabel metal1 18262 8602 18262 8602 0 NN4BEG[13]
rlabel metal1 18630 8602 18630 8602 0 NN4BEG[14]
rlabel metal1 19136 8602 19136 8602 0 NN4BEG[15]
rlabel metal1 13800 8602 13800 8602 0 NN4BEG[1]
rlabel metal2 14398 9591 14398 9591 0 NN4BEG[2]
rlabel metal1 14536 8602 14536 8602 0 NN4BEG[3]
rlabel metal1 14904 8602 14904 8602 0 NN4BEG[4]
rlabel metal1 15364 8602 15364 8602 0 NN4BEG[5]
rlabel metal1 15640 8602 15640 8602 0 NN4BEG[6]
rlabel metal1 16008 8602 16008 8602 0 NN4BEG[7]
rlabel metal1 16376 8602 16376 8602 0 NN4BEG[8]
rlabel metal1 16836 8602 16836 8602 0 NN4BEG[9]
rlabel metal2 19274 10213 19274 10213 0 S1END[0]
rlabel metal1 17618 3502 17618 3502 0 S1END[1]
rlabel metal2 20010 10825 20010 10825 0 S1END[2]
rlabel metal2 17526 3706 17526 3706 0 S1END[3]
rlabel metal2 23690 8938 23690 8938 0 S2END[0]
rlabel metal2 24058 8700 24058 8700 0 S2END[1]
rlabel metal2 24426 8190 24426 8190 0 S2END[2]
rlabel metal2 24794 8156 24794 8156 0 S2END[3]
rlabel metal2 25162 8394 25162 8394 0 S2END[4]
rlabel metal2 25530 8938 25530 8938 0 S2END[5]
rlabel metal2 25898 9516 25898 9516 0 S2END[6]
rlabel metal2 26266 10281 26266 10281 0 S2END[7]
rlabel metal2 20746 11046 20746 11046 0 S2MID[0]
rlabel metal2 20976 4148 20976 4148 0 S2MID[1]
rlabel metal1 19964 4726 19964 4726 0 S2MID[2]
rlabel metal1 20332 4658 20332 4658 0 S2MID[3]
rlabel metal2 22218 8394 22218 8394 0 S2MID[4]
rlabel metal1 19596 6290 19596 6290 0 S2MID[5]
rlabel metal1 20378 6732 20378 6732 0 S2MID[6]
rlabel metal2 23322 9244 23322 9244 0 S2MID[7]
rlabel metal2 26634 11097 26634 11097 0 S4END[0]
rlabel metal2 30314 8989 30314 8989 0 S4END[10]
rlabel metal2 30682 7850 30682 7850 0 S4END[11]
rlabel metal1 32729 5202 32729 5202 0 S4END[12]
rlabel metal2 31418 8394 31418 8394 0 S4END[13]
rlabel metal2 31786 8700 31786 8700 0 S4END[14]
rlabel metal2 32154 11097 32154 11097 0 S4END[15]
rlabel metal2 10166 8551 10166 8551 0 S4END[1]
rlabel metal1 10350 7718 10350 7718 0 S4END[2]
rlabel metal2 15502 9316 15502 9316 0 S4END[3]
rlabel metal2 28106 9482 28106 9482 0 S4END[4]
rlabel metal2 28474 9482 28474 9482 0 S4END[5]
rlabel metal2 28842 9244 28842 9244 0 S4END[6]
rlabel metal2 29210 8700 29210 8700 0 S4END[7]
rlabel metal2 29578 8394 29578 8394 0 S4END[8]
rlabel metal2 29946 9669 29946 9669 0 S4END[9]
rlabel metal2 32522 8768 32522 8768 0 SS4END[0]
rlabel metal1 20286 6698 20286 6698 0 SS4END[10]
rlabel metal1 13340 6766 13340 6766 0 SS4END[11]
rlabel metal1 12696 6766 12696 6766 0 SS4END[12]
rlabel metal2 21390 10064 21390 10064 0 SS4END[13]
rlabel via2 37674 11097 37674 11097 0 SS4END[14]
rlabel metal1 14398 8976 14398 8976 0 SS4END[15]
rlabel metal2 32890 9278 32890 9278 0 SS4END[1]
rlabel metal2 33258 11097 33258 11097 0 SS4END[2]
rlabel metal2 33626 9516 33626 9516 0 SS4END[3]
rlabel metal2 18078 9452 18078 9452 0 SS4END[4]
rlabel metal2 16974 8636 16974 8636 0 SS4END[5]
rlabel metal2 16606 9520 16606 9520 0 SS4END[6]
rlabel metal2 15778 8381 15778 8381 0 SS4END[7]
rlabel metal1 15456 7446 15456 7446 0 SS4END[8]
rlabel metal2 14582 7174 14582 7174 0 SS4END[9]
rlabel metal2 1794 55 1794 55 0 UserCLK
rlabel metal1 38456 8602 38456 8602 0 UserCLKo
rlabel metal2 2162 3264 2162 3264 0 net1
rlabel via2 15318 5627 15318 5627 0 net10
rlabel metal1 14582 6630 14582 6630 0 net100
rlabel metal1 15088 7514 15088 7514 0 net101
rlabel metal1 15686 7514 15686 7514 0 net102
rlabel metal1 16100 8058 16100 8058 0 net103
rlabel metal2 16514 8262 16514 8262 0 net104
rlabel metal1 36846 3162 36846 3162 0 net105
rlabel metal2 25714 4760 25714 4760 0 net11
rlabel metal1 43194 2380 43194 2380 0 net12
rlabel metal1 20516 2822 20516 2822 0 net13
rlabel metal2 17710 3502 17710 3502 0 net14
rlabel metal1 39422 4488 39422 4488 0 net15
rlabel metal1 36570 6290 36570 6290 0 net16
rlabel metal1 42320 6970 42320 6970 0 net17
rlabel metal2 41170 6392 41170 6392 0 net18
rlabel metal1 42182 7446 42182 7446 0 net19
rlabel metal2 25898 3485 25898 3485 0 net2
rlabel metal1 30498 5576 30498 5576 0 net20
rlabel metal2 43930 6460 43930 6460 0 net21
rlabel via2 5290 7803 5290 7803 0 net22
rlabel metal2 19826 2958 19826 2958 0 net23
rlabel metal1 36570 7480 36570 7480 0 net24
rlabel metal2 42826 7446 42826 7446 0 net25
rlabel metal2 40158 2975 40158 2975 0 net26
rlabel metal2 18078 2652 18078 2652 0 net27
rlabel metal1 43286 2312 43286 2312 0 net28
rlabel metal2 40066 3281 40066 3281 0 net29
rlabel metal2 24610 3757 24610 3757 0 net3
rlabel via2 23690 3995 23690 3995 0 net30
rlabel metal2 36570 3740 36570 3740 0 net31
rlabel metal2 20010 4352 20010 4352 0 net32
rlabel metal1 37950 2890 37950 2890 0 net33
rlabel metal2 26726 5610 26726 5610 0 net34
rlabel metal2 40066 8466 40066 8466 0 net35
rlabel metal1 36294 3060 36294 3060 0 net36
rlabel metal2 40802 8500 40802 8500 0 net37
rlabel metal1 43884 7854 43884 7854 0 net38
rlabel metal2 36662 7616 36662 7616 0 net39
rlabel metal2 41078 4794 41078 4794 0 net4
rlabel metal2 42182 7242 42182 7242 0 net40
rlabel metal2 41262 7548 41262 7548 0 net41
rlabel metal2 44298 6630 44298 6630 0 net42
rlabel metal1 43562 6732 43562 6732 0 net43
rlabel metal2 38318 5780 38318 5780 0 net44
rlabel metal2 20930 3400 20930 3400 0 net45
rlabel metal2 9982 3400 9982 3400 0 net46
rlabel metal1 18262 2924 18262 2924 0 net47
rlabel metal1 21298 3060 21298 3060 0 net48
rlabel metal1 19320 2822 19320 2822 0 net49
rlabel metal2 21942 6188 21942 6188 0 net5
rlabel metal1 20194 3400 20194 3400 0 net50
rlabel metal2 39974 5848 39974 5848 0 net51
rlabel metal2 32706 6086 32706 6086 0 net52
rlabel metal2 2346 7378 2346 7378 0 net53
rlabel metal1 2231 7378 2231 7378 0 net54
rlabel metal2 2438 7412 2438 7412 0 net55
rlabel metal1 1702 7888 1702 7888 0 net56
rlabel metal1 1794 8398 1794 8398 0 net57
rlabel metal1 20194 6664 20194 6664 0 net58
rlabel metal1 19366 6188 19366 6188 0 net59
rlabel metal2 19090 5678 19090 5678 0 net6
rlabel metal1 14858 5848 14858 5848 0 net60
rlabel metal2 11454 6851 11454 6851 0 net61
rlabel metal2 8326 6766 8326 6766 0 net62
rlabel metal2 17986 5508 17986 5508 0 net63
rlabel metal2 10350 6596 10350 6596 0 net64
rlabel metal2 14674 7616 14674 7616 0 net65
rlabel metal2 20378 8143 20378 8143 0 net66
rlabel metal1 12650 8466 12650 8466 0 net67
rlabel metal1 16560 5644 16560 5644 0 net68
rlabel metal2 6210 6732 6210 6732 0 net69
rlabel metal1 44298 5270 44298 5270 0 net7
rlabel metal2 9798 6562 9798 6562 0 net70
rlabel metal1 16560 6392 16560 6392 0 net71
rlabel metal2 7314 7004 7314 7004 0 net72
rlabel metal3 16560 7208 16560 7208 0 net73
rlabel metal2 22034 7888 22034 7888 0 net74
rlabel metal1 21390 8024 21390 8024 0 net75
rlabel metal1 10166 7514 10166 7514 0 net76
rlabel metal1 10120 7990 10120 7990 0 net77
rlabel metal1 10442 7956 10442 7956 0 net78
rlabel metal1 13202 8500 13202 8500 0 net79
rlabel metal2 20470 5984 20470 5984 0 net8
rlabel metal3 16560 6256 16560 6256 0 net80
rlabel metal2 14950 6630 14950 6630 0 net81
rlabel metal2 14582 5304 14582 5304 0 net82
rlabel metal2 9522 6188 9522 6188 0 net83
rlabel metal2 9890 6001 9890 6001 0 net84
rlabel metal2 31142 7140 31142 7140 0 net85
rlabel metal2 14858 6324 14858 6324 0 net86
rlabel metal1 19182 6120 19182 6120 0 net87
rlabel metal2 10994 7854 10994 7854 0 net88
rlabel metal2 13294 8126 13294 8126 0 net89
rlabel metal2 27278 5916 27278 5916 0 net9
rlabel metal1 17342 8058 17342 8058 0 net90
rlabel metal1 17848 8058 17848 8058 0 net91
rlabel metal2 18170 8364 18170 8364 0 net92
rlabel via1 19366 7939 19366 7939 0 net93
rlabel metal2 18906 7888 18906 7888 0 net94
rlabel metal1 20102 8466 20102 8466 0 net95
rlabel metal1 12466 8024 12466 8024 0 net96
rlabel metal2 12650 7684 12650 7684 0 net97
rlabel metal1 13340 8330 13340 8330 0 net98
rlabel metal1 14168 6834 14168 6834 0 net99
<< properties >>
string FIXED_BBOX 0 0 46000 11152
<< end >>
