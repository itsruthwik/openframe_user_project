magic
tech sky130A
magscale 1 2
timestamp 1746698478
<< viali >>
rect 2697 8585 2731 8619
rect 3065 8585 3099 8619
rect 4169 8585 4203 8619
rect 4537 8585 4571 8619
rect 4905 8585 4939 8619
rect 5273 8585 5307 8619
rect 5733 8585 5767 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 7941 8585 7975 8619
rect 8217 8585 8251 8619
rect 8585 8585 8619 8619
rect 9321 8585 9355 8619
rect 9689 8585 9723 8619
rect 10057 8585 10091 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 11161 8585 11195 8619
rect 11897 8585 11931 8619
rect 12265 8585 12299 8619
rect 12633 8585 12667 8619
rect 13001 8585 13035 8619
rect 13737 8585 13771 8619
rect 14473 8585 14507 8619
rect 14841 8585 14875 8619
rect 15209 8585 15243 8619
rect 15577 8585 15611 8619
rect 15945 8585 15979 8619
rect 16313 8585 16347 8619
rect 17049 8585 17083 8619
rect 31585 8585 31619 8619
rect 32321 8585 32355 8619
rect 33057 8585 33091 8619
rect 33425 8585 33459 8619
rect 34897 8585 34931 8619
rect 36001 8585 36035 8619
rect 37473 8585 37507 8619
rect 37841 8585 37875 8619
rect 2881 8449 2915 8483
rect 3249 8449 3283 8483
rect 3617 8449 3651 8483
rect 4353 8449 4387 8483
rect 4721 8449 4755 8483
rect 5101 8449 5135 8483
rect 5450 8449 5484 8483
rect 5549 8449 5583 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 7757 8449 7791 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10253 8449 10287 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 11345 8449 11379 8483
rect 12081 8449 12115 8483
rect 12449 8449 12483 8483
rect 12817 8449 12851 8483
rect 13185 8449 13219 8483
rect 13553 8449 13587 8483
rect 13933 8449 13967 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 15393 8449 15427 8483
rect 15761 8449 15795 8483
rect 16129 8449 16163 8483
rect 16497 8449 16531 8483
rect 17233 8449 17267 8483
rect 17601 8449 17635 8483
rect 31769 8449 31803 8483
rect 32137 8449 32171 8483
rect 32505 8449 32539 8483
rect 32873 8449 32907 8483
rect 33241 8449 33275 8483
rect 33609 8449 33643 8483
rect 33977 8449 34011 8483
rect 34713 8449 34747 8483
rect 35081 8449 35115 8483
rect 35449 8449 35483 8483
rect 35817 8449 35851 8483
rect 36185 8449 36219 8483
rect 36553 8449 36587 8483
rect 37289 8449 37323 8483
rect 37657 8449 37691 8483
rect 38209 8449 38243 8483
rect 3433 8313 3467 8347
rect 13369 8313 13403 8347
rect 17417 8313 17451 8347
rect 32689 8313 32723 8347
rect 33793 8313 33827 8347
rect 34161 8313 34195 8347
rect 35265 8313 35299 8347
rect 35633 8313 35667 8347
rect 36369 8313 36403 8347
rect 36737 8313 36771 8347
rect 38393 8313 38427 8347
rect 3249 8041 3283 8075
rect 3893 8041 3927 8075
rect 4353 8041 4387 8075
rect 5457 8041 5491 8075
rect 6285 8041 6319 8075
rect 6837 8041 6871 8075
rect 7665 8041 7699 8075
rect 8493 8041 8527 8075
rect 9321 8041 9355 8075
rect 9873 8041 9907 8075
rect 10977 8041 11011 8075
rect 11529 8041 11563 8075
rect 12081 8041 12115 8075
rect 13185 8041 13219 8075
rect 13737 8041 13771 8075
rect 14565 8041 14599 8075
rect 15393 8041 15427 8075
rect 33701 8041 33735 8075
rect 34069 8041 34103 8075
rect 35081 8041 35115 8075
rect 36185 8041 36219 8075
rect 36553 8041 36587 8075
rect 36921 8041 36955 8075
rect 37289 8041 37323 8075
rect 37657 8041 37691 8075
rect 3433 7837 3467 7871
rect 4077 7837 4111 7871
rect 4537 7837 4571 7871
rect 5641 7837 5675 7871
rect 6469 7837 6503 7871
rect 7021 7837 7055 7871
rect 7849 7837 7883 7871
rect 8677 7837 8711 7871
rect 9505 7837 9539 7871
rect 10057 7837 10091 7871
rect 11161 7837 11195 7871
rect 11713 7837 11747 7871
rect 12265 7837 12299 7871
rect 13369 7837 13403 7871
rect 13921 7837 13955 7871
rect 14749 7837 14783 7871
rect 15577 7837 15611 7871
rect 33517 7837 33551 7871
rect 33885 7837 33919 7871
rect 34897 7837 34931 7871
rect 36001 7837 36035 7871
rect 36369 7837 36403 7871
rect 36737 7837 36771 7871
rect 37105 7837 37139 7871
rect 37473 7837 37507 7871
rect 37841 7837 37875 7871
rect 38209 7837 38243 7871
rect 38025 7701 38059 7735
rect 38393 7701 38427 7735
rect 5181 7497 5215 7531
rect 5457 7497 5491 7531
rect 5733 7497 5767 7531
rect 6009 7497 6043 7531
rect 6837 7497 6871 7531
rect 7113 7497 7147 7531
rect 7665 7497 7699 7531
rect 14197 7497 14231 7531
rect 14933 7497 14967 7531
rect 15393 7497 15427 7531
rect 15761 7497 15795 7531
rect 16773 7497 16807 7531
rect 17049 7497 17083 7531
rect 19901 7497 19935 7531
rect 22293 7497 22327 7531
rect 22477 7497 22511 7531
rect 22845 7497 22879 7531
rect 28825 7497 28859 7531
rect 37657 7497 37691 7531
rect 38025 7497 38059 7531
rect 5365 7361 5399 7395
rect 5641 7361 5675 7395
rect 5917 7361 5951 7395
rect 6193 7361 6227 7395
rect 6745 7361 6779 7395
rect 7021 7361 7055 7395
rect 7297 7361 7331 7395
rect 7849 7361 7883 7395
rect 13001 7361 13035 7395
rect 13277 7361 13311 7395
rect 14105 7361 14139 7395
rect 14381 7361 14415 7395
rect 14657 7361 14691 7395
rect 15117 7361 15151 7395
rect 15577 7361 15611 7395
rect 15945 7361 15979 7395
rect 16957 7361 16991 7395
rect 17233 7361 17267 7395
rect 18797 7361 18831 7395
rect 18889 7361 18923 7395
rect 19717 7361 19751 7395
rect 19993 7361 20027 7395
rect 20361 7361 20395 7395
rect 20545 7361 20579 7395
rect 20637 7361 20671 7395
rect 20913 7361 20947 7395
rect 21281 7361 21315 7395
rect 21557 7361 21591 7395
rect 21833 7361 21867 7395
rect 22109 7361 22143 7395
rect 22569 7361 22603 7395
rect 22661 7361 22695 7395
rect 22937 7361 22971 7395
rect 23213 7361 23247 7395
rect 24409 7361 24443 7395
rect 29009 7361 29043 7395
rect 29469 7361 29503 7395
rect 29745 7361 29779 7395
rect 30021 7361 30055 7395
rect 30297 7361 30331 7395
rect 36829 7361 36863 7395
rect 37473 7361 37507 7395
rect 37841 7361 37875 7395
rect 38209 7361 38243 7395
rect 6561 7225 6595 7259
rect 13093 7225 13127 7259
rect 14473 7225 14507 7259
rect 20453 7225 20487 7259
rect 20821 7225 20855 7259
rect 21097 7225 21131 7259
rect 24225 7225 24259 7259
rect 37013 7225 37047 7259
rect 13921 7157 13955 7191
rect 18705 7157 18739 7191
rect 19073 7157 19107 7191
rect 20177 7157 20211 7191
rect 21465 7157 21499 7191
rect 22017 7157 22051 7191
rect 23121 7157 23155 7191
rect 29285 7157 29319 7191
rect 29561 7157 29595 7191
rect 29837 7157 29871 7191
rect 30113 7157 30147 7191
rect 38393 7157 38427 7191
rect 8309 6953 8343 6987
rect 9965 6953 9999 6987
rect 13645 6953 13679 6987
rect 9597 6885 9631 6919
rect 13093 6885 13127 6919
rect 14381 6885 14415 6919
rect 19717 6885 19751 6919
rect 25697 6885 25731 6919
rect 25973 6885 26007 6919
rect 26893 6885 26927 6919
rect 22201 6817 22235 6851
rect 22753 6817 22787 6851
rect 6469 6749 6503 6783
rect 7389 6749 7423 6783
rect 7757 6749 7791 6783
rect 8033 6749 8067 6783
rect 8493 6749 8527 6783
rect 8769 6749 8803 6783
rect 9229 6749 9263 6783
rect 9505 6749 9539 6783
rect 9781 6749 9815 6783
rect 10149 6749 10183 6783
rect 10425 6749 10459 6783
rect 13001 6749 13035 6783
rect 13277 6749 13311 6783
rect 13553 6749 13587 6783
rect 13829 6749 13863 6783
rect 14289 6749 14323 6783
rect 14565 6749 14599 6783
rect 17969 6749 18003 6783
rect 19441 6749 19475 6783
rect 19533 6749 19567 6783
rect 20269 6749 20303 6783
rect 20361 6749 20395 6783
rect 21005 6749 21039 6783
rect 21189 6749 21223 6783
rect 22293 6749 22327 6783
rect 22385 6749 22419 6783
rect 22845 6749 22879 6783
rect 22937 6749 22971 6783
rect 25605 6749 25639 6783
rect 25881 6749 25915 6783
rect 26157 6749 26191 6783
rect 26433 6749 26467 6783
rect 27077 6749 27111 6783
rect 27353 6749 27387 6783
rect 27629 6749 27663 6783
rect 28089 6749 28123 6783
rect 28365 6749 28399 6783
rect 28733 6749 28767 6783
rect 37473 6749 37507 6783
rect 37841 6749 37875 6783
rect 38209 6749 38243 6783
rect 20177 6681 20211 6715
rect 6285 6613 6319 6647
rect 7573 6613 7607 6647
rect 7849 6613 7883 6647
rect 8585 6613 8619 6647
rect 9321 6613 9355 6647
rect 10241 6613 10275 6647
rect 12817 6613 12851 6647
rect 13369 6613 13403 6647
rect 14105 6613 14139 6647
rect 17785 6613 17819 6647
rect 18153 6613 18187 6647
rect 19349 6613 19383 6647
rect 20545 6613 20579 6647
rect 21373 6613 21407 6647
rect 22569 6613 22603 6647
rect 23121 6613 23155 6647
rect 25421 6613 25455 6647
rect 26249 6613 26283 6647
rect 27169 6613 27203 6647
rect 27445 6613 27479 6647
rect 27905 6613 27939 6647
rect 28181 6613 28215 6647
rect 28549 6613 28583 6647
rect 37657 6613 37691 6647
rect 38025 6613 38059 6647
rect 38393 6613 38427 6647
rect 10241 6409 10275 6443
rect 10609 6409 10643 6443
rect 13185 6409 13219 6443
rect 17049 6409 17083 6443
rect 28457 6409 28491 6443
rect 29469 6409 29503 6443
rect 38393 6409 38427 6443
rect 8309 6273 8343 6307
rect 10417 6273 10451 6307
rect 10793 6273 10827 6307
rect 13369 6273 13403 6307
rect 16773 6273 16807 6307
rect 16865 6273 16899 6307
rect 22293 6273 22327 6307
rect 28273 6273 28307 6307
rect 29285 6273 29319 6307
rect 37841 6273 37875 6307
rect 38209 6273 38243 6307
rect 38025 6137 38059 6171
rect 8125 6069 8159 6103
rect 10149 6069 10183 6103
rect 22477 6069 22511 6103
rect 31401 5865 31435 5899
rect 34897 5865 34931 5899
rect 37105 5865 37139 5899
rect 37381 5865 37415 5899
rect 28365 5797 28399 5831
rect 33333 5797 33367 5831
rect 36093 5797 36127 5831
rect 38393 5797 38427 5831
rect 28181 5661 28215 5695
rect 31217 5661 31251 5695
rect 33149 5661 33183 5695
rect 34713 5661 34747 5695
rect 35909 5661 35943 5695
rect 36921 5661 36955 5695
rect 37189 5661 37223 5695
rect 37841 5661 37875 5695
rect 38209 5661 38243 5695
rect 38025 5525 38059 5559
rect 38393 5321 38427 5355
rect 19625 5185 19659 5219
rect 19717 5185 19751 5219
rect 28089 5185 28123 5219
rect 37841 5185 37875 5219
rect 38209 5185 38243 5219
rect 19901 5049 19935 5083
rect 28273 4981 28307 5015
rect 38025 4981 38059 5015
rect 38393 4709 38427 4743
rect 21925 4641 21959 4675
rect 21281 4573 21315 4607
rect 21373 4573 21407 4607
rect 22017 4573 22051 4607
rect 22109 4573 22143 4607
rect 37841 4573 37875 4607
rect 38209 4573 38243 4607
rect 21189 4505 21223 4539
rect 21557 4437 21591 4471
rect 22293 4437 22327 4471
rect 38025 4437 38059 4471
rect 15393 4233 15427 4267
rect 15209 4097 15243 4131
rect 15485 4097 15519 4131
rect 16129 4097 16163 4131
rect 16497 4097 16531 4131
rect 16681 4097 16715 4131
rect 17049 4097 17083 4131
rect 17509 4097 17543 4131
rect 17601 4097 17635 4131
rect 18337 4097 18371 4131
rect 18429 4097 18463 4131
rect 18705 4097 18739 4131
rect 18981 4097 19015 4131
rect 19441 4097 19475 4131
rect 20453 4097 20487 4131
rect 21189 4097 21223 4131
rect 21281 4097 21315 4131
rect 21833 4097 21867 4131
rect 22293 4097 22327 4131
rect 22385 4097 22419 4131
rect 22661 4097 22695 4131
rect 22937 4097 22971 4131
rect 26985 4097 27019 4131
rect 37841 4097 37875 4131
rect 38209 4097 38243 4131
rect 17877 3961 17911 3995
rect 18613 3961 18647 3995
rect 21465 3961 21499 3995
rect 22017 3961 22051 3995
rect 38393 3961 38427 3995
rect 15669 3893 15703 3927
rect 16313 3893 16347 3927
rect 16405 3893 16439 3927
rect 16865 3893 16899 3927
rect 17233 3893 17267 3927
rect 17417 3893 17451 3927
rect 17785 3893 17819 3927
rect 18245 3893 18279 3927
rect 18889 3893 18923 3927
rect 19625 3893 19659 3927
rect 20637 3893 20671 3927
rect 21097 3893 21131 3927
rect 21557 3893 21591 3927
rect 22201 3893 22235 3927
rect 22569 3893 22603 3927
rect 22845 3893 22879 3927
rect 27169 3893 27203 3927
rect 38025 3893 38059 3927
rect 18061 3689 18095 3723
rect 26893 3621 26927 3655
rect 27445 3621 27479 3655
rect 38393 3621 38427 3655
rect 17877 3485 17911 3519
rect 21741 3485 21775 3519
rect 21925 3485 21959 3519
rect 25329 3485 25363 3519
rect 25421 3485 25455 3519
rect 26157 3485 26191 3519
rect 26617 3485 26651 3519
rect 26709 3485 26743 3519
rect 26985 3485 27019 3519
rect 27261 3485 27295 3519
rect 37841 3485 37875 3519
rect 38209 3485 38243 3519
rect 22109 3349 22143 3383
rect 25237 3349 25271 3383
rect 25605 3349 25639 3383
rect 26341 3349 26375 3383
rect 26525 3349 26559 3383
rect 27169 3349 27203 3383
rect 38025 3349 38059 3383
rect 38393 3145 38427 3179
rect 37473 3009 37507 3043
rect 37841 3009 37875 3043
rect 38209 3009 38243 3043
rect 37657 2805 37691 2839
rect 38025 2805 38059 2839
rect 36645 2533 36679 2567
rect 37013 2533 37047 2567
rect 38393 2533 38427 2567
rect 36461 2397 36495 2431
rect 36829 2397 36863 2431
rect 37473 2397 37507 2431
rect 37841 2397 37875 2431
rect 38209 2397 38243 2431
rect 37657 2261 37691 2295
rect 38025 2261 38059 2295
<< metal1 >>
rect 10428 11104 22232 11132
rect 10428 11076 10456 11104
rect 22204 11076 22232 11104
rect 10410 11024 10416 11076
rect 10468 11024 10474 11076
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11020 11036 22094 11064
rect 11020 11024 11026 11036
rect 7374 10956 7380 11008
rect 7432 10996 7438 11008
rect 17954 10996 17960 11008
rect 7432 10968 17960 10996
rect 7432 10956 7438 10968
rect 17954 10956 17960 10968
rect 18012 10956 18018 11008
rect 22066 10996 22094 11036
rect 22186 11024 22192 11076
rect 22244 11024 22250 11076
rect 22370 10996 22376 11008
rect 22066 10968 22376 10996
rect 22370 10956 22376 10968
rect 22428 10956 22434 11008
rect 11422 10888 11428 10940
rect 11480 10928 11486 10940
rect 21542 10928 21548 10940
rect 11480 10900 21548 10928
rect 11480 10888 11486 10900
rect 21542 10888 21548 10900
rect 21600 10888 21606 10940
rect 14458 10820 14464 10872
rect 14516 10860 14522 10872
rect 23198 10860 23204 10872
rect 14516 10832 23204 10860
rect 14516 10820 14522 10832
rect 23198 10820 23204 10832
rect 23256 10820 23262 10872
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 20714 10792 20720 10804
rect 11572 10764 20720 10792
rect 11572 10752 11578 10764
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 23382 10140 23388 10192
rect 23440 10180 23446 10192
rect 25958 10180 25964 10192
rect 23440 10152 25964 10180
rect 23440 10140 23446 10152
rect 25958 10140 25964 10152
rect 26016 10140 26022 10192
rect 21542 10072 21548 10124
rect 21600 10112 21606 10124
rect 24578 10112 24584 10124
rect 21600 10084 24584 10112
rect 21600 10072 21606 10084
rect 24578 10072 24584 10084
rect 24636 10072 24642 10124
rect 25866 10004 25872 10056
rect 25924 10044 25930 10056
rect 31202 10044 31208 10056
rect 25924 10016 31208 10044
rect 25924 10004 25930 10016
rect 31202 10004 31208 10016
rect 31260 10004 31266 10056
rect 13354 9936 13360 9988
rect 13412 9976 13418 9988
rect 18506 9976 18512 9988
rect 13412 9948 18512 9976
rect 13412 9936 13418 9948
rect 18506 9936 18512 9948
rect 18564 9936 18570 9988
rect 13630 9868 13636 9920
rect 13688 9908 13694 9920
rect 17678 9908 17684 9920
rect 13688 9880 17684 9908
rect 13688 9868 13694 9880
rect 17678 9868 17684 9880
rect 17736 9868 17742 9920
rect 25590 9868 25596 9920
rect 25648 9908 25654 9920
rect 30926 9908 30932 9920
rect 25648 9880 30932 9908
rect 25648 9868 25654 9880
rect 30926 9868 30932 9880
rect 30984 9868 30990 9920
rect 16666 9800 16672 9852
rect 16724 9840 16730 9852
rect 25682 9840 25688 9852
rect 16724 9812 25688 9840
rect 16724 9800 16730 9812
rect 25682 9800 25688 9812
rect 25740 9800 25746 9852
rect 13906 9732 13912 9784
rect 13964 9772 13970 9784
rect 18782 9772 18788 9784
rect 13964 9744 18788 9772
rect 13964 9732 13970 9744
rect 18782 9732 18788 9744
rect 18840 9732 18846 9784
rect 30374 9772 30380 9784
rect 25700 9744 30380 9772
rect 25700 9716 25728 9744
rect 30374 9732 30380 9744
rect 30432 9732 30438 9784
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 21818 9704 21824 9716
rect 1360 9676 21824 9704
rect 1360 9664 1366 9676
rect 21818 9664 21824 9676
rect 21876 9664 21882 9716
rect 25682 9664 25688 9716
rect 25740 9664 25746 9716
rect 25774 9664 25780 9716
rect 25832 9704 25838 9716
rect 30650 9704 30656 9716
rect 25832 9676 30656 9704
rect 25832 9664 25838 9676
rect 30650 9664 30656 9676
rect 30708 9664 30714 9716
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 17402 9568 17408 9580
rect 14608 9540 17408 9568
rect 14608 9528 14614 9540
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 14182 9392 14188 9444
rect 14240 9432 14246 9444
rect 26602 9432 26608 9444
rect 14240 9404 26608 9432
rect 14240 9392 14246 9404
rect 26602 9392 26608 9404
rect 26660 9392 26666 9444
rect 16114 9324 16120 9376
rect 16172 9364 16178 9376
rect 28810 9364 28816 9376
rect 16172 9336 28816 9364
rect 16172 9324 16178 9336
rect 28810 9324 28816 9336
rect 28868 9324 28874 9376
rect 10686 9256 10692 9308
rect 10744 9296 10750 9308
rect 15838 9296 15844 9308
rect 10744 9268 15844 9296
rect 10744 9256 10750 9268
rect 15838 9256 15844 9268
rect 15896 9256 15902 9308
rect 15930 9256 15936 9308
rect 15988 9296 15994 9308
rect 28902 9296 28908 9308
rect 15988 9268 28908 9296
rect 15988 9256 15994 9268
rect 28902 9256 28908 9268
rect 28960 9256 28966 9308
rect 11974 9188 11980 9240
rect 12032 9228 12038 9240
rect 13906 9228 13912 9240
rect 12032 9200 13912 9228
rect 12032 9188 12038 9200
rect 13906 9188 13912 9200
rect 13964 9188 13970 9240
rect 15654 9188 15660 9240
rect 15712 9228 15718 9240
rect 29362 9228 29368 9240
rect 15712 9200 29368 9228
rect 15712 9188 15718 9200
rect 29362 9188 29368 9200
rect 29420 9188 29426 9240
rect 1118 9120 1124 9172
rect 1176 9160 1182 9172
rect 22094 9160 22100 9172
rect 1176 9132 22100 9160
rect 1176 9120 1182 9132
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 27430 9120 27436 9172
rect 27488 9160 27494 9172
rect 34882 9160 34888 9172
rect 27488 9132 34888 9160
rect 27488 9120 27494 9132
rect 34882 9120 34888 9132
rect 34940 9120 34946 9172
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 17034 9092 17040 9104
rect 8444 9064 17040 9092
rect 8444 9052 8450 9064
rect 17034 9052 17040 9064
rect 17092 9052 17098 9104
rect 24670 9052 24676 9104
rect 24728 9092 24734 9104
rect 32122 9092 32128 9104
rect 24728 9064 32128 9092
rect 24728 9052 24734 9064
rect 32122 9052 32128 9064
rect 32180 9052 32186 9104
rect 13170 8984 13176 9036
rect 13228 9024 13234 9036
rect 15562 9024 15568 9036
rect 13228 8996 15568 9024
rect 13228 8984 13234 8996
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 19886 9024 19892 9036
rect 16264 8996 19892 9024
rect 16264 8984 16270 8996
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 28442 8984 28448 9036
rect 28500 9024 28506 9036
rect 35802 9024 35808 9036
rect 28500 8996 35808 9024
rect 28500 8984 28506 8996
rect 35802 8984 35808 8996
rect 35860 8984 35866 9036
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 18230 8956 18236 8968
rect 7892 8928 18236 8956
rect 7892 8916 7898 8928
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 22278 8916 22284 8968
rect 22336 8956 22342 8968
rect 38194 8956 38200 8968
rect 22336 8928 38200 8956
rect 22336 8916 22342 8928
rect 38194 8916 38200 8928
rect 38252 8916 38258 8968
rect 4246 8848 4252 8900
rect 4304 8888 4310 8900
rect 10134 8888 10140 8900
rect 4304 8860 10140 8888
rect 4304 8848 4310 8860
rect 10134 8848 10140 8860
rect 10192 8848 10198 8900
rect 12802 8848 12808 8900
rect 12860 8888 12866 8900
rect 24210 8888 24216 8900
rect 12860 8860 24216 8888
rect 12860 8848 12866 8860
rect 24210 8848 24216 8860
rect 24268 8848 24274 8900
rect 31846 8848 31852 8900
rect 31904 8888 31910 8900
rect 33594 8888 33600 8900
rect 31904 8860 33600 8888
rect 31904 8848 31910 8860
rect 33594 8848 33600 8860
rect 33652 8848 33658 8900
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 6454 8820 6460 8832
rect 4948 8792 6460 8820
rect 4948 8780 4954 8792
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 9490 8780 9496 8832
rect 9548 8820 9554 8832
rect 14826 8820 14832 8832
rect 9548 8792 14832 8820
rect 9548 8780 9554 8792
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 19610 8820 19616 8832
rect 17644 8792 19616 8820
rect 17644 8780 17650 8792
rect 19610 8780 19616 8792
rect 19668 8780 19674 8832
rect 33134 8780 33140 8832
rect 33192 8820 33198 8832
rect 34146 8820 34152 8832
rect 33192 8792 34152 8820
rect 33192 8780 33198 8792
rect 34146 8780 34152 8792
rect 34204 8780 34210 8832
rect 35342 8780 35348 8832
rect 35400 8820 35406 8832
rect 35710 8820 35716 8832
rect 35400 8792 35716 8820
rect 35400 8780 35406 8792
rect 35710 8780 35716 8792
rect 35768 8780 35774 8832
rect 1104 8730 38824 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 38824 8730
rect 1104 8656 38824 8678
rect 2685 8619 2743 8625
rect 2685 8585 2697 8619
rect 2731 8616 2743 8619
rect 2774 8616 2780 8628
rect 2731 8588 2780 8616
rect 2731 8585 2743 8588
rect 2685 8579 2743 8585
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 3053 8619 3111 8625
rect 3053 8585 3065 8619
rect 3099 8616 3111 8619
rect 3418 8616 3424 8628
rect 3099 8588 3424 8616
rect 3099 8585 3111 8588
rect 3053 8579 3111 8585
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4430 8616 4436 8628
rect 4203 8588 4436 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4706 8616 4712 8628
rect 4571 8588 4712 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 4982 8616 4988 8628
rect 4939 8588 4988 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 5534 8616 5540 8628
rect 5307 8588 5540 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5810 8616 5816 8628
rect 5767 8588 5816 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6362 8616 6368 8628
rect 6043 8588 6368 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 6914 8616 6920 8628
rect 6779 8588 6920 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7190 8616 7196 8628
rect 7147 8588 7196 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7742 8616 7748 8628
rect 7515 8588 7748 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8018 8616 8024 8628
rect 7975 8588 8024 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8478 8616 8484 8628
rect 8251 8588 8484 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 8754 8616 8760 8628
rect 8619 8588 8760 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9398 8616 9404 8628
rect 9355 8588 9404 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 9950 8616 9956 8628
rect 9723 8588 9956 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10226 8616 10232 8628
rect 10091 8588 10232 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10502 8616 10508 8628
rect 10459 8588 10508 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 11054 8616 11060 8628
rect 10827 8588 11060 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11606 8616 11612 8628
rect 11195 8588 11612 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12158 8616 12164 8628
rect 11931 8588 12164 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12434 8616 12440 8628
rect 12299 8588 12440 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12621 8619 12679 8625
rect 12621 8585 12633 8619
rect 12667 8616 12679 8619
rect 12710 8616 12716 8628
rect 12667 8588 12716 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 12989 8619 13047 8625
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13262 8616 13268 8628
rect 13035 8588 13268 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 14090 8616 14096 8628
rect 13771 8588 14096 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 14461 8619 14519 8625
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14642 8616 14648 8628
rect 14507 8588 14648 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14642 8576 14648 8588
rect 14700 8576 14706 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 14918 8616 14924 8628
rect 14875 8588 14924 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15470 8616 15476 8628
rect 15243 8588 15476 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15746 8616 15752 8628
rect 15611 8588 15752 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16022 8616 16028 8628
rect 15979 8588 16028 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16022 8576 16028 8588
rect 16080 8576 16086 8628
rect 16298 8576 16304 8628
rect 16356 8576 16362 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16908 8588 17049 8616
rect 16908 8576 16914 8588
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 17420 8588 17632 8616
rect 6822 8548 6828 8560
rect 5368 8520 6828 8548
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 4246 8480 4252 8492
rect 3651 8452 4252 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 1210 8304 1216 8356
rect 1268 8344 1274 8356
rect 1670 8344 1676 8356
rect 1268 8316 1676 8344
rect 1268 8304 1274 8316
rect 1670 8304 1676 8316
rect 1728 8304 1734 8356
rect 2884 8344 2912 8443
rect 3252 8412 3280 8443
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8480 4767 8483
rect 4890 8480 4896 8492
rect 4755 8452 4896 8480
rect 4755 8449 4767 8452
rect 4709 8443 4767 8449
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5089 8483 5147 8489
rect 5089 8449 5101 8483
rect 5135 8480 5147 8483
rect 5368 8480 5396 8520
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 10686 8548 10692 8560
rect 8772 8520 10692 8548
rect 5442 8489 5448 8492
rect 5135 8452 5396 8480
rect 5135 8449 5147 8452
rect 5089 8443 5147 8449
rect 5438 8443 5448 8489
rect 5442 8440 5448 8443
rect 5500 8440 5506 8492
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8480 6975 8483
rect 7190 8480 7196 8492
rect 6963 8452 7196 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 5350 8412 5356 8424
rect 3252 8384 5356 8412
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 6196 8412 6224 8443
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 6196 8384 7512 8412
rect 3421 8347 3479 8353
rect 2884 8316 3372 8344
rect 3344 8276 3372 8316
rect 3421 8313 3433 8347
rect 3467 8344 3479 8347
rect 3878 8344 3884 8356
rect 3467 8316 3884 8344
rect 3467 8313 3479 8316
rect 3421 8307 3479 8313
rect 3878 8304 3884 8316
rect 3936 8304 3942 8356
rect 6362 8344 6368 8356
rect 3988 8316 6368 8344
rect 3988 8276 4016 8316
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 7484 8344 7512 8384
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 7760 8412 7788 8443
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8772 8489 8800 8520
rect 10686 8508 10692 8520
rect 10744 8508 10750 8560
rect 14274 8548 14280 8560
rect 12084 8520 14280 8548
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 10241 8483 10299 8489
rect 10241 8449 10253 8483
rect 10287 8480 10299 8483
rect 10287 8452 10364 8480
rect 10287 8449 10299 8452
rect 10241 8443 10299 8449
rect 7616 8384 7788 8412
rect 7616 8372 7622 8384
rect 9582 8344 9588 8356
rect 7484 8316 9588 8344
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 9876 8344 9904 8443
rect 10336 8344 10364 8452
rect 10594 8440 10600 8492
rect 10652 8440 10658 8492
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11238 8480 11244 8492
rect 11011 8452 11244 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 11790 8480 11796 8492
rect 11379 8452 11796 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 12084 8489 12112 8520
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 17420 8548 17448 8588
rect 14660 8520 16344 8548
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12452 8412 12480 8443
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 13170 8440 13176 8492
rect 13228 8440 13234 8492
rect 14660 8489 14688 8520
rect 16316 8492 16344 8520
rect 16500 8520 17448 8548
rect 17604 8548 17632 8588
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 25406 8616 25412 8628
rect 17736 8588 25412 8616
rect 17736 8576 17742 8588
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 31478 8576 31484 8628
rect 31536 8616 31542 8628
rect 31573 8619 31631 8625
rect 31573 8616 31585 8619
rect 31536 8588 31585 8616
rect 31536 8576 31542 8588
rect 31573 8585 31585 8588
rect 31619 8585 31631 8619
rect 31573 8579 31631 8585
rect 31754 8576 31760 8628
rect 31812 8616 31818 8628
rect 32309 8619 32367 8625
rect 32309 8616 32321 8619
rect 31812 8588 32321 8616
rect 31812 8576 31818 8588
rect 32309 8585 32321 8588
rect 32355 8585 32367 8619
rect 32309 8579 32367 8585
rect 32398 8576 32404 8628
rect 32456 8616 32462 8628
rect 33045 8619 33103 8625
rect 33045 8616 33057 8619
rect 32456 8588 33057 8616
rect 32456 8576 32462 8588
rect 33045 8585 33057 8588
rect 33091 8585 33103 8619
rect 33045 8579 33103 8585
rect 33413 8619 33471 8625
rect 33413 8585 33425 8619
rect 33459 8585 33471 8619
rect 33413 8579 33471 8585
rect 27982 8548 27988 8560
rect 17604 8520 27988 8548
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8480 13599 8483
rect 13921 8483 13979 8489
rect 13587 8452 13860 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 13446 8412 13452 8424
rect 12452 8384 13452 8412
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 13832 8412 13860 8452
rect 13921 8449 13933 8483
rect 13967 8480 13979 8483
rect 14645 8483 14703 8489
rect 13967 8452 14044 8480
rect 13967 8449 13979 8452
rect 13921 8443 13979 8449
rect 14016 8412 14044 8452
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8480 15439 8483
rect 15654 8480 15660 8492
rect 15427 8452 15660 8480
rect 15427 8449 15439 8452
rect 15381 8443 15439 8449
rect 14182 8412 14188 8424
rect 13832 8384 13952 8412
rect 14016 8384 14188 8412
rect 13170 8344 13176 8356
rect 9876 8316 10272 8344
rect 10336 8316 13176 8344
rect 3344 8248 4016 8276
rect 5810 8236 5816 8288
rect 5868 8276 5874 8288
rect 9858 8276 9864 8288
rect 5868 8248 9864 8276
rect 5868 8236 5874 8248
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10244 8276 10272 8316
rect 13170 8304 13176 8316
rect 13228 8304 13234 8356
rect 13357 8347 13415 8353
rect 13357 8313 13369 8347
rect 13403 8344 13415 8347
rect 13814 8344 13820 8356
rect 13403 8316 13820 8344
rect 13403 8313 13415 8316
rect 13357 8307 13415 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 13924 8344 13952 8384
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 15028 8412 15056 8443
rect 15654 8440 15660 8452
rect 15712 8440 15718 8492
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8480 15807 8483
rect 15930 8480 15936 8492
rect 15795 8452 15936 8480
rect 15795 8449 15807 8452
rect 15749 8443 15807 8449
rect 15930 8440 15936 8452
rect 15988 8440 15994 8492
rect 16114 8440 16120 8492
rect 16172 8440 16178 8492
rect 16298 8440 16304 8492
rect 16356 8440 16362 8492
rect 16500 8489 16528 8520
rect 27982 8508 27988 8520
rect 28040 8508 28046 8560
rect 32582 8508 32588 8560
rect 32640 8548 32646 8560
rect 33428 8548 33456 8579
rect 33962 8576 33968 8628
rect 34020 8616 34026 8628
rect 34885 8619 34943 8625
rect 34885 8616 34897 8619
rect 34020 8588 34897 8616
rect 34020 8576 34026 8588
rect 34885 8585 34897 8588
rect 34931 8585 34943 8619
rect 34885 8579 34943 8585
rect 35066 8576 35072 8628
rect 35124 8616 35130 8628
rect 35989 8619 36047 8625
rect 35989 8616 36001 8619
rect 35124 8588 36001 8616
rect 35124 8576 35130 8588
rect 35989 8585 36001 8588
rect 36035 8585 36047 8619
rect 35989 8579 36047 8585
rect 36446 8576 36452 8628
rect 36504 8616 36510 8628
rect 37461 8619 37519 8625
rect 37461 8616 37473 8619
rect 36504 8588 37473 8616
rect 36504 8576 36510 8588
rect 37461 8585 37473 8588
rect 37507 8585 37519 8619
rect 37461 8579 37519 8585
rect 37829 8619 37887 8625
rect 37829 8585 37841 8619
rect 37875 8585 37887 8619
rect 37829 8579 37887 8585
rect 32640 8520 33456 8548
rect 34072 8520 36584 8548
rect 32640 8508 32646 8520
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8449 16543 8483
rect 16485 8443 16543 8449
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8480 17279 8483
rect 17494 8480 17500 8492
rect 17267 8452 17500 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 17589 8483 17647 8489
rect 17589 8449 17601 8483
rect 17635 8480 17647 8483
rect 17635 8452 22094 8480
rect 17635 8449 17647 8452
rect 17589 8443 17647 8449
rect 22066 8412 22094 8452
rect 23014 8440 23020 8492
rect 23072 8480 23078 8492
rect 31757 8483 31815 8489
rect 31757 8480 31769 8483
rect 23072 8452 31769 8480
rect 23072 8440 23078 8452
rect 31757 8449 31769 8452
rect 31803 8449 31815 8483
rect 31757 8443 31815 8449
rect 32122 8440 32128 8492
rect 32180 8440 32186 8492
rect 32490 8440 32496 8492
rect 32548 8440 32554 8492
rect 32674 8440 32680 8492
rect 32732 8480 32738 8492
rect 32861 8483 32919 8489
rect 32861 8480 32873 8483
rect 32732 8452 32873 8480
rect 32732 8440 32738 8452
rect 32861 8449 32873 8452
rect 32907 8449 32919 8483
rect 32861 8443 32919 8449
rect 33229 8483 33287 8489
rect 33229 8449 33241 8483
rect 33275 8480 33287 8483
rect 33502 8480 33508 8492
rect 33275 8452 33508 8480
rect 33275 8449 33287 8452
rect 33229 8443 33287 8449
rect 33502 8440 33508 8452
rect 33560 8440 33566 8492
rect 33594 8440 33600 8492
rect 33652 8440 33658 8492
rect 33965 8483 34023 8489
rect 33965 8449 33977 8483
rect 34011 8449 34023 8483
rect 33965 8443 34023 8449
rect 26142 8412 26148 8424
rect 15028 8384 17908 8412
rect 22066 8384 26148 8412
rect 16114 8344 16120 8356
rect 13924 8316 16120 8344
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 17405 8347 17463 8353
rect 17405 8344 17417 8347
rect 16632 8316 17417 8344
rect 16632 8304 16638 8316
rect 17405 8313 17417 8316
rect 17451 8313 17463 8347
rect 17405 8307 17463 8313
rect 11054 8276 11060 8288
rect 10244 8248 11060 8276
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 17770 8276 17776 8288
rect 12676 8248 17776 8276
rect 12676 8236 12682 8248
rect 17770 8236 17776 8248
rect 17828 8236 17834 8288
rect 17880 8276 17908 8384
rect 26142 8372 26148 8384
rect 26200 8372 26206 8424
rect 26418 8372 26424 8424
rect 26476 8412 26482 8424
rect 33980 8412 34008 8443
rect 26476 8384 34008 8412
rect 26476 8372 26482 8384
rect 27706 8304 27712 8356
rect 27764 8344 27770 8356
rect 28350 8344 28356 8356
rect 27764 8316 28356 8344
rect 27764 8304 27770 8316
rect 28350 8304 28356 8316
rect 28408 8304 28414 8356
rect 32030 8304 32036 8356
rect 32088 8344 32094 8356
rect 32677 8347 32735 8353
rect 32677 8344 32689 8347
rect 32088 8316 32689 8344
rect 32088 8304 32094 8316
rect 32677 8313 32689 8316
rect 32723 8313 32735 8347
rect 32677 8307 32735 8313
rect 32858 8304 32864 8356
rect 32916 8344 32922 8356
rect 33781 8347 33839 8353
rect 33781 8344 33793 8347
rect 32916 8316 33793 8344
rect 32916 8304 32922 8316
rect 33781 8313 33793 8316
rect 33827 8313 33839 8347
rect 34072 8344 34100 8520
rect 34606 8440 34612 8492
rect 34664 8480 34670 8492
rect 34701 8483 34759 8489
rect 34701 8480 34713 8483
rect 34664 8452 34713 8480
rect 34664 8440 34670 8452
rect 34701 8449 34713 8452
rect 34747 8449 34759 8483
rect 34701 8443 34759 8449
rect 34882 8440 34888 8492
rect 34940 8480 34946 8492
rect 35069 8483 35127 8489
rect 35069 8480 35081 8483
rect 34940 8452 35081 8480
rect 34940 8440 34946 8452
rect 35069 8449 35081 8452
rect 35115 8449 35127 8483
rect 35069 8443 35127 8449
rect 35434 8440 35440 8492
rect 35492 8440 35498 8492
rect 35618 8440 35624 8492
rect 35676 8480 35682 8492
rect 35676 8452 35756 8480
rect 35676 8440 35682 8452
rect 34514 8372 34520 8424
rect 34572 8412 34578 8424
rect 35728 8412 35756 8452
rect 35802 8440 35808 8492
rect 35860 8440 35866 8492
rect 35986 8440 35992 8492
rect 36044 8480 36050 8492
rect 36556 8489 36584 8520
rect 36722 8508 36728 8560
rect 36780 8548 36786 8560
rect 37844 8548 37872 8579
rect 36780 8520 37872 8548
rect 36780 8508 36786 8520
rect 36173 8483 36231 8489
rect 36173 8480 36185 8483
rect 36044 8452 36185 8480
rect 36044 8440 36050 8452
rect 36173 8449 36185 8452
rect 36219 8449 36231 8483
rect 36173 8443 36231 8449
rect 36541 8483 36599 8489
rect 36541 8449 36553 8483
rect 36587 8449 36599 8483
rect 36541 8443 36599 8449
rect 37274 8440 37280 8492
rect 37332 8440 37338 8492
rect 37366 8440 37372 8492
rect 37424 8480 37430 8492
rect 37645 8483 37703 8489
rect 37645 8480 37657 8483
rect 37424 8452 37657 8480
rect 37424 8440 37430 8452
rect 37645 8449 37657 8452
rect 37691 8449 37703 8483
rect 37645 8443 37703 8449
rect 38194 8440 38200 8492
rect 38252 8440 38258 8492
rect 34572 8384 35664 8412
rect 35728 8384 36768 8412
rect 34572 8372 34578 8384
rect 33781 8307 33839 8313
rect 33888 8316 34100 8344
rect 29638 8276 29644 8288
rect 17880 8248 29644 8276
rect 29638 8236 29644 8248
rect 29696 8236 29702 8288
rect 32950 8236 32956 8288
rect 33008 8276 33014 8288
rect 33888 8276 33916 8316
rect 34146 8304 34152 8356
rect 34204 8304 34210 8356
rect 34238 8304 34244 8356
rect 34296 8344 34302 8356
rect 35636 8353 35664 8384
rect 35253 8347 35311 8353
rect 35253 8344 35265 8347
rect 34296 8316 35265 8344
rect 34296 8304 34302 8316
rect 35253 8313 35265 8316
rect 35299 8313 35311 8347
rect 35253 8307 35311 8313
rect 35621 8347 35679 8353
rect 35621 8313 35633 8347
rect 35667 8313 35679 8347
rect 35621 8307 35679 8313
rect 35710 8304 35716 8356
rect 35768 8344 35774 8356
rect 36740 8353 36768 8384
rect 36357 8347 36415 8353
rect 36357 8344 36369 8347
rect 35768 8316 36369 8344
rect 35768 8304 35774 8316
rect 36357 8313 36369 8316
rect 36403 8313 36415 8347
rect 36357 8307 36415 8313
rect 36725 8347 36783 8353
rect 36725 8313 36737 8347
rect 36771 8313 36783 8347
rect 36725 8307 36783 8313
rect 38378 8304 38384 8356
rect 38436 8304 38442 8356
rect 33008 8248 33916 8276
rect 33008 8236 33014 8248
rect 1104 8186 38824 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 38824 8186
rect 1104 8112 38824 8134
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 3237 8075 3295 8081
rect 3237 8072 3249 8075
rect 2924 8044 3249 8072
rect 2924 8032 2930 8044
rect 3237 8041 3249 8044
rect 3283 8041 3295 8075
rect 3237 8035 3295 8041
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 3881 8075 3939 8081
rect 3881 8072 3893 8075
rect 3660 8044 3893 8072
rect 3660 8032 3666 8044
rect 3881 8041 3893 8044
rect 3927 8041 3939 8075
rect 3881 8035 3939 8041
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 4212 8044 4353 8072
rect 4212 8032 4218 8044
rect 4341 8041 4353 8044
rect 4387 8041 4399 8075
rect 4341 8035 4399 8041
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 5316 8044 5457 8072
rect 5316 8032 5322 8044
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6273 8075 6331 8081
rect 6273 8072 6285 8075
rect 6144 8044 6285 8072
rect 6144 8032 6150 8044
rect 6273 8041 6285 8044
rect 6319 8041 6331 8075
rect 6273 8035 6331 8041
rect 6638 8032 6644 8084
rect 6696 8072 6702 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6696 8044 6837 8072
rect 6696 8032 6702 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 7524 8044 7665 8072
rect 7524 8032 7530 8044
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 7653 8035 7711 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8481 8075 8539 8081
rect 8481 8072 8493 8075
rect 8352 8044 8493 8072
rect 8352 8032 8358 8044
rect 8481 8041 8493 8044
rect 8527 8041 8539 8075
rect 8481 8035 8539 8041
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 8904 8044 9321 8072
rect 8904 8032 8910 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 9309 8035 9367 8041
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 9732 8044 9873 8072
rect 9732 8032 9738 8044
rect 9861 8041 9873 8044
rect 9907 8041 9919 8075
rect 9861 8035 9919 8041
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 10965 8075 11023 8081
rect 10965 8072 10977 8075
rect 10836 8044 10977 8072
rect 10836 8032 10842 8044
rect 10965 8041 10977 8044
rect 11011 8041 11023 8075
rect 10965 8035 11023 8041
rect 11330 8032 11336 8084
rect 11388 8072 11394 8084
rect 11517 8075 11575 8081
rect 11517 8072 11529 8075
rect 11388 8044 11529 8072
rect 11388 8032 11394 8044
rect 11517 8041 11529 8044
rect 11563 8041 11575 8075
rect 11517 8035 11575 8041
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 12069 8075 12127 8081
rect 12069 8072 12081 8075
rect 11940 8044 12081 8072
rect 11940 8032 11946 8044
rect 12069 8041 12081 8044
rect 12115 8041 12127 8075
rect 12069 8035 12127 8041
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13173 8075 13231 8081
rect 13173 8072 13185 8075
rect 13044 8044 13185 8072
rect 13044 8032 13050 8044
rect 13173 8041 13185 8044
rect 13219 8041 13231 8075
rect 13173 8035 13231 8041
rect 13538 8032 13544 8084
rect 13596 8072 13602 8084
rect 13725 8075 13783 8081
rect 13725 8072 13737 8075
rect 13596 8044 13737 8072
rect 13596 8032 13602 8044
rect 13725 8041 13737 8044
rect 13771 8041 13783 8075
rect 13725 8035 13783 8041
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14553 8075 14611 8081
rect 14553 8072 14565 8075
rect 14424 8044 14565 8072
rect 14424 8032 14430 8044
rect 14553 8041 14565 8044
rect 14599 8041 14611 8075
rect 14553 8035 14611 8041
rect 15378 8032 15384 8084
rect 15436 8032 15442 8084
rect 17770 8032 17776 8084
rect 17828 8072 17834 8084
rect 19058 8072 19064 8084
rect 17828 8044 19064 8072
rect 17828 8032 17834 8044
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 28994 8032 29000 8084
rect 29052 8072 29058 8084
rect 29914 8072 29920 8084
rect 29052 8044 29920 8072
rect 29052 8032 29058 8044
rect 29914 8032 29920 8044
rect 29972 8032 29978 8084
rect 33410 8032 33416 8084
rect 33468 8072 33474 8084
rect 33689 8075 33747 8081
rect 33689 8072 33701 8075
rect 33468 8044 33701 8072
rect 33468 8032 33474 8044
rect 33689 8041 33701 8044
rect 33735 8041 33747 8075
rect 33689 8035 33747 8041
rect 33778 8032 33784 8084
rect 33836 8072 33842 8084
rect 34057 8075 34115 8081
rect 34057 8072 34069 8075
rect 33836 8044 34069 8072
rect 33836 8032 33842 8044
rect 34057 8041 34069 8044
rect 34103 8041 34115 8075
rect 34057 8035 34115 8041
rect 34790 8032 34796 8084
rect 34848 8072 34854 8084
rect 35069 8075 35127 8081
rect 35069 8072 35081 8075
rect 34848 8044 35081 8072
rect 34848 8032 34854 8044
rect 35069 8041 35081 8044
rect 35115 8041 35127 8075
rect 35069 8035 35127 8041
rect 35894 8032 35900 8084
rect 35952 8072 35958 8084
rect 36173 8075 36231 8081
rect 36173 8072 36185 8075
rect 35952 8044 36185 8072
rect 35952 8032 35958 8044
rect 36173 8041 36185 8044
rect 36219 8041 36231 8075
rect 36173 8035 36231 8041
rect 36262 8032 36268 8084
rect 36320 8072 36326 8084
rect 36541 8075 36599 8081
rect 36541 8072 36553 8075
rect 36320 8044 36553 8072
rect 36320 8032 36326 8044
rect 36541 8041 36553 8044
rect 36587 8041 36599 8075
rect 36541 8035 36599 8041
rect 36906 8032 36912 8084
rect 36964 8032 36970 8084
rect 36998 8032 37004 8084
rect 37056 8072 37062 8084
rect 37277 8075 37335 8081
rect 37277 8072 37289 8075
rect 37056 8044 37289 8072
rect 37056 8032 37062 8044
rect 37277 8041 37289 8044
rect 37323 8041 37335 8075
rect 37277 8035 37335 8041
rect 37645 8075 37703 8081
rect 37645 8041 37657 8075
rect 37691 8072 37703 8075
rect 38654 8072 38660 8084
rect 37691 8044 38660 8072
rect 37691 8041 37703 8044
rect 37645 8035 37703 8041
rect 38654 8032 38660 8044
rect 38712 8032 38718 8084
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 14642 8004 14648 8016
rect 5684 7976 14648 8004
rect 5684 7964 5690 7976
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 6730 7936 6736 7948
rect 4540 7908 6736 7936
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3436 7800 3464 7831
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 4540 7877 4568 7908
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 8478 7936 8484 7948
rect 7024 7908 8484 7936
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7868 5687 7871
rect 5994 7868 6000 7880
rect 5675 7840 6000 7868
rect 5675 7837 5687 7840
rect 5629 7831 5687 7837
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7868 6515 7871
rect 6914 7868 6920 7880
rect 6503 7840 6920 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7024 7877 7052 7908
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 16758 7936 16764 7948
rect 8680 7908 16764 7936
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 8294 7868 8300 7880
rect 7883 7840 8300 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 8680 7877 8708 7908
rect 16758 7896 16764 7908
rect 16816 7896 16822 7948
rect 32766 7896 32772 7948
rect 32824 7936 32830 7948
rect 32824 7908 34928 7936
rect 32824 7896 32830 7908
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7837 8723 7871
rect 8665 7831 8723 7837
rect 9490 7828 9496 7880
rect 9548 7828 9554 7880
rect 10042 7828 10048 7880
rect 10100 7828 10106 7880
rect 11146 7828 11152 7880
rect 11204 7828 11210 7880
rect 11698 7828 11704 7880
rect 11756 7828 11762 7880
rect 12250 7828 12256 7880
rect 12308 7828 12314 7880
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 13722 7868 13728 7880
rect 13403 7840 13728 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7868 13967 7871
rect 14642 7868 14648 7880
rect 13955 7840 14648 7868
rect 13955 7837 13967 7840
rect 13909 7831 13967 7837
rect 14642 7828 14648 7840
rect 14700 7828 14706 7880
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7868 15623 7871
rect 30006 7868 30012 7880
rect 15611 7840 30012 7868
rect 15611 7837 15623 7840
rect 15565 7831 15623 7837
rect 6086 7800 6092 7812
rect 3436 7772 6092 7800
rect 6086 7760 6092 7772
rect 6144 7760 6150 7812
rect 6178 7760 6184 7812
rect 6236 7800 6242 7812
rect 11974 7800 11980 7812
rect 6236 7772 11980 7800
rect 6236 7760 6242 7772
rect 11974 7760 11980 7772
rect 12032 7760 12038 7812
rect 14752 7800 14780 7831
rect 30006 7828 30012 7840
rect 30064 7828 30070 7880
rect 32398 7828 32404 7880
rect 32456 7868 32462 7880
rect 34900 7877 34928 7908
rect 34974 7896 34980 7948
rect 35032 7936 35038 7948
rect 35032 7908 37872 7936
rect 35032 7896 35038 7908
rect 33505 7871 33563 7877
rect 33505 7868 33517 7871
rect 32456 7840 33517 7868
rect 32456 7828 32462 7840
rect 33505 7837 33517 7840
rect 33551 7837 33563 7871
rect 33505 7831 33563 7837
rect 33873 7871 33931 7877
rect 33873 7837 33885 7871
rect 33919 7837 33931 7871
rect 33873 7831 33931 7837
rect 34885 7871 34943 7877
rect 34885 7837 34897 7871
rect 34931 7837 34943 7871
rect 34885 7831 34943 7837
rect 18414 7800 18420 7812
rect 14752 7772 18420 7800
rect 18414 7760 18420 7772
rect 18472 7760 18478 7812
rect 22002 7760 22008 7812
rect 22060 7800 22066 7812
rect 33778 7800 33784 7812
rect 22060 7772 33784 7800
rect 22060 7760 22066 7772
rect 33778 7760 33784 7772
rect 33836 7760 33842 7812
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 13630 7732 13636 7744
rect 7064 7704 13636 7732
rect 7064 7692 7070 7704
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 15562 7692 15568 7744
rect 15620 7732 15626 7744
rect 23382 7732 23388 7744
rect 15620 7704 23388 7732
rect 15620 7692 15626 7704
rect 23382 7692 23388 7704
rect 23440 7692 23446 7744
rect 31754 7692 31760 7744
rect 31812 7732 31818 7744
rect 33888 7732 33916 7831
rect 35066 7828 35072 7880
rect 35124 7868 35130 7880
rect 35989 7871 36047 7877
rect 35989 7868 36001 7871
rect 35124 7840 36001 7868
rect 35124 7828 35130 7840
rect 35989 7837 36001 7840
rect 36035 7837 36047 7871
rect 35989 7831 36047 7837
rect 36354 7828 36360 7880
rect 36412 7828 36418 7880
rect 36722 7828 36728 7880
rect 36780 7828 36786 7880
rect 37090 7828 37096 7880
rect 37148 7828 37154 7880
rect 37458 7828 37464 7880
rect 37516 7828 37522 7880
rect 37844 7877 37872 7908
rect 37829 7871 37887 7877
rect 37829 7837 37841 7871
rect 37875 7837 37887 7871
rect 37829 7831 37887 7837
rect 38197 7871 38255 7877
rect 38197 7837 38209 7871
rect 38243 7837 38255 7871
rect 38197 7831 38255 7837
rect 35158 7760 35164 7812
rect 35216 7800 35222 7812
rect 38212 7800 38240 7831
rect 35216 7772 38240 7800
rect 35216 7760 35222 7772
rect 31812 7704 33916 7732
rect 31812 7692 31818 7704
rect 38010 7692 38016 7744
rect 38068 7692 38074 7744
rect 38378 7692 38384 7744
rect 38436 7692 38442 7744
rect 1104 7642 38824 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 38824 7642
rect 1104 7568 38824 7590
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 5169 7531 5227 7537
rect 5169 7528 5181 7531
rect 4120 7500 5181 7528
rect 4120 7488 4126 7500
rect 5169 7497 5181 7500
rect 5215 7497 5227 7531
rect 5169 7491 5227 7497
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5445 7531 5503 7537
rect 5445 7528 5457 7531
rect 5408 7500 5457 7528
rect 5408 7488 5414 7500
rect 5445 7497 5457 7500
rect 5491 7497 5503 7531
rect 5445 7491 5503 7497
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 5592 7500 5733 7528
rect 5592 7488 5598 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 5994 7488 6000 7540
rect 6052 7488 6058 7540
rect 6086 7488 6092 7540
rect 6144 7528 6150 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6144 7500 6837 7528
rect 6144 7488 6150 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 7101 7531 7159 7537
rect 7101 7528 7113 7531
rect 6972 7500 7113 7528
rect 6972 7488 6978 7500
rect 7101 7497 7113 7500
rect 7147 7497 7159 7531
rect 7101 7491 7159 7497
rect 7653 7531 7711 7537
rect 7653 7497 7665 7531
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 5810 7460 5816 7472
rect 5368 7432 5816 7460
rect 5368 7401 5396 7432
rect 5810 7420 5816 7432
rect 5868 7420 5874 7472
rect 6454 7420 6460 7472
rect 6512 7460 6518 7472
rect 7668 7460 7696 7491
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 14185 7531 14243 7537
rect 14185 7528 14197 7531
rect 10100 7500 14197 7528
rect 10100 7488 10106 7500
rect 14185 7497 14197 7500
rect 14231 7497 14243 7531
rect 14185 7491 14243 7497
rect 14826 7488 14832 7540
rect 14884 7528 14890 7540
rect 14921 7531 14979 7537
rect 14921 7528 14933 7531
rect 14884 7500 14933 7528
rect 14884 7488 14890 7500
rect 14921 7497 14933 7500
rect 14967 7497 14979 7531
rect 14921 7491 14979 7497
rect 15381 7531 15439 7537
rect 15381 7497 15393 7531
rect 15427 7497 15439 7531
rect 15381 7491 15439 7497
rect 15749 7531 15807 7537
rect 15749 7497 15761 7531
rect 15795 7528 15807 7531
rect 15838 7528 15844 7540
rect 15795 7500 15844 7528
rect 15795 7497 15807 7500
rect 15749 7491 15807 7497
rect 6512 7432 7696 7460
rect 6512 7420 6518 7432
rect 9490 7420 9496 7472
rect 9548 7460 9554 7472
rect 15396 7460 15424 7491
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 16758 7488 16764 7540
rect 16816 7488 16822 7540
rect 17034 7488 17040 7540
rect 17092 7488 17098 7540
rect 19889 7531 19947 7537
rect 19889 7497 19901 7531
rect 19935 7528 19947 7531
rect 20990 7528 20996 7540
rect 19935 7500 20996 7528
rect 19935 7497 19947 7500
rect 19889 7491 19947 7497
rect 20990 7488 20996 7500
rect 21048 7488 21054 7540
rect 22278 7488 22284 7540
rect 22336 7488 22342 7540
rect 22462 7488 22468 7540
rect 22520 7488 22526 7540
rect 22833 7531 22891 7537
rect 22833 7497 22845 7531
rect 22879 7528 22891 7531
rect 22879 7500 27292 7528
rect 22879 7497 22891 7500
rect 22833 7491 22891 7497
rect 16666 7460 16672 7472
rect 9548 7432 15424 7460
rect 15488 7432 16672 7460
rect 9548 7420 9554 7432
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 5920 7324 5948 7355
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 6914 7392 6920 7404
rect 6779 7364 6920 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 10134 7392 10140 7404
rect 7883 7364 10140 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 7300 7324 7328 7355
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7392 13047 7395
rect 13265 7395 13323 7401
rect 13265 7392 13277 7395
rect 13035 7364 13277 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13265 7361 13277 7364
rect 13311 7392 13323 7395
rect 13722 7392 13728 7404
rect 13311 7364 13728 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 12618 7324 12624 7336
rect 5920 7296 7236 7324
rect 7300 7296 12624 7324
rect 6362 7216 6368 7268
rect 6420 7256 6426 7268
rect 6549 7259 6607 7265
rect 6549 7256 6561 7259
rect 6420 7228 6561 7256
rect 6420 7216 6426 7228
rect 6549 7225 6561 7228
rect 6595 7225 6607 7259
rect 7208 7256 7236 7296
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 14108 7324 14136 7355
rect 14366 7352 14372 7404
rect 14424 7352 14430 7404
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7392 14703 7395
rect 14734 7392 14740 7404
rect 14691 7364 14740 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15488 7392 15516 7432
rect 16666 7420 16672 7432
rect 16724 7420 16730 7472
rect 19518 7460 19524 7472
rect 16960 7432 19524 7460
rect 15151 7364 15516 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 15562 7352 15568 7404
rect 15620 7352 15626 7404
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7392 15991 7395
rect 16482 7392 16488 7404
rect 15979 7364 16488 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16960 7401 16988 7432
rect 19518 7420 19524 7432
rect 19576 7420 19582 7472
rect 26786 7460 26792 7472
rect 20456 7432 20944 7460
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17218 7352 17224 7404
rect 17276 7352 17282 7404
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7392 18843 7395
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 18831 7364 18889 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 18877 7361 18889 7364
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 19702 7352 19708 7404
rect 19760 7352 19766 7404
rect 19978 7352 19984 7404
rect 20036 7352 20042 7404
rect 20346 7352 20352 7404
rect 20404 7392 20410 7404
rect 20456 7392 20484 7432
rect 20916 7401 20944 7432
rect 21008 7432 26792 7460
rect 20404 7364 20484 7392
rect 20533 7395 20591 7401
rect 20404 7352 20410 7364
rect 20533 7361 20545 7395
rect 20579 7392 20591 7395
rect 20625 7395 20683 7401
rect 20625 7392 20637 7395
rect 20579 7364 20637 7392
rect 20579 7361 20591 7364
rect 20533 7355 20591 7361
rect 20625 7361 20637 7364
rect 20671 7361 20683 7395
rect 20625 7355 20683 7361
rect 20901 7395 20959 7401
rect 20901 7361 20913 7395
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 20714 7324 20720 7336
rect 14108 7296 20720 7324
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 21008 7324 21036 7432
rect 26786 7420 26792 7432
rect 26844 7420 26850 7472
rect 27264 7460 27292 7500
rect 28810 7488 28816 7540
rect 28868 7488 28874 7540
rect 37458 7528 37464 7540
rect 30116 7500 37464 7528
rect 30116 7460 30144 7500
rect 37458 7488 37464 7500
rect 37516 7488 37522 7540
rect 37642 7488 37648 7540
rect 37700 7488 37706 7540
rect 38013 7531 38071 7537
rect 38013 7497 38025 7531
rect 38059 7528 38071 7531
rect 38286 7528 38292 7540
rect 38059 7500 38292 7528
rect 38059 7497 38071 7500
rect 38013 7491 38071 7497
rect 38286 7488 38292 7500
rect 38344 7488 38350 7540
rect 27264 7432 30144 7460
rect 33778 7420 33784 7472
rect 33836 7460 33842 7472
rect 33836 7432 37872 7460
rect 33836 7420 33842 7432
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7392 21327 7395
rect 21358 7392 21364 7404
rect 21315 7364 21364 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 21358 7352 21364 7364
rect 21416 7392 21422 7404
rect 21545 7395 21603 7401
rect 21545 7392 21557 7395
rect 21416 7364 21557 7392
rect 21416 7352 21422 7364
rect 21545 7361 21557 7364
rect 21591 7361 21603 7395
rect 21545 7355 21603 7361
rect 21818 7352 21824 7404
rect 21876 7352 21882 7404
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7392 22615 7395
rect 22649 7395 22707 7401
rect 22649 7392 22661 7395
rect 22603 7364 22661 7392
rect 22603 7361 22615 7364
rect 22557 7355 22615 7361
rect 22649 7361 22661 7364
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 22922 7352 22928 7404
rect 22980 7392 22986 7404
rect 23201 7395 23259 7401
rect 23201 7392 23213 7395
rect 22980 7364 23213 7392
rect 22980 7352 22986 7364
rect 23201 7361 23213 7364
rect 23247 7361 23259 7395
rect 23201 7355 23259 7361
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7392 24455 7395
rect 25866 7392 25872 7404
rect 24443 7364 25872 7392
rect 24443 7361 24455 7364
rect 24397 7355 24455 7361
rect 25866 7352 25872 7364
rect 25924 7352 25930 7404
rect 27890 7352 27896 7404
rect 27948 7392 27954 7404
rect 28997 7395 29055 7401
rect 28997 7392 29009 7395
rect 27948 7364 29009 7392
rect 27948 7352 27954 7364
rect 28997 7361 29009 7364
rect 29043 7361 29055 7395
rect 28997 7355 29055 7361
rect 29454 7352 29460 7404
rect 29512 7352 29518 7404
rect 29730 7352 29736 7404
rect 29788 7352 29794 7404
rect 29914 7352 29920 7404
rect 29972 7392 29978 7404
rect 30009 7395 30067 7401
rect 30009 7392 30021 7395
rect 29972 7364 30021 7392
rect 29972 7352 29978 7364
rect 30009 7361 30021 7364
rect 30055 7361 30067 7395
rect 30009 7355 30067 7361
rect 30282 7352 30288 7404
rect 30340 7352 30346 7404
rect 34238 7352 34244 7404
rect 34296 7392 34302 7404
rect 37844 7401 37872 7432
rect 36817 7395 36875 7401
rect 36817 7392 36829 7395
rect 34296 7364 36829 7392
rect 34296 7352 34302 7364
rect 36817 7361 36829 7364
rect 36863 7361 36875 7395
rect 36817 7355 36875 7361
rect 37461 7395 37519 7401
rect 37461 7361 37473 7395
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 37829 7395 37887 7401
rect 37829 7361 37841 7395
rect 37875 7361 37887 7395
rect 37829 7355 37887 7361
rect 38197 7395 38255 7401
rect 38197 7361 38209 7395
rect 38243 7361 38255 7395
rect 38197 7355 38255 7361
rect 37476 7324 37504 7355
rect 20824 7296 21036 7324
rect 21100 7296 37504 7324
rect 7834 7256 7840 7268
rect 7208 7228 7840 7256
rect 6549 7219 6607 7225
rect 7834 7216 7840 7228
rect 7892 7216 7898 7268
rect 11238 7216 11244 7268
rect 11296 7256 11302 7268
rect 13081 7259 13139 7265
rect 13081 7256 13093 7259
rect 11296 7228 13093 7256
rect 11296 7216 11302 7228
rect 13081 7225 13093 7228
rect 13127 7225 13139 7259
rect 13081 7219 13139 7225
rect 13446 7216 13452 7268
rect 13504 7256 13510 7268
rect 14461 7259 14519 7265
rect 14461 7256 14473 7259
rect 13504 7228 14473 7256
rect 13504 7216 13510 7228
rect 14461 7225 14473 7228
rect 14507 7225 14519 7259
rect 16390 7256 16396 7268
rect 14461 7219 14519 7225
rect 14568 7228 16396 7256
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7374 7188 7380 7200
rect 6972 7160 7380 7188
rect 6972 7148 6978 7160
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 13909 7191 13967 7197
rect 13909 7188 13921 7191
rect 11112 7160 13921 7188
rect 11112 7148 11118 7160
rect 13909 7157 13921 7160
rect 13955 7157 13967 7191
rect 13909 7151 13967 7157
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 14568 7188 14596 7228
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 19334 7216 19340 7268
rect 19392 7256 19398 7268
rect 20824 7265 20852 7296
rect 21100 7265 21128 7296
rect 20441 7259 20499 7265
rect 20441 7256 20453 7259
rect 19392 7228 20453 7256
rect 19392 7216 19398 7228
rect 20441 7225 20453 7228
rect 20487 7225 20499 7259
rect 20441 7219 20499 7225
rect 20809 7259 20867 7265
rect 20809 7225 20821 7259
rect 20855 7225 20867 7259
rect 20809 7219 20867 7225
rect 21085 7259 21143 7265
rect 21085 7225 21097 7259
rect 21131 7225 21143 7259
rect 23382 7256 23388 7268
rect 21085 7219 21143 7225
rect 21192 7228 23388 7256
rect 14424 7160 14596 7188
rect 14424 7148 14430 7160
rect 14642 7148 14648 7200
rect 14700 7188 14706 7200
rect 17678 7188 17684 7200
rect 14700 7160 17684 7188
rect 14700 7148 14706 7160
rect 17678 7148 17684 7160
rect 17736 7148 17742 7200
rect 18690 7148 18696 7200
rect 18748 7148 18754 7200
rect 19058 7148 19064 7200
rect 19116 7148 19122 7200
rect 20165 7191 20223 7197
rect 20165 7157 20177 7191
rect 20211 7188 20223 7191
rect 21192 7188 21220 7228
rect 23382 7216 23388 7228
rect 23440 7216 23446 7268
rect 24210 7216 24216 7268
rect 24268 7216 24274 7268
rect 26786 7216 26792 7268
rect 26844 7256 26850 7268
rect 34974 7256 34980 7268
rect 26844 7228 34980 7256
rect 26844 7216 26850 7228
rect 34974 7216 34980 7228
rect 35032 7216 35038 7268
rect 36998 7216 37004 7268
rect 37056 7216 37062 7268
rect 20211 7160 21220 7188
rect 20211 7157 20223 7160
rect 20165 7151 20223 7157
rect 21450 7148 21456 7200
rect 21508 7148 21514 7200
rect 22002 7148 22008 7200
rect 22060 7148 22066 7200
rect 23109 7191 23167 7197
rect 23109 7157 23121 7191
rect 23155 7188 23167 7191
rect 24762 7188 24768 7200
rect 23155 7160 24768 7188
rect 23155 7157 23167 7160
rect 23109 7151 23167 7157
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 28902 7148 28908 7200
rect 28960 7188 28966 7200
rect 29273 7191 29331 7197
rect 29273 7188 29285 7191
rect 28960 7160 29285 7188
rect 28960 7148 28966 7160
rect 29273 7157 29285 7160
rect 29319 7157 29331 7191
rect 29273 7151 29331 7157
rect 29362 7148 29368 7200
rect 29420 7188 29426 7200
rect 29549 7191 29607 7197
rect 29549 7188 29561 7191
rect 29420 7160 29561 7188
rect 29420 7148 29426 7160
rect 29549 7157 29561 7160
rect 29595 7157 29607 7191
rect 29549 7151 29607 7157
rect 29638 7148 29644 7200
rect 29696 7188 29702 7200
rect 29825 7191 29883 7197
rect 29825 7188 29837 7191
rect 29696 7160 29837 7188
rect 29696 7148 29702 7160
rect 29825 7157 29837 7160
rect 29871 7157 29883 7191
rect 29825 7151 29883 7157
rect 30006 7148 30012 7200
rect 30064 7188 30070 7200
rect 30101 7191 30159 7197
rect 30101 7188 30113 7191
rect 30064 7160 30113 7188
rect 30064 7148 30070 7160
rect 30101 7157 30113 7160
rect 30147 7157 30159 7191
rect 30101 7151 30159 7157
rect 34698 7148 34704 7200
rect 34756 7188 34762 7200
rect 38212 7188 38240 7355
rect 34756 7160 38240 7188
rect 34756 7148 34762 7160
rect 38378 7148 38384 7200
rect 38436 7148 38442 7200
rect 1104 7098 38824 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 38824 7098
rect 1104 7024 38824 7046
rect 8294 6944 8300 6996
rect 8352 6944 8358 6996
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 9953 6987 10011 6993
rect 9953 6984 9965 6987
rect 8536 6956 9965 6984
rect 8536 6944 8542 6956
rect 9953 6953 9965 6956
rect 9999 6953 10011 6987
rect 9953 6947 10011 6953
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 12308 6956 13645 6984
rect 12308 6944 12314 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 20806 6984 20812 6996
rect 13780 6956 20812 6984
rect 13780 6944 13786 6956
rect 20806 6944 20812 6956
rect 20864 6944 20870 6996
rect 36722 6984 36728 6996
rect 22066 6956 36728 6984
rect 9585 6919 9643 6925
rect 9585 6916 9597 6919
rect 8404 6888 9597 6916
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 8404 6848 8432 6888
rect 9585 6885 9597 6888
rect 9631 6885 9643 6919
rect 9585 6879 9643 6885
rect 13081 6919 13139 6925
rect 13081 6885 13093 6919
rect 13127 6885 13139 6919
rect 13081 6879 13139 6885
rect 14369 6919 14427 6925
rect 14369 6885 14381 6919
rect 14415 6885 14427 6919
rect 14369 6879 14427 6885
rect 19705 6919 19763 6925
rect 19705 6885 19717 6919
rect 19751 6885 19763 6919
rect 19705 6879 19763 6885
rect 11054 6848 11060 6860
rect 7340 6820 8432 6848
rect 8496 6820 11060 6848
rect 7340 6808 7346 6820
rect 6454 6740 6460 6792
rect 6512 6740 6518 6792
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 7834 6780 7840 6792
rect 7791 6752 7840 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 7834 6740 7840 6752
rect 7892 6780 7898 6792
rect 8496 6789 8524 6820
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 13096 6848 13124 6879
rect 11204 6820 13124 6848
rect 11204 6808 11210 6820
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 14384 6848 14412 6879
rect 13228 6820 14412 6848
rect 19720 6848 19748 6879
rect 21450 6876 21456 6928
rect 21508 6916 21514 6928
rect 22066 6916 22094 6956
rect 36722 6944 36728 6956
rect 36780 6944 36786 6996
rect 25685 6919 25743 6925
rect 25685 6916 25697 6919
rect 21508 6888 22094 6916
rect 25424 6888 25697 6916
rect 21508 6876 21514 6888
rect 22094 6848 22100 6860
rect 19720 6820 22100 6848
rect 13228 6808 13234 6820
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 22186 6808 22192 6860
rect 22244 6808 22250 6860
rect 22738 6808 22744 6860
rect 22796 6808 22802 6860
rect 23842 6808 23848 6860
rect 23900 6848 23906 6860
rect 25424 6848 25452 6888
rect 25685 6885 25697 6888
rect 25731 6885 25743 6919
rect 25685 6879 25743 6885
rect 25961 6919 26019 6925
rect 25961 6885 25973 6919
rect 26007 6916 26019 6919
rect 26142 6916 26148 6928
rect 26007 6888 26148 6916
rect 26007 6885 26019 6888
rect 25961 6879 26019 6885
rect 26142 6876 26148 6888
rect 26200 6876 26206 6928
rect 26881 6919 26939 6925
rect 26881 6885 26893 6919
rect 26927 6885 26939 6919
rect 26881 6879 26939 6885
rect 23900 6820 25452 6848
rect 23900 6808 23906 6820
rect 25774 6808 25780 6860
rect 25832 6848 25838 6860
rect 25832 6820 26004 6848
rect 25832 6808 25838 6820
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7892 6752 8033 6780
rect 7892 6740 7898 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9263 6752 9505 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 6730 6672 6736 6724
rect 6788 6712 6794 6724
rect 6788 6684 7972 6712
rect 6788 6672 6794 6684
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 6273 6647 6331 6653
rect 6273 6644 6285 6647
rect 5500 6616 6285 6644
rect 5500 6604 5506 6616
rect 6273 6613 6285 6616
rect 6319 6613 6331 6647
rect 6273 6607 6331 6613
rect 7558 6604 7564 6656
rect 7616 6604 7622 6656
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7800 6616 7849 6644
rect 7800 6604 7806 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7944 6644 7972 6684
rect 8573 6647 8631 6653
rect 8573 6644 8585 6647
rect 7944 6616 8585 6644
rect 7837 6607 7895 6613
rect 8573 6613 8585 6616
rect 8619 6613 8631 6647
rect 8573 6607 8631 6613
rect 9309 6647 9367 6653
rect 9309 6613 9321 6647
rect 9355 6644 9367 6647
rect 9398 6644 9404 6656
rect 9355 6616 9404 6644
rect 9355 6613 9367 6616
rect 9309 6607 9367 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9508 6644 9536 6743
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6780 10195 6783
rect 10318 6780 10324 6792
rect 10183 6752 10324 6780
rect 10183 6749 10195 6752
rect 10137 6743 10195 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10428 6712 10456 6743
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 10652 6752 12940 6780
rect 10652 6740 10658 6752
rect 12710 6712 12716 6724
rect 9876 6684 10364 6712
rect 10428 6684 12716 6712
rect 9876 6644 9904 6684
rect 9508 6616 9904 6644
rect 10226 6604 10232 6656
rect 10284 6604 10290 6656
rect 10336 6644 10364 6684
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 12912 6712 12940 6752
rect 12986 6740 12992 6792
rect 13044 6740 13050 6792
rect 13262 6740 13268 6792
rect 13320 6740 13326 6792
rect 13538 6740 13544 6792
rect 13596 6740 13602 6792
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 13832 6712 13860 6743
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 17862 6780 17868 6792
rect 14599 6752 17868 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19521 6783 19579 6789
rect 19521 6780 19533 6783
rect 19475 6752 19533 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19521 6749 19533 6752
rect 19567 6749 19579 6783
rect 19521 6743 19579 6749
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6780 20315 6783
rect 20349 6783 20407 6789
rect 20349 6780 20361 6783
rect 20303 6752 20361 6780
rect 20303 6749 20315 6752
rect 20257 6743 20315 6749
rect 20349 6749 20361 6752
rect 20395 6749 20407 6783
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20349 6743 20407 6749
rect 20456 6752 21005 6780
rect 14458 6712 14464 6724
rect 12912 6684 13400 6712
rect 13832 6684 14464 6712
rect 11422 6644 11428 6656
rect 10336 6616 11428 6644
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 13372 6653 13400 6684
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 17972 6712 18000 6743
rect 17788 6684 18000 6712
rect 17788 6656 17816 6684
rect 19242 6672 19248 6724
rect 19300 6712 19306 6724
rect 20165 6715 20223 6721
rect 20165 6712 20177 6715
rect 19300 6684 20177 6712
rect 19300 6672 19306 6684
rect 20165 6681 20177 6684
rect 20211 6681 20223 6715
rect 20165 6675 20223 6681
rect 12805 6647 12863 6653
rect 12805 6644 12817 6647
rect 11848 6616 12817 6644
rect 11848 6604 11854 6616
rect 12805 6613 12817 6616
rect 12851 6613 12863 6647
rect 12805 6607 12863 6613
rect 13357 6647 13415 6653
rect 13357 6613 13369 6647
rect 13403 6613 13415 6647
rect 13357 6607 13415 6613
rect 14093 6647 14151 6653
rect 14093 6613 14105 6647
rect 14139 6644 14151 6647
rect 14182 6644 14188 6656
rect 14139 6616 14188 6644
rect 14139 6613 14151 6616
rect 14093 6607 14151 6613
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 17770 6604 17776 6656
rect 17828 6604 17834 6656
rect 18138 6604 18144 6656
rect 18196 6604 18202 6656
rect 19334 6604 19340 6656
rect 19392 6604 19398 6656
rect 19518 6604 19524 6656
rect 19576 6644 19582 6656
rect 20456 6644 20484 6752
rect 20993 6749 21005 6752
rect 21039 6780 21051 6783
rect 21177 6783 21235 6789
rect 21177 6780 21189 6783
rect 21039 6752 21189 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21177 6749 21189 6752
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 22281 6783 22339 6789
rect 22281 6749 22293 6783
rect 22327 6780 22339 6783
rect 22373 6783 22431 6789
rect 22373 6780 22385 6783
rect 22327 6752 22385 6780
rect 22327 6749 22339 6752
rect 22281 6743 22339 6749
rect 22373 6749 22385 6752
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6780 22891 6783
rect 22925 6783 22983 6789
rect 22925 6780 22937 6783
rect 22879 6752 22937 6780
rect 22879 6749 22891 6752
rect 22833 6743 22891 6749
rect 22925 6749 22937 6752
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 25590 6740 25596 6792
rect 25648 6740 25654 6792
rect 25682 6740 25688 6792
rect 25740 6780 25746 6792
rect 25869 6783 25927 6789
rect 25869 6780 25881 6783
rect 25740 6752 25881 6780
rect 25740 6740 25746 6752
rect 25869 6749 25881 6752
rect 25915 6749 25927 6783
rect 25976 6780 26004 6820
rect 26326 6808 26332 6860
rect 26384 6848 26390 6860
rect 26896 6848 26924 6879
rect 28258 6876 28264 6928
rect 28316 6916 28322 6928
rect 28316 6888 28994 6916
rect 28316 6876 28322 6888
rect 26384 6820 26924 6848
rect 28966 6848 28994 6888
rect 29822 6848 29828 6860
rect 28966 6820 29828 6848
rect 26384 6808 26390 6820
rect 29822 6808 29828 6820
rect 29880 6808 29886 6860
rect 34974 6808 34980 6860
rect 35032 6848 35038 6860
rect 35032 6820 38240 6848
rect 35032 6808 35038 6820
rect 26145 6783 26203 6789
rect 26145 6780 26157 6783
rect 25976 6752 26157 6780
rect 25869 6743 25927 6749
rect 26145 6749 26157 6752
rect 26191 6749 26203 6783
rect 26145 6743 26203 6749
rect 26421 6783 26479 6789
rect 26421 6749 26433 6783
rect 26467 6780 26479 6783
rect 26878 6780 26884 6792
rect 26467 6752 26884 6780
rect 26467 6749 26479 6752
rect 26421 6743 26479 6749
rect 26878 6740 26884 6752
rect 26936 6740 26942 6792
rect 27065 6783 27123 6789
rect 27065 6749 27077 6783
rect 27111 6780 27123 6783
rect 27246 6780 27252 6792
rect 27111 6752 27252 6780
rect 27111 6749 27123 6752
rect 27065 6743 27123 6749
rect 27246 6740 27252 6752
rect 27304 6740 27310 6792
rect 27341 6783 27399 6789
rect 27341 6749 27353 6783
rect 27387 6749 27399 6783
rect 27341 6743 27399 6749
rect 26050 6712 26056 6724
rect 20548 6684 26056 6712
rect 20548 6653 20576 6684
rect 26050 6672 26056 6684
rect 26108 6672 26114 6724
rect 27356 6712 27384 6743
rect 27614 6740 27620 6792
rect 27672 6740 27678 6792
rect 28077 6783 28135 6789
rect 28077 6749 28089 6783
rect 28123 6776 28135 6783
rect 28123 6749 28304 6776
rect 28077 6748 28304 6749
rect 28077 6743 28135 6748
rect 28276 6712 28304 6748
rect 28350 6740 28356 6792
rect 28408 6740 28414 6792
rect 28721 6783 28779 6789
rect 28721 6749 28733 6783
rect 28767 6780 28779 6783
rect 29270 6780 29276 6792
rect 28767 6752 29276 6780
rect 28767 6749 28779 6752
rect 28721 6743 28779 6749
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 37458 6740 37464 6792
rect 37516 6740 37522 6792
rect 37550 6740 37556 6792
rect 37608 6780 37614 6792
rect 38212 6789 38240 6820
rect 37829 6783 37887 6789
rect 37829 6780 37841 6783
rect 37608 6752 37841 6780
rect 37608 6740 37614 6752
rect 37829 6749 37841 6752
rect 37875 6749 37887 6783
rect 37829 6743 37887 6749
rect 38197 6783 38255 6789
rect 38197 6749 38209 6783
rect 38243 6749 38255 6783
rect 38197 6743 38255 6749
rect 29546 6712 29552 6724
rect 27356 6684 28120 6712
rect 28276 6684 29552 6712
rect 28092 6656 28120 6684
rect 29546 6672 29552 6684
rect 29604 6672 29610 6724
rect 38562 6712 38568 6724
rect 38028 6684 38568 6712
rect 19576 6616 20484 6644
rect 20533 6647 20591 6653
rect 19576 6604 19582 6616
rect 20533 6613 20545 6647
rect 20579 6613 20591 6647
rect 20533 6607 20591 6613
rect 21361 6647 21419 6653
rect 21361 6613 21373 6647
rect 21407 6644 21419 6647
rect 22094 6644 22100 6656
rect 21407 6616 22100 6644
rect 21407 6613 21419 6616
rect 21361 6607 21419 6613
rect 22094 6604 22100 6616
rect 22152 6604 22158 6656
rect 22554 6604 22560 6656
rect 22612 6604 22618 6656
rect 23106 6604 23112 6656
rect 23164 6604 23170 6656
rect 25406 6604 25412 6656
rect 25464 6604 25470 6656
rect 25498 6604 25504 6656
rect 25556 6644 25562 6656
rect 26237 6647 26295 6653
rect 26237 6644 26249 6647
rect 25556 6616 26249 6644
rect 25556 6604 25562 6616
rect 26237 6613 26249 6616
rect 26283 6613 26295 6647
rect 26237 6607 26295 6613
rect 26602 6604 26608 6656
rect 26660 6644 26666 6656
rect 27157 6647 27215 6653
rect 27157 6644 27169 6647
rect 26660 6616 27169 6644
rect 26660 6604 26666 6616
rect 27157 6613 27169 6616
rect 27203 6613 27215 6647
rect 27157 6607 27215 6613
rect 27430 6604 27436 6656
rect 27488 6604 27494 6656
rect 27890 6604 27896 6656
rect 27948 6604 27954 6656
rect 28074 6604 28080 6656
rect 28132 6604 28138 6656
rect 28169 6647 28227 6653
rect 28169 6613 28181 6647
rect 28215 6644 28227 6647
rect 28350 6644 28356 6656
rect 28215 6616 28356 6644
rect 28215 6613 28227 6616
rect 28169 6607 28227 6613
rect 28350 6604 28356 6616
rect 28408 6604 28414 6656
rect 28534 6604 28540 6656
rect 28592 6604 28598 6656
rect 37642 6604 37648 6656
rect 37700 6604 37706 6656
rect 38028 6653 38056 6684
rect 38562 6672 38568 6684
rect 38620 6672 38626 6724
rect 38013 6647 38071 6653
rect 38013 6613 38025 6647
rect 38059 6613 38071 6647
rect 38013 6607 38071 6613
rect 38381 6647 38439 6653
rect 38381 6613 38393 6647
rect 38427 6644 38439 6647
rect 38470 6644 38476 6656
rect 38427 6616 38476 6644
rect 38427 6613 38439 6616
rect 38381 6607 38439 6613
rect 38470 6604 38476 6616
rect 38528 6604 38534 6656
rect 1104 6554 38824 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 38824 6554
rect 1104 6480 38824 6502
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 9398 6440 9404 6452
rect 7248 6412 9404 6440
rect 7248 6400 7254 6412
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 9582 6400 9588 6452
rect 9640 6440 9646 6452
rect 10229 6443 10287 6449
rect 10229 6440 10241 6443
rect 9640 6412 10241 6440
rect 9640 6400 9646 6412
rect 10229 6409 10241 6412
rect 10275 6409 10287 6443
rect 10229 6403 10287 6409
rect 10318 6400 10324 6452
rect 10376 6440 10382 6452
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 10376 6412 10609 6440
rect 10376 6400 10382 6412
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 11756 6412 13185 6440
rect 11756 6400 11762 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 16850 6440 16856 6452
rect 13173 6403 13231 6409
rect 13372 6412 16856 6440
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 9950 6304 9956 6316
rect 8812 6276 9956 6304
rect 8812 6264 8818 6276
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 10410 6313 10416 6316
rect 10405 6267 10416 6313
rect 10468 6304 10474 6316
rect 10781 6307 10839 6313
rect 10468 6276 10505 6304
rect 10410 6264 10416 6267
rect 10468 6264 10474 6276
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 10962 6304 10968 6316
rect 10827 6276 10968 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 13372 6313 13400 6412
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17083 6412 17264 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17236 6372 17264 6412
rect 17310 6400 17316 6452
rect 17368 6440 17374 6452
rect 22094 6440 22100 6452
rect 17368 6412 22100 6440
rect 17368 6400 17374 6412
rect 22094 6400 22100 6412
rect 22152 6400 22158 6452
rect 22186 6400 22192 6452
rect 22244 6440 22250 6452
rect 22244 6412 28028 6440
rect 22244 6400 22250 6412
rect 18230 6372 18236 6384
rect 17236 6344 18236 6372
rect 18230 6332 18236 6344
rect 18288 6332 18294 6384
rect 18414 6332 18420 6384
rect 18472 6372 18478 6384
rect 27890 6372 27896 6384
rect 18472 6344 27896 6372
rect 18472 6332 18478 6344
rect 27890 6332 27896 6344
rect 27948 6332 27954 6384
rect 28000 6372 28028 6412
rect 28442 6400 28448 6452
rect 28500 6400 28506 6452
rect 29457 6443 29515 6449
rect 29457 6409 29469 6443
rect 29503 6440 29515 6443
rect 35986 6440 35992 6452
rect 29503 6412 35992 6440
rect 29503 6409 29515 6412
rect 29457 6403 29515 6409
rect 35986 6400 35992 6412
rect 36044 6400 36050 6452
rect 38378 6400 38384 6452
rect 38436 6400 38442 6452
rect 37458 6372 37464 6384
rect 28000 6344 37464 6372
rect 37458 6332 37464 6344
rect 37516 6332 37522 6384
rect 37734 6332 37740 6384
rect 37792 6372 37798 6384
rect 37792 6344 38240 6372
rect 37792 6332 37798 6344
rect 13357 6307 13415 6313
rect 13357 6273 13369 6307
rect 13403 6273 13415 6307
rect 13357 6267 13415 6273
rect 16758 6264 16764 6316
rect 16816 6304 16822 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16816 6276 16865 6304
rect 16816 6264 16822 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 16960 6276 17172 6304
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 10226 6236 10232 6248
rect 7156 6208 10232 6236
rect 7156 6196 7162 6208
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 16960 6236 16988 6276
rect 12768 6208 16988 6236
rect 17144 6236 17172 6276
rect 17218 6264 17224 6316
rect 17276 6304 17282 6316
rect 21542 6304 21548 6316
rect 17276 6276 21548 6304
rect 17276 6264 17282 6276
rect 21542 6264 21548 6276
rect 21600 6264 21606 6316
rect 21634 6264 21640 6316
rect 21692 6304 21698 6316
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 21692 6276 22293 6304
rect 21692 6264 21698 6276
rect 22281 6273 22293 6276
rect 22327 6273 22339 6307
rect 23750 6304 23756 6316
rect 22281 6267 22339 6273
rect 22480 6276 23756 6304
rect 19794 6236 19800 6248
rect 17144 6208 19800 6236
rect 12768 6196 12774 6208
rect 19794 6196 19800 6208
rect 19852 6196 19858 6248
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 22480 6236 22508 6276
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 25498 6264 25504 6316
rect 25556 6304 25562 6316
rect 28261 6307 28319 6313
rect 28261 6304 28273 6307
rect 25556 6276 28273 6304
rect 25556 6264 25562 6276
rect 28261 6273 28273 6276
rect 28307 6273 28319 6307
rect 28261 6267 28319 6273
rect 29270 6264 29276 6316
rect 29328 6264 29334 6316
rect 35158 6304 35164 6316
rect 29380 6276 35164 6304
rect 22152 6208 22508 6236
rect 22152 6196 22158 6208
rect 22554 6196 22560 6248
rect 22612 6236 22618 6248
rect 29380 6236 29408 6276
rect 35158 6264 35164 6276
rect 35216 6264 35222 6316
rect 37826 6264 37832 6316
rect 37884 6264 37890 6316
rect 38212 6313 38240 6344
rect 38197 6307 38255 6313
rect 38197 6273 38209 6307
rect 38243 6273 38255 6307
rect 38197 6267 38255 6273
rect 22612 6208 29408 6236
rect 22612 6196 22618 6208
rect 29454 6196 29460 6248
rect 29512 6236 29518 6248
rect 37550 6236 37556 6248
rect 29512 6208 37556 6236
rect 29512 6196 29518 6208
rect 37550 6196 37556 6208
rect 37608 6196 37614 6248
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 10042 6168 10048 6180
rect 7432 6140 10048 6168
rect 7432 6128 7438 6140
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 13814 6128 13820 6180
rect 13872 6168 13878 6180
rect 25406 6168 25412 6180
rect 13872 6140 25412 6168
rect 13872 6128 13878 6140
rect 25406 6128 25412 6140
rect 25464 6128 25470 6180
rect 27614 6128 27620 6180
rect 27672 6168 27678 6180
rect 30098 6168 30104 6180
rect 27672 6140 30104 6168
rect 27672 6128 27678 6140
rect 30098 6128 30104 6140
rect 30156 6128 30162 6180
rect 38013 6171 38071 6177
rect 38013 6137 38025 6171
rect 38059 6168 38071 6171
rect 39574 6168 39580 6180
rect 38059 6140 39580 6168
rect 38059 6137 38071 6140
rect 38013 6131 38071 6137
rect 39574 6128 39580 6140
rect 39632 6128 39638 6180
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 8113 6103 8171 6109
rect 8113 6100 8125 6103
rect 4396 6072 8125 6100
rect 4396 6060 4402 6072
rect 8113 6069 8125 6072
rect 8159 6069 8171 6103
rect 8113 6063 8171 6069
rect 10137 6103 10195 6109
rect 10137 6069 10149 6103
rect 10183 6100 10195 6103
rect 10410 6100 10416 6112
rect 10183 6072 10416 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 20438 6100 20444 6112
rect 10560 6072 20444 6100
rect 10560 6060 10566 6072
rect 20438 6060 20444 6072
rect 20496 6060 20502 6112
rect 22462 6060 22468 6112
rect 22520 6060 22526 6112
rect 26050 6060 26056 6112
rect 26108 6100 26114 6112
rect 34238 6100 34244 6112
rect 26108 6072 34244 6100
rect 26108 6060 26114 6072
rect 34238 6060 34244 6072
rect 34296 6060 34302 6112
rect 36906 6060 36912 6112
rect 36964 6100 36970 6112
rect 38286 6100 38292 6112
rect 36964 6072 38292 6100
rect 36964 6060 36970 6072
rect 38286 6060 38292 6072
rect 38344 6060 38350 6112
rect 1104 6010 38824 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 38824 6010
rect 1104 5936 38824 5958
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 11514 5896 11520 5908
rect 7892 5868 11520 5896
rect 7892 5856 7898 5868
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 17678 5856 17684 5908
rect 17736 5896 17742 5908
rect 23842 5896 23848 5908
rect 17736 5868 23848 5896
rect 17736 5856 17742 5868
rect 23842 5856 23848 5868
rect 23900 5856 23906 5908
rect 29454 5896 29460 5908
rect 28276 5868 29460 5896
rect 8294 5788 8300 5840
rect 8352 5828 8358 5840
rect 17586 5828 17592 5840
rect 8352 5800 17592 5828
rect 8352 5788 8358 5800
rect 17586 5788 17592 5800
rect 17644 5788 17650 5840
rect 23474 5828 23480 5840
rect 22066 5800 23480 5828
rect 12986 5720 12992 5772
rect 13044 5760 13050 5772
rect 22066 5760 22094 5800
rect 23474 5788 23480 5800
rect 23532 5788 23538 5840
rect 24762 5788 24768 5840
rect 24820 5828 24826 5840
rect 28276 5828 28304 5868
rect 29454 5856 29460 5868
rect 29512 5856 29518 5908
rect 31389 5899 31447 5905
rect 31389 5865 31401 5899
rect 31435 5896 31447 5899
rect 32858 5896 32864 5908
rect 31435 5868 32864 5896
rect 31435 5865 31447 5868
rect 31389 5859 31447 5865
rect 32858 5856 32864 5868
rect 32916 5856 32922 5908
rect 34885 5899 34943 5905
rect 34885 5865 34897 5899
rect 34931 5896 34943 5899
rect 36354 5896 36360 5908
rect 34931 5868 36360 5896
rect 34931 5865 34943 5868
rect 34885 5859 34943 5865
rect 36354 5856 36360 5868
rect 36412 5856 36418 5908
rect 37090 5856 37096 5908
rect 37148 5856 37154 5908
rect 37366 5856 37372 5908
rect 37424 5856 37430 5908
rect 24820 5800 28304 5828
rect 28353 5831 28411 5837
rect 24820 5788 24826 5800
rect 28353 5797 28365 5831
rect 28399 5828 28411 5831
rect 32766 5828 32772 5840
rect 28399 5800 32772 5828
rect 28399 5797 28411 5800
rect 28353 5791 28411 5797
rect 32766 5788 32772 5800
rect 32824 5788 32830 5840
rect 33321 5831 33379 5837
rect 33321 5797 33333 5831
rect 33367 5828 33379 5831
rect 35066 5828 35072 5840
rect 33367 5800 35072 5828
rect 33367 5797 33379 5800
rect 33321 5791 33379 5797
rect 35066 5788 35072 5800
rect 35124 5788 35130 5840
rect 36081 5831 36139 5837
rect 36081 5797 36093 5831
rect 36127 5828 36139 5831
rect 37274 5828 37280 5840
rect 36127 5800 37280 5828
rect 36127 5797 36139 5800
rect 36081 5791 36139 5797
rect 37274 5788 37280 5800
rect 37332 5788 37338 5840
rect 38378 5788 38384 5840
rect 38436 5788 38442 5840
rect 13044 5732 22094 5760
rect 13044 5720 13050 5732
rect 22462 5720 22468 5772
rect 22520 5760 22526 5772
rect 22520 5732 38240 5760
rect 22520 5720 22526 5732
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13320 5664 22094 5692
rect 13320 5652 13326 5664
rect 6454 5584 6460 5636
rect 6512 5624 6518 5636
rect 13354 5624 13360 5636
rect 6512 5596 13360 5624
rect 6512 5584 6518 5596
rect 13354 5584 13360 5596
rect 13412 5584 13418 5636
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 21634 5624 21640 5636
rect 19484 5596 21640 5624
rect 19484 5584 19490 5596
rect 21634 5584 21640 5596
rect 21692 5584 21698 5636
rect 22066 5624 22094 5664
rect 23566 5652 23572 5704
rect 23624 5692 23630 5704
rect 28169 5695 28227 5701
rect 28169 5692 28181 5695
rect 23624 5664 28181 5692
rect 23624 5652 23630 5664
rect 28169 5661 28181 5664
rect 28215 5661 28227 5695
rect 28169 5655 28227 5661
rect 29086 5652 29092 5704
rect 29144 5692 29150 5704
rect 31205 5695 31263 5701
rect 31205 5692 31217 5695
rect 29144 5664 31217 5692
rect 29144 5652 29150 5664
rect 31205 5661 31217 5664
rect 31251 5661 31263 5695
rect 33137 5695 33195 5701
rect 33137 5692 33149 5695
rect 31205 5655 31263 5661
rect 31726 5664 33149 5692
rect 24302 5624 24308 5636
rect 22066 5596 24308 5624
rect 24302 5584 24308 5596
rect 24360 5584 24366 5636
rect 30926 5584 30932 5636
rect 30984 5624 30990 5636
rect 31726 5624 31754 5664
rect 33137 5661 33149 5664
rect 33183 5661 33195 5695
rect 34701 5695 34759 5701
rect 34701 5692 34713 5695
rect 33137 5655 33195 5661
rect 33244 5664 34713 5692
rect 30984 5596 31754 5624
rect 30984 5584 30990 5596
rect 32766 5584 32772 5636
rect 32824 5624 32830 5636
rect 33244 5624 33272 5664
rect 34701 5661 34713 5664
rect 34747 5661 34759 5695
rect 34701 5655 34759 5661
rect 35897 5695 35955 5701
rect 35897 5661 35909 5695
rect 35943 5661 35955 5695
rect 35897 5655 35955 5661
rect 32824 5596 33272 5624
rect 32824 5584 32830 5596
rect 34606 5584 34612 5636
rect 34664 5624 34670 5636
rect 35912 5624 35940 5655
rect 36906 5652 36912 5704
rect 36964 5652 36970 5704
rect 38212 5701 38240 5732
rect 37177 5695 37235 5701
rect 37177 5692 37189 5695
rect 37016 5664 37189 5692
rect 34664 5596 35940 5624
rect 36004 5596 36216 5624
rect 34664 5584 34670 5596
rect 14274 5516 14280 5568
rect 14332 5556 14338 5568
rect 22830 5556 22836 5568
rect 14332 5528 22836 5556
rect 14332 5516 14338 5528
rect 22830 5516 22836 5528
rect 22888 5516 22894 5568
rect 23106 5516 23112 5568
rect 23164 5556 23170 5568
rect 34698 5556 34704 5568
rect 23164 5528 34704 5556
rect 23164 5516 23170 5528
rect 34698 5516 34704 5528
rect 34756 5516 34762 5568
rect 34790 5516 34796 5568
rect 34848 5556 34854 5568
rect 36004 5556 36032 5596
rect 34848 5528 36032 5556
rect 36188 5556 36216 5596
rect 36446 5584 36452 5636
rect 36504 5624 36510 5636
rect 37016 5624 37044 5664
rect 37177 5661 37189 5664
rect 37223 5661 37235 5695
rect 37177 5655 37235 5661
rect 37829 5695 37887 5701
rect 37829 5661 37841 5695
rect 37875 5661 37887 5695
rect 37829 5655 37887 5661
rect 38197 5695 38255 5701
rect 38197 5661 38209 5695
rect 38243 5661 38255 5695
rect 38197 5655 38255 5661
rect 36504 5596 37044 5624
rect 36504 5584 36510 5596
rect 37844 5556 37872 5655
rect 36188 5528 37872 5556
rect 34848 5516 34854 5528
rect 38010 5516 38016 5568
rect 38068 5516 38074 5568
rect 1104 5466 38824 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 38824 5466
rect 1104 5392 38824 5414
rect 19058 5312 19064 5364
rect 19116 5352 19122 5364
rect 37826 5352 37832 5364
rect 19116 5324 37832 5352
rect 19116 5312 19122 5324
rect 37826 5312 37832 5324
rect 37884 5312 37890 5364
rect 38378 5312 38384 5364
rect 38436 5312 38442 5364
rect 18138 5244 18144 5296
rect 18196 5284 18202 5296
rect 18196 5256 38240 5284
rect 18196 5244 18202 5256
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 19518 5216 19524 5228
rect 8444 5188 19524 5216
rect 8444 5176 8450 5188
rect 19518 5176 19524 5188
rect 19576 5176 19582 5228
rect 19610 5176 19616 5228
rect 19668 5176 19674 5228
rect 19702 5176 19708 5228
rect 19760 5176 19766 5228
rect 22002 5176 22008 5228
rect 22060 5216 22066 5228
rect 38212 5225 38240 5256
rect 28077 5219 28135 5225
rect 28077 5216 28089 5219
rect 22060 5188 28089 5216
rect 22060 5176 22066 5188
rect 28077 5185 28089 5188
rect 28123 5185 28135 5219
rect 37829 5219 37887 5225
rect 37829 5216 37841 5219
rect 28077 5179 28135 5185
rect 31726 5188 37841 5216
rect 18230 5108 18236 5160
rect 18288 5148 18294 5160
rect 31726 5148 31754 5188
rect 37829 5185 37841 5188
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 38197 5219 38255 5225
rect 38197 5185 38209 5219
rect 38243 5185 38255 5219
rect 38197 5179 38255 5185
rect 18288 5120 19564 5148
rect 18288 5108 18294 5120
rect 19536 5092 19564 5120
rect 19812 5120 31754 5148
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 19426 5080 19432 5092
rect 7616 5052 19432 5080
rect 7616 5040 7622 5052
rect 19426 5040 19432 5052
rect 19484 5040 19490 5092
rect 19518 5040 19524 5092
rect 19576 5040 19582 5092
rect 19702 5040 19708 5092
rect 19760 5080 19766 5092
rect 19812 5080 19840 5120
rect 19760 5052 19840 5080
rect 19889 5083 19947 5089
rect 19760 5040 19766 5052
rect 19889 5049 19901 5083
rect 19935 5080 19947 5083
rect 26878 5080 26884 5092
rect 19935 5052 26884 5080
rect 19935 5049 19947 5052
rect 19889 5043 19947 5049
rect 26878 5040 26884 5052
rect 26936 5040 26942 5092
rect 1118 4972 1124 5024
rect 1176 5012 1182 5024
rect 19334 5012 19340 5024
rect 1176 4984 19340 5012
rect 1176 4972 1182 4984
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 28261 5015 28319 5021
rect 28261 4981 28273 5015
rect 28307 5012 28319 5015
rect 35434 5012 35440 5024
rect 28307 4984 35440 5012
rect 28307 4981 28319 4984
rect 28261 4975 28319 4981
rect 35434 4972 35440 4984
rect 35492 4972 35498 5024
rect 38013 5015 38071 5021
rect 38013 4981 38025 5015
rect 38059 5012 38071 5015
rect 39114 5012 39120 5024
rect 38059 4984 39120 5012
rect 38059 4981 38071 4984
rect 38013 4975 38071 4981
rect 39114 4972 39120 4984
rect 39172 4972 39178 5024
rect 1104 4922 38824 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 38824 4922
rect 1104 4848 38824 4870
rect 38378 4700 38384 4752
rect 38436 4700 38442 4752
rect 13722 4632 13728 4684
rect 13780 4672 13786 4684
rect 21913 4675 21971 4681
rect 21913 4672 21925 4675
rect 13780 4644 21925 4672
rect 13780 4632 13786 4644
rect 21913 4641 21925 4644
rect 21959 4641 21971 4675
rect 21913 4635 21971 4641
rect 26878 4632 26884 4684
rect 26936 4672 26942 4684
rect 26936 4644 38240 4672
rect 26936 4632 26942 4644
rect 38212 4613 38240 4644
rect 21269 4607 21327 4613
rect 21269 4573 21281 4607
rect 21315 4604 21327 4607
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 21315 4576 21373 4604
rect 21315 4573 21327 4576
rect 21269 4567 21327 4573
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4604 22063 4607
rect 22097 4607 22155 4613
rect 22097 4604 22109 4607
rect 22051 4576 22109 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 22097 4573 22109 4576
rect 22143 4573 22155 4607
rect 37829 4607 37887 4613
rect 37829 4604 37841 4607
rect 22097 4567 22155 4573
rect 31726 4576 37841 4604
rect 21174 4496 21180 4548
rect 21232 4496 21238 4548
rect 31726 4536 31754 4576
rect 37829 4573 37841 4576
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 38197 4607 38255 4613
rect 38197 4573 38209 4607
rect 38243 4573 38255 4607
rect 38197 4567 38255 4573
rect 21560 4508 31754 4536
rect 21560 4477 21588 4508
rect 21545 4471 21603 4477
rect 21545 4437 21557 4471
rect 21591 4437 21603 4471
rect 21545 4431 21603 4437
rect 22281 4471 22339 4477
rect 22281 4437 22293 4471
rect 22327 4468 22339 4471
rect 26878 4468 26884 4480
rect 22327 4440 26884 4468
rect 22327 4437 22339 4440
rect 22281 4431 22339 4437
rect 26878 4428 26884 4440
rect 26936 4428 26942 4480
rect 38010 4428 38016 4480
rect 38068 4428 38074 4480
rect 1104 4378 38824 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 38824 4378
rect 1104 4304 38824 4326
rect 15381 4267 15439 4273
rect 15381 4233 15393 4267
rect 15427 4233 15439 4267
rect 15381 4227 15439 4233
rect 22066 4236 22600 4264
rect 15396 4140 15424 4227
rect 22066 4196 22094 4236
rect 18616 4168 19104 4196
rect 5166 4088 5172 4140
rect 5224 4128 5230 4140
rect 15197 4131 15255 4137
rect 15197 4128 15209 4131
rect 5224 4100 15209 4128
rect 5224 4088 5230 4100
rect 15197 4097 15209 4100
rect 15243 4097 15255 4131
rect 15197 4091 15255 4097
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 15470 4088 15476 4140
rect 15528 4088 15534 4140
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16531 4100 16681 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17589 4131 17647 4137
rect 17589 4128 17601 4131
rect 17543 4100 17601 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17589 4097 17601 4100
rect 17635 4097 17647 4131
rect 17589 4091 17647 4097
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4128 18383 4131
rect 18417 4131 18475 4137
rect 18417 4128 18429 4131
rect 18371 4100 18429 4128
rect 18371 4097 18383 4100
rect 18325 4091 18383 4097
rect 18417 4097 18429 4100
rect 18463 4097 18475 4131
rect 18616 4128 18644 4168
rect 18417 4091 18475 4097
rect 18524 4100 18644 4128
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 16132 4060 16160 4091
rect 3476 4032 16160 4060
rect 3476 4020 3482 4032
rect 7834 3952 7840 4004
rect 7892 3992 7898 4004
rect 15470 3992 15476 4004
rect 7892 3964 15476 3992
rect 7892 3952 7898 3964
rect 15470 3952 15476 3964
rect 15528 3952 15534 4004
rect 17052 3992 17080 4091
rect 17126 4020 17132 4072
rect 17184 4060 17190 4072
rect 18524 4060 18552 4100
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 18969 4131 19027 4137
rect 18969 4128 18981 4131
rect 18748 4100 18981 4128
rect 18748 4088 18754 4100
rect 18969 4097 18981 4100
rect 19015 4097 19027 4131
rect 19076 4128 19104 4168
rect 21744 4168 22094 4196
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19076 4100 19441 4128
rect 18969 4091 19027 4097
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19429 4091 19487 4097
rect 20438 4088 20444 4140
rect 20496 4088 20502 4140
rect 21177 4131 21235 4137
rect 21177 4097 21189 4131
rect 21223 4128 21235 4131
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 21223 4100 21281 4128
rect 21223 4097 21235 4100
rect 21177 4091 21235 4097
rect 21269 4097 21281 4100
rect 21315 4097 21327 4131
rect 21744 4128 21772 4168
rect 21269 4091 21327 4097
rect 21376 4100 21772 4128
rect 21376 4060 21404 4100
rect 21818 4088 21824 4140
rect 21876 4088 21882 4140
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 22373 4131 22431 4137
rect 22373 4128 22385 4131
rect 22327 4100 22385 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 22373 4097 22385 4100
rect 22419 4097 22431 4131
rect 22373 4091 22431 4097
rect 17184 4032 18552 4060
rect 18616 4032 21404 4060
rect 21468 4032 22232 4060
rect 17184 4020 17190 4032
rect 18616 4001 18644 4032
rect 21468 4001 21496 4032
rect 17865 3995 17923 4001
rect 17865 3992 17877 3995
rect 15580 3964 17877 3992
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15580 3924 15608 3964
rect 17865 3961 17877 3964
rect 17911 3961 17923 3995
rect 17865 3955 17923 3961
rect 18601 3995 18659 4001
rect 18601 3961 18613 3995
rect 18647 3961 18659 3995
rect 18601 3955 18659 3961
rect 21453 3995 21511 4001
rect 21453 3961 21465 3995
rect 21499 3961 21511 3995
rect 21453 3955 21511 3961
rect 22005 3995 22063 4001
rect 22005 3961 22017 3995
rect 22051 3992 22063 3995
rect 22094 3992 22100 4004
rect 22051 3964 22100 3992
rect 22051 3961 22063 3964
rect 22005 3955 22063 3961
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 22204 3992 22232 4032
rect 22462 3992 22468 4004
rect 22204 3964 22468 3992
rect 22462 3952 22468 3964
rect 22520 3952 22526 4004
rect 22572 3992 22600 4236
rect 26878 4156 26884 4208
rect 26936 4196 26942 4208
rect 26936 4168 31754 4196
rect 26936 4156 26942 4168
rect 22646 4088 22652 4140
rect 22704 4128 22710 4140
rect 22925 4131 22983 4137
rect 22925 4128 22937 4131
rect 22704 4100 22937 4128
rect 22704 4088 22710 4100
rect 22925 4097 22937 4100
rect 22971 4097 22983 4131
rect 22925 4091 22983 4097
rect 23106 4088 23112 4140
rect 23164 4128 23170 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 23164 4100 26985 4128
rect 23164 4088 23170 4100
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 31726 4060 31754 4168
rect 33778 4088 33784 4140
rect 33836 4128 33842 4140
rect 37829 4131 37887 4137
rect 37829 4128 37841 4131
rect 33836 4100 37841 4128
rect 33836 4088 33842 4100
rect 37829 4097 37841 4100
rect 37875 4097 37887 4131
rect 37829 4091 37887 4097
rect 38197 4131 38255 4137
rect 38197 4097 38209 4131
rect 38243 4097 38255 4131
rect 38197 4091 38255 4097
rect 38212 4060 38240 4091
rect 31726 4032 38240 4060
rect 37458 3992 37464 4004
rect 22572 3964 37464 3992
rect 37458 3952 37464 3964
rect 37516 3952 37522 4004
rect 38378 3952 38384 4004
rect 38436 3952 38442 4004
rect 15160 3896 15608 3924
rect 15160 3884 15166 3896
rect 15654 3884 15660 3936
rect 15712 3884 15718 3936
rect 16298 3884 16304 3936
rect 16356 3884 16362 3936
rect 16390 3884 16396 3936
rect 16448 3884 16454 3936
rect 16850 3884 16856 3936
rect 16908 3884 16914 3936
rect 17218 3884 17224 3936
rect 17276 3884 17282 3936
rect 17402 3884 17408 3936
rect 17460 3884 17466 3936
rect 17770 3884 17776 3936
rect 17828 3884 17834 3936
rect 18230 3884 18236 3936
rect 18288 3884 18294 3936
rect 18874 3884 18880 3936
rect 18932 3884 18938 3936
rect 19610 3884 19616 3936
rect 19668 3884 19674 3936
rect 20622 3884 20628 3936
rect 20680 3884 20686 3936
rect 20898 3884 20904 3936
rect 20956 3924 20962 3936
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20956 3896 21097 3924
rect 20956 3884 20962 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 21542 3884 21548 3936
rect 21600 3924 21606 3936
rect 21818 3924 21824 3936
rect 21600 3896 21824 3924
rect 21600 3884 21606 3896
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 22186 3884 22192 3936
rect 22244 3884 22250 3936
rect 22554 3884 22560 3936
rect 22612 3884 22618 3936
rect 22833 3927 22891 3933
rect 22833 3893 22845 3927
rect 22879 3924 22891 3927
rect 27062 3924 27068 3936
rect 22879 3896 27068 3924
rect 22879 3893 22891 3896
rect 22833 3887 22891 3893
rect 27062 3884 27068 3896
rect 27120 3884 27126 3936
rect 27157 3927 27215 3933
rect 27157 3893 27169 3927
rect 27203 3924 27215 3927
rect 27430 3924 27436 3936
rect 27203 3896 27436 3924
rect 27203 3893 27215 3896
rect 27157 3887 27215 3893
rect 27430 3884 27436 3896
rect 27488 3884 27494 3936
rect 38013 3927 38071 3933
rect 38013 3893 38025 3927
rect 38059 3924 38071 3927
rect 39114 3924 39120 3936
rect 38059 3896 39120 3924
rect 38059 3893 38071 3896
rect 38013 3887 38071 3893
rect 39114 3884 39120 3896
rect 39172 3884 39178 3936
rect 1104 3834 38824 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 38824 3834
rect 1104 3760 38824 3782
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 17126 3720 17132 3732
rect 8904 3692 17132 3720
rect 8904 3680 8910 3692
rect 17126 3680 17132 3692
rect 17184 3680 17190 3732
rect 18049 3723 18107 3729
rect 18049 3689 18061 3723
rect 18095 3720 18107 3723
rect 23014 3720 23020 3732
rect 18095 3692 23020 3720
rect 18095 3689 18107 3692
rect 18049 3683 18107 3689
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 37826 3720 37832 3732
rect 23124 3692 37832 3720
rect 9582 3612 9588 3664
rect 9640 3652 9646 3664
rect 18230 3652 18236 3664
rect 9640 3624 18236 3652
rect 9640 3612 9646 3624
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 22278 3612 22284 3664
rect 22336 3652 22342 3664
rect 23124 3652 23152 3692
rect 37826 3680 37832 3692
rect 37884 3680 37890 3732
rect 22336 3624 23152 3652
rect 22336 3612 22342 3624
rect 26418 3612 26424 3664
rect 26476 3652 26482 3664
rect 26881 3655 26939 3661
rect 26881 3652 26893 3655
rect 26476 3624 26893 3652
rect 26476 3612 26482 3624
rect 26881 3621 26893 3624
rect 26927 3621 26939 3655
rect 26881 3615 26939 3621
rect 27433 3655 27491 3661
rect 27433 3621 27445 3655
rect 27479 3652 27491 3655
rect 32398 3652 32404 3664
rect 27479 3624 32404 3652
rect 27479 3621 27491 3624
rect 27433 3615 27491 3621
rect 32398 3612 32404 3624
rect 32456 3612 32462 3664
rect 38378 3612 38384 3664
rect 38436 3612 38442 3664
rect 8570 3544 8576 3596
rect 8628 3584 8634 3596
rect 17402 3584 17408 3596
rect 8628 3556 17408 3584
rect 8628 3544 8634 3556
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 18046 3544 18052 3596
rect 18104 3584 18110 3596
rect 18104 3556 26188 3584
rect 18104 3544 18110 3556
rect 1486 3476 1492 3528
rect 1544 3516 1550 3528
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 1544 3488 17877 3516
rect 1544 3476 1550 3488
rect 17865 3485 17877 3488
rect 17911 3485 17923 3519
rect 17865 3479 17923 3485
rect 20346 3476 20352 3528
rect 20404 3516 20410 3528
rect 26160 3525 26188 3556
rect 27062 3544 27068 3596
rect 27120 3584 27126 3596
rect 27120 3556 31754 3584
rect 27120 3544 27126 3556
rect 21729 3519 21787 3525
rect 21729 3516 21741 3519
rect 20404 3488 21741 3516
rect 20404 3476 20410 3488
rect 21729 3485 21741 3488
rect 21775 3516 21787 3519
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21775 3488 21925 3516
rect 21775 3485 21787 3488
rect 21729 3479 21787 3485
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 25317 3519 25375 3525
rect 25317 3485 25329 3519
rect 25363 3516 25375 3519
rect 25409 3519 25467 3525
rect 25409 3516 25421 3519
rect 25363 3488 25421 3516
rect 25363 3485 25375 3488
rect 25317 3479 25375 3485
rect 25409 3485 25421 3488
rect 25455 3485 25467 3519
rect 25409 3479 25467 3485
rect 26145 3519 26203 3525
rect 26145 3485 26157 3519
rect 26191 3485 26203 3519
rect 26145 3479 26203 3485
rect 26605 3519 26663 3525
rect 26605 3485 26617 3519
rect 26651 3516 26663 3519
rect 26697 3519 26755 3525
rect 26697 3516 26709 3519
rect 26651 3488 26709 3516
rect 26651 3485 26663 3488
rect 26605 3479 26663 3485
rect 26697 3485 26709 3488
rect 26743 3485 26755 3519
rect 26697 3479 26755 3485
rect 26970 3476 26976 3528
rect 27028 3476 27034 3528
rect 27249 3519 27307 3525
rect 27249 3485 27261 3519
rect 27295 3485 27307 3519
rect 31726 3516 31754 3556
rect 37829 3519 37887 3525
rect 37829 3516 37841 3519
rect 31726 3488 37841 3516
rect 27249 3479 27307 3485
rect 37829 3485 37841 3488
rect 37875 3485 37887 3519
rect 37829 3479 37887 3485
rect 9490 3408 9496 3460
rect 9548 3448 9554 3460
rect 16390 3448 16396 3460
rect 9548 3420 16396 3448
rect 9548 3408 9554 3420
rect 16390 3408 16396 3420
rect 16448 3408 16454 3460
rect 23474 3408 23480 3460
rect 23532 3448 23538 3460
rect 27264 3448 27292 3479
rect 38194 3476 38200 3528
rect 38252 3476 38258 3528
rect 23532 3420 27292 3448
rect 23532 3408 23538 3420
rect 22094 3340 22100 3392
rect 22152 3340 22158 3392
rect 25222 3340 25228 3392
rect 25280 3340 25286 3392
rect 25590 3340 25596 3392
rect 25648 3340 25654 3392
rect 26326 3340 26332 3392
rect 26384 3340 26390 3392
rect 26510 3340 26516 3392
rect 26568 3340 26574 3392
rect 27157 3383 27215 3389
rect 27157 3349 27169 3383
rect 27203 3380 27215 3383
rect 27522 3380 27528 3392
rect 27203 3352 27528 3380
rect 27203 3349 27215 3352
rect 27157 3343 27215 3349
rect 27522 3340 27528 3352
rect 27580 3340 27586 3392
rect 38010 3340 38016 3392
rect 38068 3340 38074 3392
rect 1104 3290 38824 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 38824 3290
rect 1104 3216 38824 3238
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 38194 3176 38200 3188
rect 17276 3148 38200 3176
rect 17276 3136 17282 3148
rect 38194 3136 38200 3148
rect 38252 3136 38258 3188
rect 38378 3136 38384 3188
rect 38436 3136 38442 3188
rect 7006 3068 7012 3120
rect 7064 3108 7070 3120
rect 20438 3108 20444 3120
rect 7064 3080 20444 3108
rect 7064 3068 7070 3080
rect 20438 3068 20444 3080
rect 20496 3068 20502 3120
rect 22462 3068 22468 3120
rect 22520 3108 22526 3120
rect 22520 3080 38240 3108
rect 22520 3068 22526 3080
rect 16298 3000 16304 3052
rect 16356 3040 16362 3052
rect 24670 3040 24676 3052
rect 16356 3012 24676 3040
rect 16356 3000 16362 3012
rect 24670 3000 24676 3012
rect 24728 3000 24734 3052
rect 26234 3040 26240 3052
rect 25516 3012 26240 3040
rect 19610 2932 19616 2984
rect 19668 2972 19674 2984
rect 25516 2972 25544 3012
rect 26234 3000 26240 3012
rect 26292 3000 26298 3052
rect 26326 3000 26332 3052
rect 26384 3040 26390 3052
rect 34514 3040 34520 3052
rect 26384 3012 34520 3040
rect 26384 3000 26390 3012
rect 34514 3000 34520 3012
rect 34572 3000 34578 3052
rect 37458 3000 37464 3052
rect 37516 3000 37522 3052
rect 37826 3000 37832 3052
rect 37884 3000 37890 3052
rect 38212 3049 38240 3080
rect 38197 3043 38255 3049
rect 38197 3009 38209 3043
rect 38243 3009 38255 3043
rect 38197 3003 38255 3009
rect 19668 2944 25544 2972
rect 19668 2932 19674 2944
rect 25590 2932 25596 2984
rect 25648 2972 25654 2984
rect 31846 2972 31852 2984
rect 25648 2944 31852 2972
rect 25648 2932 25654 2944
rect 31846 2932 31852 2944
rect 31904 2932 31910 2984
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 32674 2904 32680 2916
rect 20680 2876 22140 2904
rect 20680 2864 20686 2876
rect 22112 2836 22140 2876
rect 25608 2876 32680 2904
rect 25608 2836 25636 2876
rect 32674 2864 32680 2876
rect 32732 2864 32738 2916
rect 22112 2808 25636 2836
rect 26234 2796 26240 2848
rect 26292 2836 26298 2848
rect 33502 2836 33508 2848
rect 26292 2808 33508 2836
rect 26292 2796 26298 2808
rect 33502 2796 33508 2808
rect 33560 2796 33566 2848
rect 37645 2839 37703 2845
rect 37645 2805 37657 2839
rect 37691 2836 37703 2839
rect 37826 2836 37832 2848
rect 37691 2808 37832 2836
rect 37691 2805 37703 2808
rect 37645 2799 37703 2805
rect 37826 2796 37832 2808
rect 37884 2796 37890 2848
rect 38013 2839 38071 2845
rect 38013 2805 38025 2839
rect 38059 2836 38071 2839
rect 39114 2836 39120 2848
rect 38059 2808 39120 2836
rect 38059 2805 38071 2808
rect 38013 2799 38071 2805
rect 39114 2796 39120 2808
rect 39172 2796 39178 2848
rect 1104 2746 38824 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 38824 2746
rect 1104 2672 38824 2694
rect 18874 2592 18880 2644
rect 18932 2632 18938 2644
rect 36354 2632 36360 2644
rect 18932 2604 36360 2632
rect 18932 2592 18938 2604
rect 36354 2592 36360 2604
rect 36412 2592 36418 2644
rect 17770 2524 17776 2576
rect 17828 2564 17834 2576
rect 23658 2564 23664 2576
rect 17828 2536 23664 2564
rect 17828 2524 17834 2536
rect 23658 2524 23664 2536
rect 23716 2524 23722 2576
rect 24136 2536 36584 2564
rect 16850 2456 16856 2508
rect 16908 2496 16914 2508
rect 24136 2496 24164 2536
rect 16908 2468 24164 2496
rect 36556 2496 36584 2536
rect 36630 2524 36636 2576
rect 36688 2524 36694 2576
rect 36998 2524 37004 2576
rect 37056 2524 37062 2576
rect 38378 2524 38384 2576
rect 38436 2524 38442 2576
rect 36556 2468 37872 2496
rect 16908 2456 16914 2468
rect 15654 2388 15660 2440
rect 15712 2428 15718 2440
rect 15712 2400 22094 2428
rect 15712 2388 15718 2400
rect 22066 2360 22094 2400
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 23716 2400 36308 2428
rect 23716 2388 23722 2400
rect 36280 2360 36308 2400
rect 36354 2388 36360 2440
rect 36412 2428 36418 2440
rect 37844 2437 37872 2468
rect 36449 2431 36507 2437
rect 36449 2428 36461 2431
rect 36412 2400 36461 2428
rect 36412 2388 36418 2400
rect 36449 2397 36461 2400
rect 36495 2397 36507 2431
rect 36817 2431 36875 2437
rect 36817 2428 36829 2431
rect 36449 2391 36507 2397
rect 36556 2400 36829 2428
rect 36556 2360 36584 2400
rect 36817 2397 36829 2400
rect 36863 2397 36875 2431
rect 36817 2391 36875 2397
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 37829 2431 37887 2437
rect 37829 2397 37841 2431
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 37476 2360 37504 2391
rect 38194 2388 38200 2440
rect 38252 2388 38258 2440
rect 22066 2332 36216 2360
rect 36280 2332 36584 2360
rect 36648 2332 37504 2360
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 34974 2292 34980 2304
rect 22612 2264 34980 2292
rect 22612 2252 22618 2264
rect 34974 2252 34980 2264
rect 35032 2252 35038 2304
rect 36188 2292 36216 2332
rect 36648 2292 36676 2332
rect 36188 2264 36676 2292
rect 37642 2252 37648 2304
rect 37700 2252 37706 2304
rect 38010 2252 38016 2304
rect 38068 2252 38074 2304
rect 1104 2202 38824 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 38824 2202
rect 1104 2128 38824 2150
rect 14366 2048 14372 2100
rect 14424 2088 14430 2100
rect 23474 2088 23480 2100
rect 14424 2060 23480 2088
rect 14424 2048 14430 2060
rect 23474 2048 23480 2060
rect 23532 2048 23538 2100
rect 34974 2048 34980 2100
rect 35032 2088 35038 2100
rect 38194 2088 38200 2100
rect 35032 2060 38200 2088
rect 35032 2048 35038 2060
rect 38194 2048 38200 2060
rect 38252 2048 38258 2100
rect 19886 1504 19892 1556
rect 19944 1544 19950 1556
rect 23106 1544 23112 1556
rect 19944 1516 23112 1544
rect 19944 1504 19950 1516
rect 23106 1504 23112 1516
rect 23164 1504 23170 1556
<< via1 >>
rect 10416 11024 10468 11076
rect 10968 11024 11020 11076
rect 7380 10956 7432 11008
rect 17960 10956 18012 11008
rect 22192 11024 22244 11076
rect 22376 10956 22428 11008
rect 11428 10888 11480 10940
rect 21548 10888 21600 10940
rect 14464 10820 14516 10872
rect 23204 10820 23256 10872
rect 11520 10752 11572 10804
rect 20720 10752 20772 10804
rect 23388 10140 23440 10192
rect 25964 10140 26016 10192
rect 21548 10072 21600 10124
rect 24584 10072 24636 10124
rect 25872 10004 25924 10056
rect 31208 10004 31260 10056
rect 13360 9936 13412 9988
rect 18512 9936 18564 9988
rect 13636 9868 13688 9920
rect 17684 9868 17736 9920
rect 25596 9868 25648 9920
rect 30932 9868 30984 9920
rect 16672 9800 16724 9852
rect 25688 9800 25740 9852
rect 13912 9732 13964 9784
rect 18788 9732 18840 9784
rect 30380 9732 30432 9784
rect 1308 9664 1360 9716
rect 21824 9664 21876 9716
rect 25688 9664 25740 9716
rect 25780 9664 25832 9716
rect 30656 9664 30708 9716
rect 14556 9528 14608 9580
rect 17408 9528 17460 9580
rect 14188 9392 14240 9444
rect 26608 9392 26660 9444
rect 16120 9324 16172 9376
rect 28816 9324 28868 9376
rect 10692 9256 10744 9308
rect 15844 9256 15896 9308
rect 15936 9256 15988 9308
rect 28908 9256 28960 9308
rect 11980 9188 12032 9240
rect 13912 9188 13964 9240
rect 15660 9188 15712 9240
rect 29368 9188 29420 9240
rect 1124 9120 1176 9172
rect 22100 9120 22152 9172
rect 27436 9120 27488 9172
rect 34888 9120 34940 9172
rect 8392 9052 8444 9104
rect 17040 9052 17092 9104
rect 24676 9052 24728 9104
rect 32128 9052 32180 9104
rect 13176 8984 13228 9036
rect 15568 8984 15620 9036
rect 16212 8984 16264 9036
rect 19892 8984 19944 9036
rect 28448 8984 28500 9036
rect 35808 8984 35860 9036
rect 7840 8916 7892 8968
rect 18236 8916 18288 8968
rect 22284 8916 22336 8968
rect 38200 8916 38252 8968
rect 4252 8848 4304 8900
rect 10140 8848 10192 8900
rect 12808 8848 12860 8900
rect 24216 8848 24268 8900
rect 31852 8848 31904 8900
rect 33600 8848 33652 8900
rect 4896 8780 4948 8832
rect 6460 8780 6512 8832
rect 9496 8780 9548 8832
rect 14832 8780 14884 8832
rect 17592 8780 17644 8832
rect 19616 8780 19668 8832
rect 33140 8780 33192 8832
rect 34152 8780 34204 8832
rect 35348 8780 35400 8832
rect 35716 8780 35768 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 2780 8576 2832 8628
rect 3424 8576 3476 8628
rect 4436 8576 4488 8628
rect 4712 8576 4764 8628
rect 4988 8576 5040 8628
rect 5540 8576 5592 8628
rect 5816 8576 5868 8628
rect 6368 8576 6420 8628
rect 6920 8576 6972 8628
rect 7196 8576 7248 8628
rect 7748 8576 7800 8628
rect 8024 8576 8076 8628
rect 8484 8576 8536 8628
rect 8760 8576 8812 8628
rect 9404 8576 9456 8628
rect 9956 8576 10008 8628
rect 10232 8576 10284 8628
rect 10508 8576 10560 8628
rect 11060 8576 11112 8628
rect 11612 8576 11664 8628
rect 12164 8576 12216 8628
rect 12440 8576 12492 8628
rect 12716 8576 12768 8628
rect 13268 8576 13320 8628
rect 14096 8576 14148 8628
rect 14648 8576 14700 8628
rect 14924 8576 14976 8628
rect 15476 8576 15528 8628
rect 15752 8576 15804 8628
rect 16028 8576 16080 8628
rect 16304 8619 16356 8628
rect 16304 8585 16313 8619
rect 16313 8585 16347 8619
rect 16347 8585 16356 8619
rect 16304 8576 16356 8585
rect 16856 8576 16908 8628
rect 1216 8304 1268 8356
rect 1676 8304 1728 8356
rect 4252 8440 4304 8492
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4896 8440 4948 8492
rect 6828 8508 6880 8560
rect 5448 8483 5500 8492
rect 5448 8449 5450 8483
rect 5450 8449 5484 8483
rect 5484 8449 5500 8483
rect 5448 8440 5500 8449
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 5356 8372 5408 8424
rect 7196 8440 7248 8492
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 3884 8304 3936 8356
rect 6368 8304 6420 8356
rect 7564 8372 7616 8424
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 10692 8508 10744 8560
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9588 8304 9640 8356
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 11244 8440 11296 8492
rect 11796 8440 11848 8492
rect 14280 8508 14332 8560
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 17684 8576 17736 8628
rect 25412 8576 25464 8628
rect 31484 8576 31536 8628
rect 31760 8576 31812 8628
rect 32404 8576 32456 8628
rect 13452 8372 13504 8424
rect 5816 8236 5868 8288
rect 9864 8236 9916 8288
rect 13176 8304 13228 8356
rect 13820 8304 13872 8356
rect 14188 8372 14240 8424
rect 15660 8440 15712 8492
rect 15936 8440 15988 8492
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 16304 8440 16356 8492
rect 27988 8508 28040 8560
rect 32588 8508 32640 8560
rect 33968 8576 34020 8628
rect 35072 8576 35124 8628
rect 36452 8576 36504 8628
rect 17500 8440 17552 8492
rect 23020 8440 23072 8492
rect 32128 8483 32180 8492
rect 32128 8449 32137 8483
rect 32137 8449 32171 8483
rect 32171 8449 32180 8483
rect 32128 8440 32180 8449
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 32496 8440 32548 8449
rect 32680 8440 32732 8492
rect 33508 8440 33560 8492
rect 33600 8483 33652 8492
rect 33600 8449 33609 8483
rect 33609 8449 33643 8483
rect 33643 8449 33652 8483
rect 33600 8440 33652 8449
rect 16120 8304 16172 8356
rect 16580 8304 16632 8356
rect 11060 8236 11112 8288
rect 12624 8236 12676 8288
rect 17776 8236 17828 8288
rect 26148 8372 26200 8424
rect 26424 8372 26476 8424
rect 27712 8304 27764 8356
rect 28356 8304 28408 8356
rect 32036 8304 32088 8356
rect 32864 8304 32916 8356
rect 34612 8440 34664 8492
rect 34888 8440 34940 8492
rect 35440 8483 35492 8492
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 35624 8440 35676 8492
rect 34520 8372 34572 8424
rect 35808 8483 35860 8492
rect 35808 8449 35817 8483
rect 35817 8449 35851 8483
rect 35851 8449 35860 8483
rect 35808 8440 35860 8449
rect 35992 8440 36044 8492
rect 36728 8508 36780 8560
rect 37280 8483 37332 8492
rect 37280 8449 37289 8483
rect 37289 8449 37323 8483
rect 37323 8449 37332 8483
rect 37280 8440 37332 8449
rect 37372 8440 37424 8492
rect 38200 8483 38252 8492
rect 38200 8449 38209 8483
rect 38209 8449 38243 8483
rect 38243 8449 38252 8483
rect 38200 8440 38252 8449
rect 29644 8236 29696 8288
rect 32956 8236 33008 8288
rect 34152 8347 34204 8356
rect 34152 8313 34161 8347
rect 34161 8313 34195 8347
rect 34195 8313 34204 8347
rect 34152 8304 34204 8313
rect 34244 8304 34296 8356
rect 35716 8304 35768 8356
rect 38384 8347 38436 8356
rect 38384 8313 38393 8347
rect 38393 8313 38427 8347
rect 38427 8313 38436 8347
rect 38384 8304 38436 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 2872 8032 2924 8084
rect 3608 8032 3660 8084
rect 4160 8032 4212 8084
rect 5264 8032 5316 8084
rect 6092 8032 6144 8084
rect 6644 8032 6696 8084
rect 7472 8032 7524 8084
rect 8300 8032 8352 8084
rect 8852 8032 8904 8084
rect 9680 8032 9732 8084
rect 10784 8032 10836 8084
rect 11336 8032 11388 8084
rect 11888 8032 11940 8084
rect 12992 8032 13044 8084
rect 13544 8032 13596 8084
rect 14372 8032 14424 8084
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 17776 8032 17828 8084
rect 19064 8032 19116 8084
rect 29000 8032 29052 8084
rect 29920 8032 29972 8084
rect 33416 8032 33468 8084
rect 33784 8032 33836 8084
rect 34796 8032 34848 8084
rect 35900 8032 35952 8084
rect 36268 8032 36320 8084
rect 36912 8075 36964 8084
rect 36912 8041 36921 8075
rect 36921 8041 36955 8075
rect 36955 8041 36964 8075
rect 36912 8032 36964 8041
rect 37004 8032 37056 8084
rect 38660 8032 38712 8084
rect 5632 7964 5684 8016
rect 14648 7964 14700 8016
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 6736 7896 6788 7948
rect 6000 7828 6052 7880
rect 6920 7828 6972 7880
rect 8484 7896 8536 7948
rect 8300 7828 8352 7880
rect 16764 7896 16816 7948
rect 32772 7896 32824 7948
rect 9496 7871 9548 7880
rect 9496 7837 9505 7871
rect 9505 7837 9539 7871
rect 9539 7837 9548 7871
rect 9496 7828 9548 7837
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 13728 7828 13780 7880
rect 14648 7828 14700 7880
rect 6092 7760 6144 7812
rect 6184 7760 6236 7812
rect 11980 7760 12032 7812
rect 30012 7828 30064 7880
rect 32404 7828 32456 7880
rect 34980 7896 35032 7948
rect 18420 7760 18472 7812
rect 22008 7760 22060 7812
rect 33784 7760 33836 7812
rect 7012 7692 7064 7744
rect 13636 7692 13688 7744
rect 15568 7692 15620 7744
rect 23388 7692 23440 7744
rect 31760 7692 31812 7744
rect 35072 7828 35124 7880
rect 36360 7871 36412 7880
rect 36360 7837 36369 7871
rect 36369 7837 36403 7871
rect 36403 7837 36412 7871
rect 36360 7828 36412 7837
rect 36728 7871 36780 7880
rect 36728 7837 36737 7871
rect 36737 7837 36771 7871
rect 36771 7837 36780 7871
rect 36728 7828 36780 7837
rect 37096 7871 37148 7880
rect 37096 7837 37105 7871
rect 37105 7837 37139 7871
rect 37139 7837 37148 7871
rect 37096 7828 37148 7837
rect 37464 7871 37516 7880
rect 37464 7837 37473 7871
rect 37473 7837 37507 7871
rect 37507 7837 37516 7871
rect 37464 7828 37516 7837
rect 35164 7760 35216 7812
rect 38016 7735 38068 7744
rect 38016 7701 38025 7735
rect 38025 7701 38059 7735
rect 38059 7701 38068 7735
rect 38016 7692 38068 7701
rect 38384 7735 38436 7744
rect 38384 7701 38393 7735
rect 38393 7701 38427 7735
rect 38427 7701 38436 7735
rect 38384 7692 38436 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 4068 7488 4120 7540
rect 5356 7488 5408 7540
rect 5540 7488 5592 7540
rect 6000 7531 6052 7540
rect 6000 7497 6009 7531
rect 6009 7497 6043 7531
rect 6043 7497 6052 7531
rect 6000 7488 6052 7497
rect 6092 7488 6144 7540
rect 6920 7488 6972 7540
rect 5816 7420 5868 7472
rect 6460 7420 6512 7472
rect 10048 7488 10100 7540
rect 14832 7488 14884 7540
rect 9496 7420 9548 7472
rect 15844 7488 15896 7540
rect 16764 7531 16816 7540
rect 16764 7497 16773 7531
rect 16773 7497 16807 7531
rect 16807 7497 16816 7531
rect 16764 7488 16816 7497
rect 17040 7531 17092 7540
rect 17040 7497 17049 7531
rect 17049 7497 17083 7531
rect 17083 7497 17092 7531
rect 17040 7488 17092 7497
rect 20996 7488 21048 7540
rect 22284 7531 22336 7540
rect 22284 7497 22293 7531
rect 22293 7497 22327 7531
rect 22327 7497 22336 7531
rect 22284 7488 22336 7497
rect 22468 7531 22520 7540
rect 22468 7497 22477 7531
rect 22477 7497 22511 7531
rect 22511 7497 22520 7531
rect 22468 7488 22520 7497
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6920 7352 6972 7404
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 10140 7352 10192 7404
rect 13728 7352 13780 7404
rect 6368 7216 6420 7268
rect 12624 7284 12676 7336
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 14740 7352 14792 7404
rect 16672 7420 16724 7472
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 16488 7352 16540 7404
rect 19524 7420 19576 7472
rect 17224 7395 17276 7404
rect 17224 7361 17233 7395
rect 17233 7361 17267 7395
rect 17267 7361 17276 7395
rect 17224 7352 17276 7361
rect 19708 7395 19760 7404
rect 19708 7361 19717 7395
rect 19717 7361 19751 7395
rect 19751 7361 19760 7395
rect 19708 7352 19760 7361
rect 19984 7395 20036 7404
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 20352 7395 20404 7404
rect 20352 7361 20361 7395
rect 20361 7361 20395 7395
rect 20395 7361 20404 7395
rect 20352 7352 20404 7361
rect 20720 7284 20772 7336
rect 26792 7420 26844 7472
rect 28816 7531 28868 7540
rect 28816 7497 28825 7531
rect 28825 7497 28859 7531
rect 28859 7497 28868 7531
rect 28816 7488 28868 7497
rect 37464 7488 37516 7540
rect 37648 7531 37700 7540
rect 37648 7497 37657 7531
rect 37657 7497 37691 7531
rect 37691 7497 37700 7531
rect 37648 7488 37700 7497
rect 38292 7488 38344 7540
rect 33784 7420 33836 7472
rect 21364 7352 21416 7404
rect 21824 7395 21876 7404
rect 21824 7361 21833 7395
rect 21833 7361 21867 7395
rect 21867 7361 21876 7395
rect 21824 7352 21876 7361
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 22928 7395 22980 7404
rect 22928 7361 22937 7395
rect 22937 7361 22971 7395
rect 22971 7361 22980 7395
rect 22928 7352 22980 7361
rect 25872 7352 25924 7404
rect 27896 7352 27948 7404
rect 29460 7395 29512 7404
rect 29460 7361 29469 7395
rect 29469 7361 29503 7395
rect 29503 7361 29512 7395
rect 29460 7352 29512 7361
rect 29736 7395 29788 7404
rect 29736 7361 29745 7395
rect 29745 7361 29779 7395
rect 29779 7361 29788 7395
rect 29736 7352 29788 7361
rect 29920 7352 29972 7404
rect 30288 7395 30340 7404
rect 30288 7361 30297 7395
rect 30297 7361 30331 7395
rect 30331 7361 30340 7395
rect 30288 7352 30340 7361
rect 34244 7352 34296 7404
rect 7840 7216 7892 7268
rect 11244 7216 11296 7268
rect 13452 7216 13504 7268
rect 6920 7148 6972 7200
rect 7380 7148 7432 7200
rect 11060 7148 11112 7200
rect 14372 7148 14424 7200
rect 16396 7216 16448 7268
rect 19340 7216 19392 7268
rect 14648 7148 14700 7200
rect 17684 7148 17736 7200
rect 18696 7191 18748 7200
rect 18696 7157 18705 7191
rect 18705 7157 18739 7191
rect 18739 7157 18748 7191
rect 18696 7148 18748 7157
rect 19064 7191 19116 7200
rect 19064 7157 19073 7191
rect 19073 7157 19107 7191
rect 19107 7157 19116 7191
rect 19064 7148 19116 7157
rect 23388 7216 23440 7268
rect 24216 7259 24268 7268
rect 24216 7225 24225 7259
rect 24225 7225 24259 7259
rect 24259 7225 24268 7259
rect 24216 7216 24268 7225
rect 26792 7216 26844 7268
rect 34980 7216 35032 7268
rect 37004 7259 37056 7268
rect 37004 7225 37013 7259
rect 37013 7225 37047 7259
rect 37047 7225 37056 7259
rect 37004 7216 37056 7225
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 22008 7191 22060 7200
rect 22008 7157 22017 7191
rect 22017 7157 22051 7191
rect 22051 7157 22060 7191
rect 22008 7148 22060 7157
rect 24768 7148 24820 7200
rect 28908 7148 28960 7200
rect 29368 7148 29420 7200
rect 29644 7148 29696 7200
rect 30012 7148 30064 7200
rect 34704 7148 34756 7200
rect 38384 7191 38436 7200
rect 38384 7157 38393 7191
rect 38393 7157 38427 7191
rect 38427 7157 38436 7191
rect 38384 7148 38436 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 8484 6944 8536 6996
rect 12256 6944 12308 6996
rect 13728 6944 13780 6996
rect 20812 6944 20864 6996
rect 7288 6808 7340 6860
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 7840 6740 7892 6792
rect 11060 6808 11112 6860
rect 11152 6808 11204 6860
rect 13176 6808 13228 6860
rect 21456 6876 21508 6928
rect 36728 6944 36780 6996
rect 22100 6808 22152 6860
rect 22192 6851 22244 6860
rect 22192 6817 22201 6851
rect 22201 6817 22235 6851
rect 22235 6817 22244 6851
rect 22192 6808 22244 6817
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 23848 6808 23900 6860
rect 26148 6876 26200 6928
rect 25780 6808 25832 6860
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 6736 6672 6788 6724
rect 5448 6604 5500 6656
rect 7564 6647 7616 6656
rect 7564 6613 7573 6647
rect 7573 6613 7607 6647
rect 7607 6613 7616 6647
rect 7564 6604 7616 6613
rect 7748 6604 7800 6656
rect 9404 6604 9456 6656
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 10324 6740 10376 6792
rect 10600 6740 10652 6792
rect 10232 6647 10284 6656
rect 10232 6613 10241 6647
rect 10241 6613 10275 6647
rect 10275 6613 10284 6647
rect 10232 6604 10284 6613
rect 12716 6672 12768 6724
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 12992 6740 13044 6749
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 17868 6740 17920 6792
rect 11428 6604 11480 6656
rect 11796 6604 11848 6656
rect 14464 6672 14516 6724
rect 19248 6672 19300 6724
rect 14188 6604 14240 6656
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 18144 6647 18196 6656
rect 18144 6613 18153 6647
rect 18153 6613 18187 6647
rect 18187 6613 18196 6647
rect 18144 6604 18196 6613
rect 19340 6647 19392 6656
rect 19340 6613 19349 6647
rect 19349 6613 19383 6647
rect 19383 6613 19392 6647
rect 19340 6604 19392 6613
rect 19524 6604 19576 6656
rect 25596 6783 25648 6792
rect 25596 6749 25605 6783
rect 25605 6749 25639 6783
rect 25639 6749 25648 6783
rect 25596 6740 25648 6749
rect 25688 6740 25740 6792
rect 26332 6808 26384 6860
rect 28264 6876 28316 6928
rect 29828 6808 29880 6860
rect 34980 6808 35032 6860
rect 26884 6740 26936 6792
rect 27252 6740 27304 6792
rect 26056 6672 26108 6724
rect 27620 6783 27672 6792
rect 27620 6749 27629 6783
rect 27629 6749 27663 6783
rect 27663 6749 27672 6783
rect 27620 6740 27672 6749
rect 28356 6783 28408 6792
rect 28356 6749 28365 6783
rect 28365 6749 28399 6783
rect 28399 6749 28408 6783
rect 28356 6740 28408 6749
rect 29276 6740 29328 6792
rect 37464 6783 37516 6792
rect 37464 6749 37473 6783
rect 37473 6749 37507 6783
rect 37507 6749 37516 6783
rect 37464 6740 37516 6749
rect 37556 6740 37608 6792
rect 29552 6672 29604 6724
rect 22100 6604 22152 6656
rect 22560 6647 22612 6656
rect 22560 6613 22569 6647
rect 22569 6613 22603 6647
rect 22603 6613 22612 6647
rect 22560 6604 22612 6613
rect 23112 6647 23164 6656
rect 23112 6613 23121 6647
rect 23121 6613 23155 6647
rect 23155 6613 23164 6647
rect 23112 6604 23164 6613
rect 25412 6647 25464 6656
rect 25412 6613 25421 6647
rect 25421 6613 25455 6647
rect 25455 6613 25464 6647
rect 25412 6604 25464 6613
rect 25504 6604 25556 6656
rect 26608 6604 26660 6656
rect 27436 6647 27488 6656
rect 27436 6613 27445 6647
rect 27445 6613 27479 6647
rect 27479 6613 27488 6647
rect 27436 6604 27488 6613
rect 27896 6647 27948 6656
rect 27896 6613 27905 6647
rect 27905 6613 27939 6647
rect 27939 6613 27948 6647
rect 27896 6604 27948 6613
rect 28080 6604 28132 6656
rect 28356 6604 28408 6656
rect 28540 6647 28592 6656
rect 28540 6613 28549 6647
rect 28549 6613 28583 6647
rect 28583 6613 28592 6647
rect 28540 6604 28592 6613
rect 37648 6647 37700 6656
rect 37648 6613 37657 6647
rect 37657 6613 37691 6647
rect 37691 6613 37700 6647
rect 37648 6604 37700 6613
rect 38568 6672 38620 6724
rect 38476 6604 38528 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 7196 6400 7248 6452
rect 9404 6400 9456 6452
rect 9588 6400 9640 6452
rect 10324 6400 10376 6452
rect 11704 6400 11756 6452
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8760 6264 8812 6316
rect 9956 6264 10008 6316
rect 10416 6307 10468 6316
rect 10416 6273 10417 6307
rect 10417 6273 10451 6307
rect 10451 6273 10468 6307
rect 10416 6264 10468 6273
rect 10968 6264 11020 6316
rect 16856 6400 16908 6452
rect 17316 6400 17368 6452
rect 22100 6400 22152 6452
rect 22192 6400 22244 6452
rect 18236 6332 18288 6384
rect 18420 6332 18472 6384
rect 27896 6332 27948 6384
rect 28448 6443 28500 6452
rect 28448 6409 28457 6443
rect 28457 6409 28491 6443
rect 28491 6409 28500 6443
rect 28448 6400 28500 6409
rect 35992 6400 36044 6452
rect 38384 6443 38436 6452
rect 38384 6409 38393 6443
rect 38393 6409 38427 6443
rect 38427 6409 38436 6443
rect 38384 6400 38436 6409
rect 37464 6332 37516 6384
rect 37740 6332 37792 6384
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 16764 6264 16816 6273
rect 7104 6196 7156 6248
rect 10232 6196 10284 6248
rect 12716 6196 12768 6248
rect 17224 6264 17276 6316
rect 21548 6264 21600 6316
rect 21640 6264 21692 6316
rect 19800 6196 19852 6248
rect 22100 6196 22152 6248
rect 23756 6264 23808 6316
rect 25504 6264 25556 6316
rect 29276 6307 29328 6316
rect 29276 6273 29285 6307
rect 29285 6273 29319 6307
rect 29319 6273 29328 6307
rect 29276 6264 29328 6273
rect 22560 6196 22612 6248
rect 35164 6264 35216 6316
rect 37832 6307 37884 6316
rect 37832 6273 37841 6307
rect 37841 6273 37875 6307
rect 37875 6273 37884 6307
rect 37832 6264 37884 6273
rect 29460 6196 29512 6248
rect 37556 6196 37608 6248
rect 7380 6128 7432 6180
rect 10048 6128 10100 6180
rect 13820 6128 13872 6180
rect 25412 6128 25464 6180
rect 27620 6128 27672 6180
rect 30104 6128 30156 6180
rect 39580 6128 39632 6180
rect 4344 6060 4396 6112
rect 10416 6060 10468 6112
rect 10508 6060 10560 6112
rect 20444 6060 20496 6112
rect 22468 6103 22520 6112
rect 22468 6069 22477 6103
rect 22477 6069 22511 6103
rect 22511 6069 22520 6103
rect 22468 6060 22520 6069
rect 26056 6060 26108 6112
rect 34244 6060 34296 6112
rect 36912 6060 36964 6112
rect 38292 6060 38344 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 7840 5856 7892 5908
rect 11520 5856 11572 5908
rect 17684 5856 17736 5908
rect 23848 5856 23900 5908
rect 8300 5788 8352 5840
rect 17592 5788 17644 5840
rect 12992 5720 13044 5772
rect 23480 5788 23532 5840
rect 24768 5788 24820 5840
rect 29460 5856 29512 5908
rect 32864 5856 32916 5908
rect 36360 5856 36412 5908
rect 37096 5899 37148 5908
rect 37096 5865 37105 5899
rect 37105 5865 37139 5899
rect 37139 5865 37148 5899
rect 37096 5856 37148 5865
rect 37372 5899 37424 5908
rect 37372 5865 37381 5899
rect 37381 5865 37415 5899
rect 37415 5865 37424 5899
rect 37372 5856 37424 5865
rect 32772 5788 32824 5840
rect 35072 5788 35124 5840
rect 37280 5788 37332 5840
rect 38384 5831 38436 5840
rect 38384 5797 38393 5831
rect 38393 5797 38427 5831
rect 38427 5797 38436 5831
rect 38384 5788 38436 5797
rect 22468 5720 22520 5772
rect 13268 5652 13320 5704
rect 6460 5584 6512 5636
rect 13360 5584 13412 5636
rect 19432 5584 19484 5636
rect 21640 5584 21692 5636
rect 23572 5652 23624 5704
rect 29092 5652 29144 5704
rect 24308 5584 24360 5636
rect 30932 5584 30984 5636
rect 32772 5584 32824 5636
rect 34612 5584 34664 5636
rect 36912 5695 36964 5704
rect 36912 5661 36921 5695
rect 36921 5661 36955 5695
rect 36955 5661 36964 5695
rect 36912 5652 36964 5661
rect 14280 5516 14332 5568
rect 22836 5516 22888 5568
rect 23112 5516 23164 5568
rect 34704 5516 34756 5568
rect 34796 5516 34848 5568
rect 36452 5584 36504 5636
rect 38016 5559 38068 5568
rect 38016 5525 38025 5559
rect 38025 5525 38059 5559
rect 38059 5525 38068 5559
rect 38016 5516 38068 5525
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 19064 5312 19116 5364
rect 37832 5312 37884 5364
rect 38384 5355 38436 5364
rect 38384 5321 38393 5355
rect 38393 5321 38427 5355
rect 38427 5321 38436 5355
rect 38384 5312 38436 5321
rect 18144 5244 18196 5296
rect 8392 5176 8444 5228
rect 19524 5176 19576 5228
rect 19616 5219 19668 5228
rect 19616 5185 19625 5219
rect 19625 5185 19659 5219
rect 19659 5185 19668 5219
rect 19616 5176 19668 5185
rect 19708 5219 19760 5228
rect 19708 5185 19717 5219
rect 19717 5185 19751 5219
rect 19751 5185 19760 5219
rect 19708 5176 19760 5185
rect 22008 5176 22060 5228
rect 18236 5108 18288 5160
rect 7564 5040 7616 5092
rect 19432 5040 19484 5092
rect 19524 5040 19576 5092
rect 19708 5040 19760 5092
rect 26884 5040 26936 5092
rect 1124 4972 1176 5024
rect 19340 4972 19392 5024
rect 35440 4972 35492 5024
rect 39120 4972 39172 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 38384 4743 38436 4752
rect 38384 4709 38393 4743
rect 38393 4709 38427 4743
rect 38427 4709 38436 4743
rect 38384 4700 38436 4709
rect 13728 4632 13780 4684
rect 26884 4632 26936 4684
rect 21180 4539 21232 4548
rect 21180 4505 21189 4539
rect 21189 4505 21223 4539
rect 21223 4505 21232 4539
rect 21180 4496 21232 4505
rect 26884 4428 26936 4480
rect 38016 4471 38068 4480
rect 38016 4437 38025 4471
rect 38025 4437 38059 4471
rect 38059 4437 38068 4471
rect 38016 4428 38068 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 5172 4088 5224 4140
rect 15384 4088 15436 4140
rect 15476 4131 15528 4140
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 3424 4020 3476 4072
rect 7840 3952 7892 4004
rect 15476 3952 15528 4004
rect 17132 4020 17184 4072
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 20444 4131 20496 4140
rect 20444 4097 20453 4131
rect 20453 4097 20487 4131
rect 20487 4097 20496 4131
rect 20444 4088 20496 4097
rect 21824 4131 21876 4140
rect 21824 4097 21833 4131
rect 21833 4097 21867 4131
rect 21867 4097 21876 4131
rect 21824 4088 21876 4097
rect 15108 3884 15160 3936
rect 22100 3952 22152 4004
rect 22468 3952 22520 4004
rect 26884 4156 26936 4208
rect 22652 4131 22704 4140
rect 22652 4097 22661 4131
rect 22661 4097 22695 4131
rect 22695 4097 22704 4131
rect 22652 4088 22704 4097
rect 23112 4088 23164 4140
rect 33784 4088 33836 4140
rect 37464 3952 37516 4004
rect 38384 3995 38436 4004
rect 38384 3961 38393 3995
rect 38393 3961 38427 3995
rect 38427 3961 38436 3995
rect 38384 3952 38436 3961
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 16396 3927 16448 3936
rect 16396 3893 16405 3927
rect 16405 3893 16439 3927
rect 16439 3893 16448 3927
rect 16396 3884 16448 3893
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 17224 3927 17276 3936
rect 17224 3893 17233 3927
rect 17233 3893 17267 3927
rect 17267 3893 17276 3927
rect 17224 3884 17276 3893
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 18880 3927 18932 3936
rect 18880 3893 18889 3927
rect 18889 3893 18923 3927
rect 18923 3893 18932 3927
rect 18880 3884 18932 3893
rect 19616 3927 19668 3936
rect 19616 3893 19625 3927
rect 19625 3893 19659 3927
rect 19659 3893 19668 3927
rect 19616 3884 19668 3893
rect 20628 3927 20680 3936
rect 20628 3893 20637 3927
rect 20637 3893 20671 3927
rect 20671 3893 20680 3927
rect 20628 3884 20680 3893
rect 20904 3884 20956 3936
rect 21548 3927 21600 3936
rect 21548 3893 21557 3927
rect 21557 3893 21591 3927
rect 21591 3893 21600 3927
rect 21548 3884 21600 3893
rect 21824 3884 21876 3936
rect 22192 3927 22244 3936
rect 22192 3893 22201 3927
rect 22201 3893 22235 3927
rect 22235 3893 22244 3927
rect 22192 3884 22244 3893
rect 22560 3927 22612 3936
rect 22560 3893 22569 3927
rect 22569 3893 22603 3927
rect 22603 3893 22612 3927
rect 22560 3884 22612 3893
rect 27068 3884 27120 3936
rect 27436 3884 27488 3936
rect 39120 3884 39172 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 8852 3680 8904 3732
rect 17132 3680 17184 3732
rect 23020 3680 23072 3732
rect 9588 3612 9640 3664
rect 18236 3612 18288 3664
rect 22284 3612 22336 3664
rect 37832 3680 37884 3732
rect 26424 3612 26476 3664
rect 32404 3612 32456 3664
rect 38384 3655 38436 3664
rect 38384 3621 38393 3655
rect 38393 3621 38427 3655
rect 38427 3621 38436 3655
rect 38384 3612 38436 3621
rect 8576 3544 8628 3596
rect 17408 3544 17460 3596
rect 18052 3544 18104 3596
rect 1492 3476 1544 3528
rect 20352 3476 20404 3528
rect 27068 3544 27120 3596
rect 26976 3519 27028 3528
rect 26976 3485 26985 3519
rect 26985 3485 27019 3519
rect 27019 3485 27028 3519
rect 26976 3476 27028 3485
rect 9496 3408 9548 3460
rect 16396 3408 16448 3460
rect 23480 3408 23532 3460
rect 38200 3519 38252 3528
rect 38200 3485 38209 3519
rect 38209 3485 38243 3519
rect 38243 3485 38252 3519
rect 38200 3476 38252 3485
rect 22100 3383 22152 3392
rect 22100 3349 22109 3383
rect 22109 3349 22143 3383
rect 22143 3349 22152 3383
rect 22100 3340 22152 3349
rect 25228 3383 25280 3392
rect 25228 3349 25237 3383
rect 25237 3349 25271 3383
rect 25271 3349 25280 3383
rect 25228 3340 25280 3349
rect 25596 3383 25648 3392
rect 25596 3349 25605 3383
rect 25605 3349 25639 3383
rect 25639 3349 25648 3383
rect 25596 3340 25648 3349
rect 26332 3383 26384 3392
rect 26332 3349 26341 3383
rect 26341 3349 26375 3383
rect 26375 3349 26384 3383
rect 26332 3340 26384 3349
rect 26516 3383 26568 3392
rect 26516 3349 26525 3383
rect 26525 3349 26559 3383
rect 26559 3349 26568 3383
rect 26516 3340 26568 3349
rect 27528 3340 27580 3392
rect 38016 3383 38068 3392
rect 38016 3349 38025 3383
rect 38025 3349 38059 3383
rect 38059 3349 38068 3383
rect 38016 3340 38068 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 17224 3136 17276 3188
rect 38200 3136 38252 3188
rect 38384 3179 38436 3188
rect 38384 3145 38393 3179
rect 38393 3145 38427 3179
rect 38427 3145 38436 3179
rect 38384 3136 38436 3145
rect 7012 3068 7064 3120
rect 20444 3068 20496 3120
rect 22468 3068 22520 3120
rect 16304 3000 16356 3052
rect 24676 3000 24728 3052
rect 19616 2932 19668 2984
rect 26240 3000 26292 3052
rect 26332 3000 26384 3052
rect 34520 3000 34572 3052
rect 37464 3043 37516 3052
rect 37464 3009 37473 3043
rect 37473 3009 37507 3043
rect 37507 3009 37516 3043
rect 37464 3000 37516 3009
rect 37832 3043 37884 3052
rect 37832 3009 37841 3043
rect 37841 3009 37875 3043
rect 37875 3009 37884 3043
rect 37832 3000 37884 3009
rect 25596 2932 25648 2984
rect 31852 2932 31904 2984
rect 20628 2864 20680 2916
rect 32680 2864 32732 2916
rect 26240 2796 26292 2848
rect 33508 2796 33560 2848
rect 37832 2796 37884 2848
rect 39120 2796 39172 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 18880 2592 18932 2644
rect 36360 2592 36412 2644
rect 17776 2524 17828 2576
rect 23664 2524 23716 2576
rect 16856 2456 16908 2508
rect 36636 2567 36688 2576
rect 36636 2533 36645 2567
rect 36645 2533 36679 2567
rect 36679 2533 36688 2567
rect 36636 2524 36688 2533
rect 37004 2567 37056 2576
rect 37004 2533 37013 2567
rect 37013 2533 37047 2567
rect 37047 2533 37056 2567
rect 37004 2524 37056 2533
rect 38384 2567 38436 2576
rect 38384 2533 38393 2567
rect 38393 2533 38427 2567
rect 38427 2533 38436 2567
rect 38384 2524 38436 2533
rect 15660 2388 15712 2440
rect 23664 2388 23716 2440
rect 36360 2388 36412 2440
rect 38200 2431 38252 2440
rect 38200 2397 38209 2431
rect 38209 2397 38243 2431
rect 38243 2397 38252 2431
rect 38200 2388 38252 2397
rect 22560 2252 22612 2304
rect 34980 2252 35032 2304
rect 37648 2295 37700 2304
rect 37648 2261 37657 2295
rect 37657 2261 37691 2295
rect 37691 2261 37700 2295
rect 37648 2252 37700 2261
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 14372 2048 14424 2100
rect 23480 2048 23532 2100
rect 34980 2048 35032 2100
rect 38200 2048 38252 2100
rect 19892 1504 19944 1556
rect 23112 1504 23164 1556
<< metal2 >>
rect 2778 11096 2834 11152
rect 3054 11096 3110 11152
rect 3330 11096 3386 11152
rect 3606 11096 3662 11152
rect 3882 11096 3938 11152
rect 4158 11096 4214 11152
rect 4434 11096 4490 11152
rect 4710 11096 4766 11152
rect 4986 11096 5042 11152
rect 5262 11096 5318 11152
rect 5538 11096 5594 11152
rect 5814 11096 5870 11152
rect 6090 11096 6146 11152
rect 6366 11096 6422 11152
rect 6642 11096 6698 11152
rect 6918 11096 6974 11152
rect 7194 11096 7250 11152
rect 7470 11096 7526 11152
rect 7746 11096 7802 11152
rect 8022 11096 8078 11152
rect 8298 11096 8354 11152
rect 8574 11096 8630 11152
rect 8850 11096 8906 11152
rect 9126 11096 9182 11152
rect 9402 11096 9458 11152
rect 9678 11096 9734 11152
rect 9954 11096 10010 11152
rect 10230 11096 10286 11152
rect 10322 11112 10378 11121
rect 570 10024 626 10033
rect 570 9959 626 9968
rect 584 9081 612 9959
rect 938 9888 994 9897
rect 938 9823 994 9832
rect 570 9072 626 9081
rect 570 9007 626 9016
rect 952 8809 980 9823
rect 1308 9716 1360 9722
rect 1308 9658 1360 9664
rect 1124 9172 1176 9178
rect 1124 9114 1176 9120
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 1136 7993 1164 9114
rect 1320 8537 1348 9658
rect 2792 8634 2820 11096
rect 3068 9194 3096 11096
rect 2884 9166 3096 9194
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 1306 8528 1362 8537
rect 1306 8463 1362 8472
rect 1306 8392 1362 8401
rect 1216 8356 1268 8362
rect 1306 8327 1362 8336
rect 1674 8392 1730 8401
rect 1674 8327 1676 8336
rect 1216 8298 1268 8304
rect 1122 7984 1178 7993
rect 1122 7919 1178 7928
rect 1228 7177 1256 8298
rect 1320 7721 1348 8327
rect 1728 8327 1730 8336
rect 1676 8298 1728 8304
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2884 8090 2912 9166
rect 3344 8786 3372 11096
rect 3344 8758 3464 8786
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3436 8634 3464 8758
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3620 8090 3648 11096
rect 3896 8362 3924 11096
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 4172 8090 4200 11096
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 4264 8498 4292 8842
rect 4448 8634 4476 11096
rect 4724 8634 4752 11096
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4908 8498 4936 8774
rect 5000 8634 5028 11096
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 4080 7546 4108 7822
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 1214 7168 1270 7177
rect 1214 7103 1270 7112
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1766 6760 1822 6769
rect 1766 6695 1822 6704
rect 1780 6089 1808 6695
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 4356 6118 4384 8434
rect 5276 8090 5304 11096
rect 5552 8634 5580 11096
rect 5828 8634 5856 11096
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5368 7546 5396 8366
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5460 6662 5488 8434
rect 5552 7546 5580 8434
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5644 7410 5672 7958
rect 5828 7478 5856 8230
rect 6104 8090 6132 11096
rect 6274 9480 6330 9489
rect 6274 9415 6330 9424
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6288 7993 6316 9415
rect 6380 8634 6408 11096
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6274 7984 6330 7993
rect 6274 7919 6330 7928
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6012 7546 6040 7822
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6104 7546 6132 7754
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 6196 7410 6224 7754
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6380 7274 6408 8298
rect 6472 7478 6500 8774
rect 6656 8090 6684 11096
rect 6932 8634 6960 11096
rect 7208 8634 7236 11096
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 4344 6112 4396 6118
rect 1766 6080 1822 6089
rect 4344 6054 4396 6060
rect 1766 6015 1822 6024
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 6472 5642 6500 6734
rect 6748 6730 6776 7890
rect 6840 7562 6868 8502
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6920 7880 6972 7886
rect 6972 7828 7144 7834
rect 6920 7822 7144 7828
rect 6932 7806 7144 7822
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6840 7546 6960 7562
rect 6840 7540 6972 7546
rect 6840 7534 6920 7540
rect 6920 7482 6972 7488
rect 7024 7410 7052 7686
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6932 7206 6960 7346
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 7116 6254 7144 7806
rect 7208 6458 7236 8434
rect 7300 6866 7328 8434
rect 7392 7206 7420 10950
rect 7484 8090 7512 11096
rect 7760 8634 7788 11096
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7392 6186 7420 6734
rect 7576 6662 7604 8366
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7668 6610 7696 8434
rect 7852 7274 7880 8910
rect 8036 8634 8064 11096
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8312 8090 8340 11096
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8404 8498 8432 9046
rect 8484 8628 8536 8634
rect 8588 8616 8616 11096
rect 8864 9602 8892 11096
rect 8772 9574 8892 9602
rect 8772 8634 8800 9574
rect 9140 9466 9168 11096
rect 8864 9438 9168 9466
rect 8536 8588 8616 8616
rect 8760 8628 8812 8634
rect 8484 8570 8536 8576
rect 8760 8570 8812 8576
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8864 8090 8892 9438
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 9416 8634 9444 11096
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9508 8498 9536 8774
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 8312 7002 8340 7822
rect 8496 7002 8524 7890
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9508 7478 9536 7822
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 7748 6656 7800 6662
rect 7668 6604 7748 6610
rect 7668 6598 7800 6604
rect 7668 6582 7788 6598
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7852 5914 7880 6734
rect 8772 6322 8800 6734
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9416 6458 9444 6598
rect 9600 6458 9628 8298
rect 9692 8090 9720 11096
rect 9770 10976 9826 10985
rect 9770 10911 9826 10920
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9784 6798 9812 10911
rect 9862 10160 9918 10169
rect 9862 10095 9918 10104
rect 9876 8294 9904 10095
rect 9968 8634 9996 11096
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 10152 8106 10180 8842
rect 10244 8634 10272 11096
rect 10506 11096 10562 11152
rect 10782 11096 10838 11152
rect 11058 11096 11114 11152
rect 11334 11096 11390 11152
rect 11610 11096 11666 11152
rect 11886 11096 11942 11152
rect 12162 11096 12218 11152
rect 12438 11096 12494 11152
rect 12714 11096 12770 11152
rect 12990 11096 13046 11152
rect 13266 11096 13322 11152
rect 13542 11096 13598 11152
rect 13818 11096 13874 11152
rect 14094 11096 14150 11152
rect 14370 11096 14426 11152
rect 14646 11096 14702 11152
rect 14922 11096 14978 11152
rect 15198 11096 15254 11152
rect 15474 11096 15530 11152
rect 15750 11096 15806 11152
rect 16026 11096 16082 11152
rect 16302 11096 16358 11152
rect 16578 11096 16634 11152
rect 16854 11096 16910 11152
rect 17130 11096 17186 11152
rect 17406 11096 17462 11152
rect 17682 11096 17738 11152
rect 17958 11096 18014 11152
rect 18234 11096 18290 11152
rect 18510 11096 18566 11152
rect 18786 11096 18842 11152
rect 19062 11096 19118 11152
rect 19338 11096 19394 11152
rect 19614 11096 19670 11152
rect 19890 11096 19946 11152
rect 20166 11096 20222 11152
rect 20442 11096 20498 11152
rect 20718 11096 20774 11152
rect 20994 11098 21050 11152
rect 20916 11096 21050 11098
rect 21270 11096 21326 11152
rect 21546 11096 21602 11152
rect 21822 11112 21878 11152
rect 10322 11047 10378 11056
rect 10416 11076 10468 11082
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10152 8078 10272 8106
rect 10138 7984 10194 7993
rect 10138 7919 10194 7928
rect 10048 7880 10100 7886
rect 9954 7848 10010 7857
rect 10048 7822 10100 7828
rect 9954 7783 10010 7792
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9968 6322 9996 7783
rect 10060 7546 10088 7822
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10152 7410 10180 7919
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10244 6662 10272 8078
rect 10336 6798 10364 11047
rect 10416 11018 10468 11024
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8312 5846 8340 6258
rect 10232 6248 10284 6254
rect 8390 6216 8446 6225
rect 8390 6151 8446 6160
rect 10046 6216 10102 6225
rect 10336 6236 10364 6394
rect 10428 6322 10456 11018
rect 10520 8634 10548 11096
rect 10692 9308 10744 9314
rect 10692 9250 10744 9256
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10704 8566 10732 9250
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10612 6798 10640 8434
rect 10796 8090 10824 11096
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10980 6322 11008 11018
rect 11072 8634 11100 11096
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 7206 11100 8230
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11164 6866 11192 7822
rect 11256 7274 11284 8434
rect 11348 8090 11376 11096
rect 11428 10940 11480 10946
rect 11428 10882 11480 10888
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10284 6208 10364 6236
rect 10232 6190 10284 6196
rect 10046 6151 10048 6160
rect 8300 5840 8352 5846
rect 7562 5808 7618 5817
rect 8300 5782 8352 5788
rect 7562 5743 7618 5752
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 1122 5536 1178 5545
rect 1122 5471 1178 5480
rect 1136 5030 1164 5471
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 7576 5098 7604 5743
rect 8404 5234 8432 6151
rect 10100 6151 10102 6160
rect 10048 6122 10100 6128
rect 10428 6118 10456 6258
rect 10506 6216 10562 6225
rect 10506 6151 10562 6160
rect 10520 6118 10548 6151
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 11072 5681 11100 6802
rect 11440 6662 11468 10882
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11532 5914 11560 10746
rect 11624 8634 11652 11096
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11716 6458 11744 7822
rect 11808 6662 11836 8434
rect 11900 8090 11928 11096
rect 11980 9240 12032 9246
rect 11980 9182 12032 9188
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11992 7818 12020 9182
rect 12176 8634 12204 11096
rect 12452 8634 12480 11096
rect 12728 8634 12756 11096
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12820 8498 12848 8842
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 12268 7002 12296 7822
rect 12636 7342 12664 8230
rect 13004 8090 13032 11096
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13188 8498 13216 8978
rect 13280 8634 13308 11096
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 13188 6866 13216 8298
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 12728 6254 12756 6666
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 13004 5778 13032 6734
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13280 5710 13308 6734
rect 13268 5704 13320 5710
rect 11058 5672 11114 5681
rect 13268 5646 13320 5652
rect 13372 5642 13400 9930
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13464 7274 13492 8366
rect 13556 8090 13584 11096
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13648 7750 13676 9862
rect 13832 8362 13860 11096
rect 13912 9784 13964 9790
rect 13912 9726 13964 9732
rect 13924 9246 13952 9726
rect 13912 9240 13964 9246
rect 13912 9182 13964 9188
rect 14108 8634 14136 11096
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14200 8430 14228 9386
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13740 7528 13768 7822
rect 13740 7500 13860 7528
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13740 7002 13768 7346
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13556 6225 13584 6734
rect 13542 6216 13598 6225
rect 13832 6186 13860 7500
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14292 6882 14320 8502
rect 14384 8090 14412 11096
rect 14464 10872 14516 10878
rect 14464 10814 14516 10820
rect 14476 8412 14504 10814
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14568 8514 14596 9522
rect 14660 8634 14688 11096
rect 14738 9072 14794 9081
rect 14738 9007 14794 9016
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14568 8486 14688 8514
rect 14476 8384 14596 8412
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14568 7426 14596 8384
rect 14660 8022 14688 8486
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14476 7398 14596 7426
rect 14384 7206 14412 7346
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14200 6854 14320 6882
rect 14200 6662 14228 6854
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 13542 6151 13598 6160
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 11058 5607 11114 5616
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 14292 5574 14320 6734
rect 14476 6730 14504 7398
rect 14660 7206 14688 7822
rect 14752 7410 14780 9007
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14844 7546 14872 8774
rect 14936 8634 14964 11096
rect 15212 9466 15240 11096
rect 15212 9438 15424 9466
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15396 8090 15424 9438
rect 15488 8634 15516 11096
rect 15660 9240 15712 9246
rect 15660 9182 15712 9188
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15580 7834 15608 8978
rect 15672 8498 15700 9182
rect 15764 8634 15792 11096
rect 15844 9308 15896 9314
rect 15844 9250 15896 9256
rect 15936 9308 15988 9314
rect 15936 9250 15988 9256
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15580 7806 15700 7834
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 15580 7410 15608 7686
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 15672 6497 15700 7806
rect 15856 7546 15884 9250
rect 15948 8498 15976 9250
rect 16040 8634 16068 11096
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16132 8498 16160 9318
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15658 6488 15714 6497
rect 15658 6423 15714 6432
rect 16132 5817 16160 8298
rect 16224 7857 16252 8978
rect 16316 8634 16344 11096
rect 16486 10840 16542 10849
rect 16486 10775 16542 10784
rect 16394 8936 16450 8945
rect 16394 8871 16450 8880
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16210 7848 16266 7857
rect 16210 7783 16266 7792
rect 16210 7304 16266 7313
rect 16210 7239 16266 7248
rect 16224 6361 16252 7239
rect 16316 6633 16344 8434
rect 16408 7274 16436 8871
rect 16500 7410 16528 10775
rect 16592 8362 16620 11096
rect 16672 9852 16724 9858
rect 16672 9794 16724 9800
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16684 7478 16712 9794
rect 16868 8634 16896 11096
rect 17144 10169 17172 11096
rect 17130 10160 17186 10169
rect 17130 10095 17186 10104
rect 17420 9586 17448 11096
rect 17696 9926 17724 11096
rect 17972 11014 18000 11096
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16776 7546 16804 7890
rect 17052 7546 17080 9046
rect 18248 8974 18276 11096
rect 18524 9994 18552 11096
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 18800 9790 18828 11096
rect 18788 9784 18840 9790
rect 18788 9726 18840 9732
rect 18236 8968 18288 8974
rect 17512 8894 17724 8922
rect 18236 8910 18288 8916
rect 17512 8498 17540 8894
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17222 7848 17278 7857
rect 17222 7783 17278 7792
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 17236 7410 17264 7783
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16302 6624 16358 6633
rect 16302 6559 16358 6568
rect 16868 6458 17356 6474
rect 16856 6452 17368 6458
rect 16908 6446 17316 6452
rect 16856 6394 16908 6400
rect 17316 6394 17368 6400
rect 16210 6352 16266 6361
rect 16210 6287 16266 6296
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 16118 5808 16174 5817
rect 16118 5743 16174 5752
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 16776 5137 16804 6258
rect 17236 6225 17264 6258
rect 17222 6216 17278 6225
rect 17222 6151 17278 6160
rect 17604 5846 17632 8774
rect 17696 8634 17724 8894
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17788 8090 17816 8230
rect 19076 8090 19104 11096
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19352 7993 19380 11096
rect 19628 8838 19656 11096
rect 19904 9042 19932 11096
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 20180 8922 20208 11096
rect 20350 9344 20406 9353
rect 20350 9279 20406 9288
rect 19812 8894 20208 8922
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19706 8256 19762 8265
rect 19706 8191 19762 8200
rect 19338 7984 19394 7993
rect 19338 7919 19394 7928
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17696 5914 17724 7142
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17592 5840 17644 5846
rect 17592 5782 17644 5788
rect 17788 5273 17816 6598
rect 17880 6225 17908 6734
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 17866 6216 17922 6225
rect 17866 6151 17922 6160
rect 18156 5302 18184 6598
rect 18432 6390 18460 7754
rect 19524 7472 19576 7478
rect 19338 7440 19394 7449
rect 19338 7375 19394 7384
rect 19522 7440 19524 7449
rect 19576 7440 19578 7449
rect 19720 7410 19748 8191
rect 19522 7375 19578 7384
rect 19708 7404 19760 7410
rect 19352 7274 19380 7375
rect 19708 7346 19760 7352
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18708 6769 18736 7142
rect 18694 6760 18750 6769
rect 18694 6695 18750 6704
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18144 5296 18196 5302
rect 17774 5264 17830 5273
rect 18144 5238 18196 5244
rect 17774 5199 17830 5208
rect 18248 5166 18276 6326
rect 19076 5370 19104 7142
rect 19246 6896 19302 6905
rect 19246 6831 19302 6840
rect 19260 6730 19288 6831
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18236 5160 18288 5166
rect 16762 5128 16818 5137
rect 7564 5092 7616 5098
rect 18236 5102 18288 5108
rect 16762 5063 16818 5072
rect 7564 5034 7616 5040
rect 19352 5030 19380 6598
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19444 5098 19472 5578
rect 19536 5234 19564 6598
rect 19812 6254 19840 8894
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20364 7410 20392 9279
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 19996 7313 20024 7346
rect 19982 7304 20038 7313
rect 19982 7239 20038 7248
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 20456 6118 20484 11096
rect 20732 10810 20760 11096
rect 20916 11070 21036 11096
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20810 9208 20866 9217
rect 20810 9143 20866 9152
rect 20718 8256 20774 8265
rect 20718 8191 20774 8200
rect 20732 7342 20760 8191
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20824 7002 20852 9143
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20916 6882 20944 11070
rect 21284 10985 21312 11096
rect 21270 10976 21326 10985
rect 21560 10946 21588 11096
rect 22098 11098 22154 11152
rect 22098 11096 22232 11098
rect 22374 11096 22430 11152
rect 22650 11096 22706 11152
rect 22926 11098 22982 11152
rect 22848 11096 22982 11098
rect 23202 11096 23258 11152
rect 23478 11096 23534 11152
rect 23754 11096 23810 11152
rect 24030 11096 24086 11152
rect 24306 11096 24362 11152
rect 24582 11096 24638 11152
rect 24858 11096 24914 11152
rect 25134 11096 25190 11152
rect 25410 11096 25466 11152
rect 25686 11096 25742 11152
rect 25962 11096 26018 11152
rect 26238 11096 26294 11152
rect 26514 11096 26570 11152
rect 26790 11096 26846 11152
rect 27066 11098 27122 11152
rect 26896 11096 27122 11098
rect 27342 11096 27398 11152
rect 27618 11098 27674 11152
rect 27618 11096 27752 11098
rect 27894 11096 27950 11152
rect 28170 11096 28226 11152
rect 28446 11096 28502 11152
rect 28722 11096 28778 11152
rect 28998 11096 29054 11152
rect 29274 11096 29330 11152
rect 29550 11096 29606 11152
rect 29826 11096 29882 11152
rect 30102 11096 30158 11152
rect 30378 11096 30434 11152
rect 30654 11096 30710 11152
rect 30930 11096 30986 11152
rect 31206 11096 31262 11152
rect 31482 11096 31538 11152
rect 31758 11096 31814 11152
rect 32034 11096 32090 11152
rect 32310 11096 32366 11152
rect 32586 11096 32642 11152
rect 32862 11096 32918 11152
rect 33138 11096 33194 11152
rect 33414 11096 33470 11152
rect 33690 11096 33746 11152
rect 33966 11096 34022 11152
rect 34242 11096 34298 11152
rect 34518 11096 34574 11152
rect 34794 11096 34850 11152
rect 35070 11096 35126 11152
rect 35346 11096 35402 11152
rect 35622 11096 35678 11152
rect 35898 11096 35954 11152
rect 36174 11096 36230 11152
rect 36450 11096 36506 11152
rect 36726 11096 36782 11152
rect 37002 11096 37058 11152
rect 22112 11082 22232 11096
rect 22112 11076 22244 11082
rect 22112 11070 22192 11076
rect 21822 11047 21878 11056
rect 22192 11018 22244 11024
rect 22388 11014 22416 11096
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 21270 10911 21326 10920
rect 21548 10940 21600 10946
rect 21548 10882 21600 10888
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21362 9888 21418 9897
rect 21362 9823 21418 9832
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 21008 6905 21036 7482
rect 21376 7410 21404 9823
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21468 6934 21496 7142
rect 21456 6928 21508 6934
rect 20824 6854 20944 6882
rect 20994 6896 21050 6905
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20824 5681 20852 6854
rect 21456 6870 21508 6876
rect 20994 6831 21050 6840
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 21560 6322 21588 10066
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21836 7410 21864 9658
rect 22466 9480 22522 9489
rect 22466 9415 22522 9424
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22008 7812 22060 7818
rect 22008 7754 22060 7760
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 22020 7206 22048 7754
rect 22112 7410 22140 9114
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22190 8528 22246 8537
rect 22190 8463 22246 8472
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22204 6866 22232 8463
rect 22296 7546 22324 8910
rect 22480 7546 22508 9415
rect 22664 9081 22692 11096
rect 22848 11070 22968 11096
rect 22650 9072 22706 9081
rect 22650 9007 22706 9016
rect 22742 8392 22798 8401
rect 22742 8327 22798 8336
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22756 6866 22784 8327
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22112 6746 22140 6802
rect 22112 6718 22324 6746
rect 22100 6656 22152 6662
rect 22152 6604 22232 6610
rect 22100 6598 22232 6604
rect 22112 6582 22232 6598
rect 22204 6458 22232 6582
rect 22296 6497 22324 6718
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22282 6488 22338 6497
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22192 6452 22244 6458
rect 22282 6423 22338 6432
rect 22192 6394 22244 6400
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 20810 5672 20866 5681
rect 21652 5642 21680 6258
rect 22112 6254 22140 6394
rect 22572 6254 22600 6598
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22480 5778 22508 6054
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 20810 5607 20866 5616
rect 21640 5636 21692 5642
rect 21640 5578 21692 5584
rect 22848 5574 22876 11070
rect 23216 10878 23244 11096
rect 23204 10872 23256 10878
rect 23204 10814 23256 10820
rect 23388 10192 23440 10198
rect 23388 10134 23440 10140
rect 22926 9752 22982 9761
rect 22926 9687 22982 9696
rect 22940 7410 22968 9687
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19616 5228 19668 5234
rect 19708 5228 19760 5234
rect 19668 5188 19708 5216
rect 19616 5170 19668 5176
rect 22008 5228 22060 5234
rect 19760 5188 19840 5216
rect 19708 5170 19760 5176
rect 19432 5092 19484 5098
rect 19432 5034 19484 5040
rect 19524 5092 19576 5098
rect 19708 5092 19760 5098
rect 19576 5052 19708 5080
rect 19524 5034 19576 5040
rect 19708 5034 19760 5040
rect 1124 5024 1176 5030
rect 1124 4966 1176 4972
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 19812 4729 19840 5188
rect 22008 5170 22060 5176
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19798 4720 19854 4729
rect 13728 4684 13780 4690
rect 19798 4655 19854 4664
rect 13728 4626 13780 4632
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 13740 4185 13768 4626
rect 21178 4584 21234 4593
rect 21178 4519 21180 4528
rect 21232 4519 21234 4528
rect 21180 4490 21232 4496
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 13726 4176 13782 4185
rect 5172 4140 5224 4146
rect 13726 4111 13782 4120
rect 15384 4140 15436 4146
rect 5172 4082 5224 4088
rect 15384 4082 15436 4088
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1504 56 1532 3470
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 3436 1986 3464 4014
rect 3344 1958 3464 1986
rect 3344 56 3372 1958
rect 5184 56 5212 4082
rect 15396 4049 15424 4082
rect 15382 4040 15438 4049
rect 7840 4004 7892 4010
rect 15488 4010 15516 4082
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 15382 3975 15438 3984
rect 15476 4004 15528 4010
rect 7840 3946 7892 3952
rect 15476 3946 15528 3952
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 7024 56 7052 3062
rect 7852 1193 7880 3946
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8588 1465 8616 3538
rect 8574 1456 8630 1465
rect 8574 1391 8630 1400
rect 7838 1184 7894 1193
rect 7838 1119 7894 1128
rect 8864 56 8892 3674
rect 9588 3664 9640 3670
rect 15120 3641 15148 3878
rect 9588 3606 9640 3612
rect 15106 3632 15162 3641
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 9508 2417 9536 3402
rect 9494 2408 9550 2417
rect 9494 2343 9550 2352
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9600 1737 9628 3606
rect 15106 3567 15162 3576
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 15672 2446 15700 3878
rect 16210 3360 16266 3369
rect 16210 3295 16266 3304
rect 15660 2440 15712 2446
rect 10690 2408 10746 2417
rect 15660 2382 15712 2388
rect 10690 2343 10746 2352
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 10704 56 10732 2343
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 14372 2100 14424 2106
rect 14372 2042 14424 2048
rect 12530 1864 12586 1873
rect 12530 1799 12586 1808
rect 12544 56 12572 1799
rect 14384 56 14412 2042
rect 16224 56 16252 3295
rect 16316 3058 16344 3878
rect 16408 3466 16436 3878
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16868 2514 16896 3878
rect 17144 3738 17172 4014
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 17236 3194 17264 3878
rect 17420 3602 17448 3878
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17788 2582 17816 3878
rect 18248 3670 18276 3878
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 18064 56 18092 3538
rect 18708 2009 18736 4082
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 18892 2650 18920 3878
rect 19628 2990 19656 3878
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20350 3632 20406 3641
rect 20350 3567 20406 3576
rect 20364 3534 20392 3567
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20456 3126 20484 4082
rect 21836 3942 21864 4082
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 20444 3120 20496 3126
rect 20444 3062 20496 3068
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 20640 2922 20668 3878
rect 20916 3097 20944 3878
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 20902 3088 20958 3097
rect 20902 3023 20958 3032
rect 21560 2961 21588 3878
rect 21546 2952 21602 2961
rect 20628 2916 20680 2922
rect 21546 2887 21602 2896
rect 20628 2858 20680 2864
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 18694 2000 18750 2009
rect 18694 1935 18750 1944
rect 19892 1556 19944 1562
rect 19892 1498 19944 1504
rect 19904 56 19932 1498
rect 21744 56 21864 82
rect 1490 0 1546 56
rect 3330 0 3386 56
rect 5170 0 5226 56
rect 7010 0 7066 56
rect 8850 0 8906 56
rect 10690 0 10746 56
rect 12530 0 12586 56
rect 14370 0 14426 56
rect 16210 0 16266 56
rect 18050 0 18106 56
rect 19890 0 19946 56
rect 21730 54 21864 56
rect 21730 0 21786 54
rect 21836 42 21864 54
rect 22020 42 22048 5170
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22112 4010 22324 4026
rect 22100 4004 22324 4010
rect 22152 3998 22324 4004
rect 22100 3946 22152 3952
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22098 3496 22154 3505
rect 22098 3431 22154 3440
rect 22112 3398 22140 3431
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22204 2553 22232 3878
rect 22296 3670 22324 3998
rect 22468 4004 22520 4010
rect 22468 3946 22520 3952
rect 22284 3664 22336 3670
rect 22284 3606 22336 3612
rect 22480 3126 22508 3946
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 22190 2544 22246 2553
rect 22190 2479 22246 2488
rect 22572 2310 22600 3878
rect 22664 3777 22692 4082
rect 22650 3768 22706 3777
rect 23032 3738 23060 8434
rect 23400 7750 23428 10134
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23386 7304 23442 7313
rect 23386 7239 23388 7248
rect 23440 7239 23442 7248
rect 23388 7210 23440 7216
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 23124 5574 23152 6598
rect 23492 5846 23520 11096
rect 23768 6322 23796 11096
rect 24044 9217 24072 11096
rect 24030 9208 24086 9217
rect 24030 9143 24086 9152
rect 24216 8900 24268 8906
rect 24216 8842 24268 8848
rect 24228 7274 24256 8842
rect 24216 7268 24268 7274
rect 24216 7210 24268 7216
rect 23848 6860 23900 6866
rect 23848 6802 23900 6808
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23860 5914 23888 6802
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23480 5840 23532 5846
rect 23480 5782 23532 5788
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 22650 3703 22706 3712
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 23124 1562 23152 4082
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 23492 2106 23520 3402
rect 23480 2100 23532 2106
rect 23480 2042 23532 2048
rect 23112 1556 23164 1562
rect 23112 1498 23164 1504
rect 23584 56 23612 5646
rect 24320 5642 24348 11096
rect 24596 10130 24624 11096
rect 24584 10124 24636 10130
rect 24584 10066 24636 10072
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 24688 3058 24716 9046
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24780 5846 24808 7142
rect 24872 6225 24900 11096
rect 25148 8265 25176 11096
rect 25424 8945 25452 11096
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 25410 8936 25466 8945
rect 25410 8871 25466 8880
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25134 8256 25190 8265
rect 25134 8191 25190 8200
rect 25424 6746 25452 8570
rect 25608 6798 25636 9862
rect 25700 9858 25728 11096
rect 25976 10198 26004 11096
rect 26252 10849 26280 11096
rect 26238 10840 26294 10849
rect 26238 10775 26294 10784
rect 25964 10192 26016 10198
rect 25964 10134 26016 10140
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 25688 9852 25740 9858
rect 25688 9794 25740 9800
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25700 6798 25728 9658
rect 25792 6866 25820 9658
rect 25884 7410 25912 9998
rect 26148 8424 26200 8430
rect 26424 8424 26476 8430
rect 26200 8372 26372 8378
rect 26148 8366 26372 8372
rect 26424 8366 26476 8372
rect 26160 8350 26372 8366
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 26148 6928 26200 6934
rect 25976 6876 26148 6882
rect 25976 6870 26200 6876
rect 25780 6860 25832 6866
rect 25780 6802 25832 6808
rect 25976 6854 26188 6870
rect 26344 6866 26372 8350
rect 26332 6860 26384 6866
rect 25596 6792 25648 6798
rect 25424 6718 25544 6746
rect 25596 6734 25648 6740
rect 25688 6792 25740 6798
rect 25688 6734 25740 6740
rect 25516 6662 25544 6718
rect 25412 6656 25464 6662
rect 25412 6598 25464 6604
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 24858 6216 24914 6225
rect 25424 6186 25452 6598
rect 25976 6361 26004 6854
rect 26332 6802 26384 6808
rect 26056 6724 26108 6730
rect 26056 6666 26108 6672
rect 25962 6352 26018 6361
rect 25504 6316 25556 6322
rect 25962 6287 26018 6296
rect 25504 6258 25556 6264
rect 24858 6151 24914 6160
rect 25412 6180 25464 6186
rect 25412 6122 25464 6128
rect 24768 5840 24820 5846
rect 24768 5782 24820 5788
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 24676 3052 24728 3058
rect 24676 2994 24728 3000
rect 23664 2576 23716 2582
rect 23664 2518 23716 2524
rect 23676 2446 23704 2518
rect 23664 2440 23716 2446
rect 25240 2417 25268 3334
rect 25516 2774 25544 6258
rect 26068 6118 26096 6666
rect 26056 6112 26108 6118
rect 26056 6054 26108 6060
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 26436 3670 26464 8366
rect 26528 7857 26556 11096
rect 26608 9444 26660 9450
rect 26608 9386 26660 9392
rect 26514 7848 26570 7857
rect 26514 7783 26570 7792
rect 26620 6662 26648 9386
rect 26804 9330 26832 11096
rect 26712 9302 26832 9330
rect 26896 11070 27108 11096
rect 26712 7449 26740 9302
rect 26792 7472 26844 7478
rect 26698 7440 26754 7449
rect 26792 7414 26844 7420
rect 26698 7375 26754 7384
rect 26804 7274 26832 7414
rect 26792 7268 26844 7274
rect 26792 7210 26844 7216
rect 26896 6798 26924 11070
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 27356 7426 27384 11096
rect 27632 11070 27752 11096
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27264 7398 27384 7426
rect 27264 6798 27292 7398
rect 26884 6792 26936 6798
rect 26884 6734 26936 6740
rect 27252 6792 27304 6798
rect 27448 6746 27476 9114
rect 27724 8362 27752 11070
rect 27712 8356 27764 8362
rect 27712 8298 27764 8304
rect 27908 7410 27936 11096
rect 28184 9353 28212 11096
rect 28170 9344 28226 9353
rect 28170 9279 28226 9288
rect 28460 9217 28488 11096
rect 28736 9489 28764 11096
rect 28722 9480 28778 9489
rect 28722 9415 28778 9424
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28446 9208 28502 9217
rect 28446 9143 28502 9152
rect 28448 9036 28500 9042
rect 28448 8978 28500 8984
rect 27988 8560 28040 8566
rect 27988 8502 28040 8508
rect 27896 7404 27948 7410
rect 27896 7346 27948 7352
rect 27526 7168 27582 7177
rect 27526 7103 27582 7112
rect 27252 6734 27304 6740
rect 27356 6718 27476 6746
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27356 5794 27384 6718
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 27448 5953 27476 6598
rect 27434 5944 27490 5953
rect 27434 5879 27490 5888
rect 27356 5766 27476 5794
rect 27250 5672 27306 5681
rect 27306 5630 27384 5658
rect 27250 5607 27306 5616
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 26884 5092 26936 5098
rect 26884 5034 26936 5040
rect 26896 4690 26924 5034
rect 26884 4684 26936 4690
rect 26884 4626 26936 4632
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 26896 4214 26924 4422
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 26884 4208 26936 4214
rect 26884 4150 26936 4156
rect 27068 3936 27120 3942
rect 27068 3878 27120 3884
rect 26424 3664 26476 3670
rect 26424 3606 26476 3612
rect 26974 3632 27030 3641
rect 27080 3602 27108 3878
rect 26974 3567 27030 3576
rect 27068 3596 27120 3602
rect 26988 3534 27016 3567
rect 27068 3538 27120 3544
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 25596 3392 25648 3398
rect 25596 3334 25648 3340
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26516 3392 26568 3398
rect 26516 3334 26568 3340
rect 25608 2990 25636 3334
rect 26344 3058 26372 3334
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 25596 2984 25648 2990
rect 25596 2926 25648 2932
rect 26252 2854 26280 2994
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 25424 2746 25544 2774
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 23664 2382 23716 2388
rect 25226 2408 25282 2417
rect 25226 2343 25282 2352
rect 25424 56 25452 2746
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26528 1873 26556 3334
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 26514 1864 26570 1873
rect 26514 1799 26570 1808
rect 27356 1442 27384 5630
rect 27448 3942 27476 5766
rect 27436 3936 27488 3942
rect 27436 3878 27488 3884
rect 27540 3398 27568 7103
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 27632 6186 27660 6734
rect 27896 6656 27948 6662
rect 27896 6598 27948 6604
rect 27908 6390 27936 6598
rect 28000 6474 28028 8502
rect 28356 8356 28408 8362
rect 28356 8298 28408 8304
rect 28264 6928 28316 6934
rect 28264 6870 28316 6876
rect 28080 6656 28132 6662
rect 28276 6644 28304 6870
rect 28368 6798 28396 8298
rect 28356 6792 28408 6798
rect 28356 6734 28408 6740
rect 28132 6616 28304 6644
rect 28356 6656 28408 6662
rect 28080 6598 28132 6604
rect 28356 6598 28408 6604
rect 28368 6474 28396 6598
rect 28000 6446 28396 6474
rect 28460 6458 28488 8978
rect 28828 7546 28856 9318
rect 28908 9308 28960 9314
rect 28908 9250 28960 9256
rect 28816 7540 28868 7546
rect 28816 7482 28868 7488
rect 28920 7206 28948 9250
rect 29012 8090 29040 11096
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 29288 6798 29316 11096
rect 29458 9344 29514 9353
rect 29458 9279 29514 9288
rect 29368 9240 29420 9246
rect 29368 9182 29420 9188
rect 29380 7206 29408 9182
rect 29472 7410 29500 9279
rect 29460 7404 29512 7410
rect 29460 7346 29512 7352
rect 29368 7200 29420 7206
rect 29368 7142 29420 7148
rect 29276 6792 29328 6798
rect 28538 6760 28594 6769
rect 29276 6734 29328 6740
rect 29564 6730 29592 11096
rect 29734 9208 29790 9217
rect 29734 9143 29790 9152
rect 29644 8288 29696 8294
rect 29644 8230 29696 8236
rect 29656 7206 29684 8230
rect 29748 7410 29776 9143
rect 29736 7404 29788 7410
rect 29736 7346 29788 7352
rect 29644 7200 29696 7206
rect 29644 7142 29696 7148
rect 29840 6866 29868 11096
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 29932 7410 29960 8026
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 29920 7404 29972 7410
rect 29920 7346 29972 7352
rect 30024 7206 30052 7822
rect 30012 7200 30064 7206
rect 30012 7142 30064 7148
rect 29828 6860 29880 6866
rect 29828 6802 29880 6808
rect 28538 6695 28594 6704
rect 29552 6724 29604 6730
rect 28552 6662 28580 6695
rect 29552 6666 29604 6672
rect 28540 6656 28592 6662
rect 28540 6598 28592 6604
rect 28448 6452 28500 6458
rect 28448 6394 28500 6400
rect 27896 6384 27948 6390
rect 27896 6326 27948 6332
rect 29276 6316 29328 6322
rect 29276 6258 29328 6264
rect 27620 6180 27672 6186
rect 27620 6122 27672 6128
rect 29092 5704 29144 5710
rect 29288 5681 29316 6258
rect 29460 6248 29512 6254
rect 29460 6190 29512 6196
rect 29472 5914 29500 6190
rect 30116 6186 30144 11096
rect 30392 9790 30420 11096
rect 30380 9784 30432 9790
rect 30380 9726 30432 9732
rect 30668 9722 30696 11096
rect 30944 9926 30972 11096
rect 31220 10062 31248 11096
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 30932 9920 30984 9926
rect 30932 9862 30984 9868
rect 30656 9716 30708 9722
rect 30656 9658 30708 9664
rect 30286 9480 30342 9489
rect 30286 9415 30342 9424
rect 30300 7410 30328 9415
rect 31496 8634 31524 11096
rect 31772 8634 31800 11096
rect 31852 8900 31904 8906
rect 31852 8842 31904 8848
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31760 8628 31812 8634
rect 31760 8570 31812 8576
rect 31760 7744 31812 7750
rect 31760 7686 31812 7692
rect 30288 7404 30340 7410
rect 30288 7346 30340 7352
rect 31772 7177 31800 7686
rect 31758 7168 31814 7177
rect 31758 7103 31814 7112
rect 30104 6180 30156 6186
rect 30104 6122 30156 6128
rect 29460 5908 29512 5914
rect 29460 5850 29512 5856
rect 29092 5646 29144 5652
rect 29274 5672 29330 5681
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 27264 1414 27384 1442
rect 27264 56 27292 1414
rect 29104 56 29132 5646
rect 29274 5607 29330 5616
rect 30932 5636 30984 5642
rect 30932 5578 30984 5584
rect 30944 56 30972 5578
rect 31864 2990 31892 8842
rect 32048 8362 32076 11096
rect 32128 9104 32180 9110
rect 32128 9046 32180 9052
rect 32140 8498 32168 9046
rect 32324 8616 32352 11096
rect 32404 8628 32456 8634
rect 32324 8588 32404 8616
rect 32404 8570 32456 8576
rect 32600 8566 32628 11096
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 32128 8492 32180 8498
rect 32128 8434 32180 8440
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32036 8356 32088 8362
rect 32036 8298 32088 8304
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 32416 3670 32444 7822
rect 32508 4049 32536 8434
rect 32494 4040 32550 4049
rect 32494 3975 32550 3984
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 31852 2984 31904 2990
rect 31852 2926 31904 2932
rect 32692 2922 32720 8434
rect 32876 8362 32904 11096
rect 33152 8838 33180 11096
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 32864 8356 32916 8362
rect 32864 8298 32916 8304
rect 32956 8288 33008 8294
rect 32956 8230 33008 8236
rect 32772 7948 32824 7954
rect 32772 7890 32824 7896
rect 32784 5846 32812 7890
rect 32968 7834 32996 8230
rect 33428 8090 33456 11096
rect 33600 8900 33652 8906
rect 33600 8842 33652 8848
rect 33612 8498 33640 8842
rect 33508 8492 33560 8498
rect 33508 8434 33560 8440
rect 33600 8492 33652 8498
rect 33600 8434 33652 8440
rect 33416 8084 33468 8090
rect 33416 8026 33468 8032
rect 32876 7806 32996 7834
rect 32876 5914 32904 7806
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 32864 5908 32916 5914
rect 32864 5850 32916 5856
rect 32772 5840 32824 5846
rect 32772 5782 32824 5788
rect 32772 5636 32824 5642
rect 32772 5578 32824 5584
rect 32680 2916 32732 2922
rect 32680 2858 32732 2864
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32784 56 32812 5578
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 33520 2854 33548 8434
rect 33704 8106 33732 11096
rect 33980 8634 34008 11096
rect 34152 8832 34204 8838
rect 34152 8774 34204 8780
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 34164 8362 34192 8774
rect 34256 8362 34284 11096
rect 34532 8430 34560 11096
rect 34612 8492 34664 8498
rect 34612 8434 34664 8440
rect 34520 8424 34572 8430
rect 34520 8366 34572 8372
rect 34152 8356 34204 8362
rect 34152 8298 34204 8304
rect 34244 8356 34296 8362
rect 34244 8298 34296 8304
rect 33704 8090 33824 8106
rect 33704 8084 33836 8090
rect 33704 8078 33784 8084
rect 33784 8026 33836 8032
rect 33784 7812 33836 7818
rect 33784 7754 33836 7760
rect 33796 7478 33824 7754
rect 33784 7472 33836 7478
rect 33784 7414 33836 7420
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 34256 6118 34284 7346
rect 34244 6112 34296 6118
rect 34244 6054 34296 6060
rect 34624 5794 34652 8434
rect 34808 8090 34836 11096
rect 34888 9172 34940 9178
rect 34888 9114 34940 9120
rect 34900 8498 34928 9114
rect 35084 8634 35112 11096
rect 35360 8838 35388 11096
rect 35348 8832 35400 8838
rect 35348 8774 35400 8780
rect 35072 8628 35124 8634
rect 35072 8570 35124 8576
rect 35636 8498 35664 11096
rect 35808 9036 35860 9042
rect 35808 8978 35860 8984
rect 35716 8832 35768 8838
rect 35716 8774 35768 8780
rect 34888 8492 34940 8498
rect 34888 8434 34940 8440
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35624 8492 35676 8498
rect 35624 8434 35676 8440
rect 34796 8084 34848 8090
rect 34796 8026 34848 8032
rect 34980 7948 35032 7954
rect 34980 7890 35032 7896
rect 34992 7274 35020 7890
rect 35072 7880 35124 7886
rect 35072 7822 35124 7828
rect 34980 7268 35032 7274
rect 34980 7210 35032 7216
rect 34704 7200 34756 7206
rect 34704 7142 34756 7148
rect 34532 5766 34652 5794
rect 33784 4140 33836 4146
rect 33784 4082 33836 4088
rect 33796 3505 33824 4082
rect 33782 3496 33838 3505
rect 33782 3431 33838 3440
rect 34532 3058 34560 5766
rect 34612 5636 34664 5642
rect 34612 5578 34664 5584
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 33508 2848 33560 2854
rect 33508 2790 33560 2796
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 34624 56 34652 5578
rect 34716 5574 34744 7142
rect 34978 6896 35034 6905
rect 34978 6831 34980 6840
rect 35032 6831 35034 6840
rect 34980 6802 35032 6808
rect 34794 6352 34850 6361
rect 34794 6287 34850 6296
rect 34808 5574 34836 6287
rect 35084 5846 35112 7822
rect 35164 7812 35216 7818
rect 35164 7754 35216 7760
rect 35176 6322 35204 7754
rect 35164 6316 35216 6322
rect 35164 6258 35216 6264
rect 35072 5840 35124 5846
rect 35072 5782 35124 5788
rect 34704 5568 34756 5574
rect 34704 5510 34756 5516
rect 34796 5568 34848 5574
rect 34796 5510 34848 5516
rect 35452 5030 35480 8434
rect 35728 8362 35756 8774
rect 35820 8498 35848 8978
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35716 8356 35768 8362
rect 35716 8298 35768 8304
rect 35912 8090 35940 11096
rect 35992 8492 36044 8498
rect 35992 8434 36044 8440
rect 35900 8084 35952 8090
rect 35900 8026 35952 8032
rect 36004 6458 36032 8434
rect 36188 8106 36216 11096
rect 36464 8634 36492 11096
rect 36452 8628 36504 8634
rect 36452 8570 36504 8576
rect 36740 8566 36768 11096
rect 36910 8800 36966 8809
rect 36910 8735 36966 8744
rect 36728 8560 36780 8566
rect 36728 8502 36780 8508
rect 36188 8090 36308 8106
rect 36924 8090 36952 8735
rect 37016 8090 37044 11096
rect 38566 9616 38622 9625
rect 38566 9551 38622 9560
rect 37646 9344 37702 9353
rect 37646 9279 37702 9288
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 37372 8492 37424 8498
rect 37372 8434 37424 8440
rect 36188 8084 36320 8090
rect 36188 8078 36268 8084
rect 36268 8026 36320 8032
rect 36912 8084 36964 8090
rect 36912 8026 36964 8032
rect 37004 8084 37056 8090
rect 37004 8026 37056 8032
rect 36360 7880 36412 7886
rect 36360 7822 36412 7828
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 37096 7880 37148 7886
rect 37096 7822 37148 7828
rect 35992 6452 36044 6458
rect 35992 6394 36044 6400
rect 36372 5914 36400 7822
rect 36740 7002 36768 7822
rect 37004 7268 37056 7274
rect 37004 7210 37056 7216
rect 36728 6996 36780 7002
rect 36728 6938 36780 6944
rect 37016 6905 37044 7210
rect 37002 6896 37058 6905
rect 37002 6831 37058 6840
rect 36912 6112 36964 6118
rect 36912 6054 36964 6060
rect 36360 5908 36412 5914
rect 36360 5850 36412 5856
rect 36924 5710 36952 6054
rect 37108 5914 37136 7822
rect 37096 5908 37148 5914
rect 37096 5850 37148 5856
rect 37292 5846 37320 8434
rect 37384 5914 37412 8434
rect 37464 7880 37516 7886
rect 37464 7822 37516 7828
rect 37476 7546 37504 7822
rect 37660 7546 37688 9279
rect 38474 9072 38530 9081
rect 38474 9007 38530 9016
rect 38200 8968 38252 8974
rect 38200 8910 38252 8916
rect 38212 8498 38240 8910
rect 38290 8528 38346 8537
rect 38200 8492 38252 8498
rect 38290 8463 38346 8472
rect 38200 8434 38252 8440
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 38016 7744 38068 7750
rect 38016 7686 38068 7692
rect 37464 7540 37516 7546
rect 37464 7482 37516 7488
rect 37648 7540 37700 7546
rect 37648 7482 37700 7488
rect 38028 7449 38056 7686
rect 38304 7546 38332 8463
rect 38384 8356 38436 8362
rect 38384 8298 38436 8304
rect 38396 7993 38424 8298
rect 38382 7984 38438 7993
rect 38382 7919 38438 7928
rect 38384 7744 38436 7750
rect 38382 7712 38384 7721
rect 38436 7712 38438 7721
rect 38382 7647 38438 7656
rect 38292 7540 38344 7546
rect 38292 7482 38344 7488
rect 38014 7440 38070 7449
rect 38014 7375 38070 7384
rect 37738 7304 37794 7313
rect 37738 7239 37794 7248
rect 37464 6792 37516 6798
rect 37464 6734 37516 6740
rect 37556 6792 37608 6798
rect 37556 6734 37608 6740
rect 37476 6390 37504 6734
rect 37464 6384 37516 6390
rect 37464 6326 37516 6332
rect 37568 6254 37596 6734
rect 37648 6656 37700 6662
rect 37648 6598 37700 6604
rect 37660 6361 37688 6598
rect 37752 6390 37780 7239
rect 38384 7200 38436 7206
rect 38382 7168 38384 7177
rect 38436 7168 38438 7177
rect 37950 7100 38258 7109
rect 38382 7103 38438 7112
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38488 6662 38516 9007
rect 38580 6730 38608 9551
rect 38658 8256 38714 8265
rect 38658 8191 38714 8200
rect 38672 8090 38700 8191
rect 38660 8084 38712 8090
rect 38660 8026 38712 8032
rect 38568 6724 38620 6730
rect 38568 6666 38620 6672
rect 38476 6656 38528 6662
rect 38382 6624 38438 6633
rect 38476 6598 38528 6604
rect 38382 6559 38438 6568
rect 38396 6458 38424 6559
rect 38384 6452 38436 6458
rect 38384 6394 38436 6400
rect 37740 6384 37792 6390
rect 37646 6352 37702 6361
rect 37740 6326 37792 6332
rect 37646 6287 37702 6296
rect 37832 6316 37884 6322
rect 37832 6258 37884 6264
rect 37556 6248 37608 6254
rect 37556 6190 37608 6196
rect 37372 5908 37424 5914
rect 37372 5850 37424 5856
rect 37280 5840 37332 5846
rect 37280 5782 37332 5788
rect 36912 5704 36964 5710
rect 36912 5646 36964 5652
rect 36452 5636 36504 5642
rect 36452 5578 36504 5584
rect 35440 5024 35492 5030
rect 35440 4966 35492 4972
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 36372 2446 36400 2586
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 34980 2304 35032 2310
rect 34980 2246 35032 2252
rect 34992 2106 35020 2246
rect 34980 2100 35032 2106
rect 34980 2042 35032 2048
rect 36464 56 36492 5578
rect 37844 5370 37872 6258
rect 39580 6180 39632 6186
rect 39580 6122 39632 6128
rect 38292 6112 38344 6118
rect 39592 6089 39620 6122
rect 38292 6054 38344 6060
rect 39578 6080 39634 6089
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 38016 5568 38068 5574
rect 38014 5536 38016 5545
rect 38068 5536 38070 5545
rect 38014 5471 38070 5480
rect 37832 5364 37884 5370
rect 37832 5306 37884 5312
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 38016 4480 38068 4486
rect 38014 4448 38016 4457
rect 38068 4448 38070 4457
rect 38014 4383 38070 4392
rect 37464 4004 37516 4010
rect 37464 3946 37516 3952
rect 37476 3058 37504 3946
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 37832 3732 37884 3738
rect 37832 3674 37884 3680
rect 37844 3058 37872 3674
rect 38200 3528 38252 3534
rect 38200 3470 38252 3476
rect 38016 3392 38068 3398
rect 38014 3360 38016 3369
rect 38068 3360 38070 3369
rect 38014 3295 38070 3304
rect 38212 3194 38240 3470
rect 38200 3188 38252 3194
rect 38200 3130 38252 3136
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 37832 3052 37884 3058
rect 37832 2994 37884 3000
rect 37832 2848 37884 2854
rect 37832 2790 37884 2796
rect 36636 2576 36688 2582
rect 36636 2518 36688 2524
rect 37004 2576 37056 2582
rect 37004 2518 37056 2524
rect 36648 2009 36676 2518
rect 36634 2000 36690 2009
rect 36634 1935 36690 1944
rect 37016 1465 37044 2518
rect 37648 2304 37700 2310
rect 37648 2246 37700 2252
rect 37002 1456 37058 1465
rect 37002 1391 37058 1400
rect 37660 1193 37688 2246
rect 37844 1737 37872 2790
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38200 2440 38252 2446
rect 38200 2382 38252 2388
rect 38016 2304 38068 2310
rect 38014 2272 38016 2281
rect 38068 2272 38070 2281
rect 38014 2207 38070 2216
rect 38212 2106 38240 2382
rect 38200 2100 38252 2106
rect 38200 2042 38252 2048
rect 37830 1728 37886 1737
rect 37830 1663 37886 1672
rect 37646 1184 37702 1193
rect 37646 1119 37702 1128
rect 38304 56 38332 6054
rect 39578 6015 39634 6024
rect 38384 5840 38436 5846
rect 38382 5808 38384 5817
rect 38436 5808 38438 5817
rect 38382 5743 38438 5752
rect 38384 5364 38436 5370
rect 38384 5306 38436 5312
rect 38396 5273 38424 5306
rect 38382 5264 38438 5273
rect 38382 5199 38438 5208
rect 39120 5024 39172 5030
rect 39118 4992 39120 5001
rect 39172 4992 39174 5001
rect 39118 4927 39174 4936
rect 38384 4752 38436 4758
rect 38382 4720 38384 4729
rect 38436 4720 38438 4729
rect 38382 4655 38438 4664
rect 38382 4176 38438 4185
rect 38382 4111 38438 4120
rect 38396 4010 38424 4111
rect 38384 4004 38436 4010
rect 38384 3946 38436 3952
rect 39120 3936 39172 3942
rect 39118 3904 39120 3913
rect 39172 3904 39174 3913
rect 39118 3839 39174 3848
rect 38384 3664 38436 3670
rect 38382 3632 38384 3641
rect 38436 3632 38438 3641
rect 38382 3567 38438 3576
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38396 3097 38424 3130
rect 38382 3088 38438 3097
rect 38382 3023 38438 3032
rect 39120 2848 39172 2854
rect 39118 2816 39120 2825
rect 39172 2816 39174 2825
rect 39118 2751 39174 2760
rect 38384 2576 38436 2582
rect 38382 2544 38384 2553
rect 38436 2544 38438 2553
rect 38382 2479 38438 2488
rect 21836 14 22048 42
rect 23570 0 23626 56
rect 25410 0 25466 56
rect 27250 0 27306 56
rect 29090 0 29146 56
rect 30930 0 30986 56
rect 32770 0 32826 56
rect 34610 0 34666 56
rect 36450 0 36506 56
rect 38290 0 38346 56
<< via2 >>
rect 570 9968 626 10024
rect 938 9832 994 9888
rect 570 9016 626 9072
rect 938 8744 994 8800
rect 1306 8472 1362 8528
rect 1306 8336 1362 8392
rect 1674 8356 1730 8392
rect 1674 8336 1676 8356
rect 1676 8336 1728 8356
rect 1728 8336 1730 8356
rect 1122 7928 1178 7984
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 1306 7656 1362 7712
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 1214 7112 1270 7168
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1766 6704 1822 6760
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 6274 9424 6330 9480
rect 6274 7928 6330 7984
rect 1766 6024 1822 6080
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9770 10920 9826 10976
rect 9862 10104 9918 10160
rect 10322 11056 10378 11112
rect 10138 7928 10194 7984
rect 9954 7792 10010 7848
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 8390 6160 8446 6216
rect 10046 6180 10102 6216
rect 10046 6160 10048 6180
rect 10048 6160 10100 6180
rect 10100 6160 10102 6180
rect 7562 5752 7618 5808
rect 1122 5480 1178 5536
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 10506 6160 10562 6216
rect 11058 5616 11114 5672
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 13542 6160 13598 6216
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 14738 9016 14794 9072
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 15658 6432 15714 6488
rect 16486 10784 16542 10840
rect 16394 8880 16450 8936
rect 16210 7792 16266 7848
rect 16210 7248 16266 7304
rect 17130 10104 17186 10160
rect 17222 7792 17278 7848
rect 16302 6568 16358 6624
rect 16210 6296 16266 6352
rect 16118 5752 16174 5808
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 17222 6160 17278 6216
rect 20350 9288 20406 9344
rect 19706 8200 19762 8256
rect 19338 7928 19394 7984
rect 17866 6160 17922 6216
rect 19338 7384 19394 7440
rect 19522 7420 19524 7440
rect 19524 7420 19576 7440
rect 19576 7420 19578 7440
rect 19522 7384 19578 7420
rect 18694 6704 18750 6760
rect 17774 5208 17830 5264
rect 19246 6840 19302 6896
rect 16762 5072 16818 5128
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19982 7248 20038 7304
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 20810 9152 20866 9208
rect 20718 8200 20774 8256
rect 21270 10920 21326 10976
rect 21822 11056 21878 11112
rect 21362 9832 21418 9888
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 20994 6840 21050 6896
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 22466 9424 22522 9480
rect 22190 8472 22246 8528
rect 22650 9016 22706 9072
rect 22742 8336 22798 8392
rect 22282 6432 22338 6488
rect 20810 5616 20866 5672
rect 22926 9696 22982 9752
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19798 4664 19854 4720
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 21178 4548 21234 4584
rect 21178 4528 21180 4548
rect 21180 4528 21232 4548
rect 21232 4528 21234 4548
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 13726 4120 13782 4176
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 15382 3984 15438 4040
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 8574 1400 8630 1456
rect 7838 1128 7894 1184
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9494 2352 9550 2408
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 15106 3576 15162 3632
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 16210 3304 16266 3360
rect 10690 2352 10746 2408
rect 9586 1672 9642 1728
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 12530 1808 12586 1864
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 20350 3576 20406 3632
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 20902 3032 20958 3088
rect 21546 2896 21602 2952
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 18694 1944 18750 2000
rect 22098 3440 22154 3496
rect 22190 2488 22246 2544
rect 22650 3712 22706 3768
rect 23386 7268 23442 7304
rect 23386 7248 23388 7268
rect 23388 7248 23440 7268
rect 23440 7248 23442 7268
rect 24030 9152 24086 9208
rect 25410 8880 25466 8936
rect 25134 8200 25190 8256
rect 26238 10784 26294 10840
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 24858 6160 24914 6216
rect 25962 6296 26018 6352
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 26514 7792 26570 7848
rect 26698 7384 26754 7440
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 28170 9288 28226 9344
rect 28722 9424 28778 9480
rect 28446 9152 28502 9208
rect 27526 7112 27582 7168
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27434 5888 27490 5944
rect 27250 5616 27306 5672
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 26974 3576 27030 3632
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25226 2352 25282 2408
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 26514 1808 26570 1864
rect 29458 9288 29514 9344
rect 28538 6704 28594 6760
rect 29734 9152 29790 9208
rect 30286 9424 30342 9480
rect 31758 7112 31814 7168
rect 29274 5616 29330 5672
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 32494 3984 32550 4040
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 33782 3440 33838 3496
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 34978 6860 35034 6896
rect 34978 6840 34980 6860
rect 34980 6840 35032 6860
rect 35032 6840 35034 6860
rect 34794 6296 34850 6352
rect 36910 8744 36966 8800
rect 38566 9560 38622 9616
rect 37646 9288 37702 9344
rect 37002 6840 37058 6896
rect 38474 9016 38530 9072
rect 38290 8472 38346 8528
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 38382 7928 38438 7984
rect 38382 7692 38384 7712
rect 38384 7692 38436 7712
rect 38436 7692 38438 7712
rect 38382 7656 38438 7692
rect 38014 7384 38070 7440
rect 37738 7248 37794 7304
rect 38382 7148 38384 7168
rect 38384 7148 38436 7168
rect 38436 7148 38438 7168
rect 38382 7112 38438 7148
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 38658 8200 38714 8256
rect 38382 6568 38438 6624
rect 37646 6296 37702 6352
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 38014 5516 38016 5536
rect 38016 5516 38068 5536
rect 38068 5516 38070 5536
rect 38014 5480 38070 5516
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 38014 4428 38016 4448
rect 38016 4428 38068 4448
rect 38068 4428 38070 4448
rect 38014 4392 38070 4428
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 38014 3340 38016 3360
rect 38016 3340 38068 3360
rect 38068 3340 38070 3360
rect 38014 3304 38070 3340
rect 36634 1944 36690 2000
rect 37002 1400 37058 1456
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 38014 2252 38016 2272
rect 38016 2252 38068 2272
rect 38068 2252 38070 2272
rect 38014 2216 38070 2252
rect 37830 1672 37886 1728
rect 37646 1128 37702 1184
rect 39578 6024 39634 6080
rect 38382 5788 38384 5808
rect 38384 5788 38436 5808
rect 38436 5788 38438 5808
rect 38382 5752 38438 5788
rect 38382 5208 38438 5264
rect 39118 4972 39120 4992
rect 39120 4972 39172 4992
rect 39172 4972 39174 4992
rect 39118 4936 39174 4972
rect 38382 4700 38384 4720
rect 38384 4700 38436 4720
rect 38436 4700 38438 4720
rect 38382 4664 38438 4700
rect 38382 4120 38438 4176
rect 39118 3884 39120 3904
rect 39120 3884 39172 3904
rect 39172 3884 39174 3904
rect 39118 3848 39174 3884
rect 38382 3612 38384 3632
rect 38384 3612 38436 3632
rect 38436 3612 38438 3632
rect 38382 3576 38438 3612
rect 38382 3032 38438 3088
rect 39118 2796 39120 2816
rect 39120 2796 39172 2816
rect 39172 2796 39174 2816
rect 39118 2760 39174 2796
rect 38382 2524 38384 2544
rect 38384 2524 38436 2544
rect 38436 2524 38438 2544
rect 38382 2488 38438 2524
<< metal3 >>
rect 10317 11114 10383 11117
rect 21817 11114 21883 11117
rect 10317 11112 21883 11114
rect 10317 11056 10322 11112
rect 10378 11056 21822 11112
rect 21878 11056 21883 11112
rect 10317 11054 21883 11056
rect 10317 11051 10383 11054
rect 21817 11051 21883 11054
rect 9765 10978 9831 10981
rect 21265 10978 21331 10981
rect 9765 10976 21331 10978
rect 9765 10920 9770 10976
rect 9826 10920 21270 10976
rect 21326 10920 21331 10976
rect 9765 10918 21331 10920
rect 9765 10915 9831 10918
rect 21265 10915 21331 10918
rect 16481 10842 16547 10845
rect 26233 10842 26299 10845
rect 16481 10840 26299 10842
rect 16481 10784 16486 10840
rect 16542 10784 26238 10840
rect 26294 10784 26299 10840
rect 16481 10782 26299 10784
rect 16481 10779 16547 10782
rect 26233 10779 26299 10782
rect 9857 10162 9923 10165
rect 17125 10162 17191 10165
rect 9857 10160 17191 10162
rect 9857 10104 9862 10160
rect 9918 10104 17130 10160
rect 17186 10104 17191 10160
rect 9857 10102 17191 10104
rect 9857 10099 9923 10102
rect 17125 10099 17191 10102
rect 565 10026 631 10029
rect 19374 10026 19380 10028
rect 565 10024 19380 10026
rect 565 9968 570 10024
rect 626 9968 19380 10024
rect 565 9966 19380 9968
rect 565 9963 631 9966
rect 19374 9964 19380 9966
rect 19444 9964 19450 10028
rect 933 9890 999 9893
rect 21357 9890 21423 9893
rect 933 9888 21423 9890
rect 933 9832 938 9888
rect 994 9832 21362 9888
rect 21418 9832 21423 9888
rect 933 9830 21423 9832
rect 933 9827 999 9830
rect 21357 9827 21423 9830
rect 22921 9754 22987 9757
rect 1350 9752 22987 9754
rect 1350 9696 22926 9752
rect 22982 9696 22987 9752
rect 1350 9694 22987 9696
rect 0 9618 120 9648
rect 1350 9618 1410 9694
rect 22921 9691 22987 9694
rect 0 9558 1410 9618
rect 38561 9618 38627 9621
rect 39808 9618 39928 9648
rect 38561 9616 39928 9618
rect 38561 9560 38566 9616
rect 38622 9560 39928 9616
rect 38561 9558 39928 9560
rect 0 9528 120 9558
rect 38561 9555 38627 9558
rect 39808 9528 39928 9558
rect 6269 9482 6335 9485
rect 22461 9482 22527 9485
rect 6269 9480 22527 9482
rect 6269 9424 6274 9480
rect 6330 9424 22466 9480
rect 22522 9424 22527 9480
rect 6269 9422 22527 9424
rect 6269 9419 6335 9422
rect 22461 9419 22527 9422
rect 28717 9482 28783 9485
rect 30281 9482 30347 9485
rect 28717 9480 30347 9482
rect 28717 9424 28722 9480
rect 28778 9424 30286 9480
rect 30342 9424 30347 9480
rect 28717 9422 30347 9424
rect 28717 9419 28783 9422
rect 30281 9419 30347 9422
rect 0 9346 120 9376
rect 20345 9346 20411 9349
rect 0 9344 20411 9346
rect 0 9288 20350 9344
rect 20406 9288 20411 9344
rect 0 9286 20411 9288
rect 0 9256 120 9286
rect 20345 9283 20411 9286
rect 28165 9346 28231 9349
rect 29453 9346 29519 9349
rect 28165 9344 29519 9346
rect 28165 9288 28170 9344
rect 28226 9288 29458 9344
rect 29514 9288 29519 9344
rect 28165 9286 29519 9288
rect 28165 9283 28231 9286
rect 29453 9283 29519 9286
rect 37641 9346 37707 9349
rect 39808 9346 39928 9376
rect 37641 9344 39928 9346
rect 37641 9288 37646 9344
rect 37702 9288 39928 9344
rect 37641 9286 39928 9288
rect 37641 9283 37707 9286
rect 39808 9256 39928 9286
rect 20805 9210 20871 9213
rect 24025 9210 24091 9213
rect 20805 9208 24091 9210
rect 20805 9152 20810 9208
rect 20866 9152 24030 9208
rect 24086 9152 24091 9208
rect 20805 9150 24091 9152
rect 20805 9147 20871 9150
rect 24025 9147 24091 9150
rect 28441 9210 28507 9213
rect 29729 9210 29795 9213
rect 28441 9208 29795 9210
rect 28441 9152 28446 9208
rect 28502 9152 29734 9208
rect 29790 9152 29795 9208
rect 28441 9150 29795 9152
rect 28441 9147 28507 9150
rect 29729 9147 29795 9150
rect 0 9074 120 9104
rect 565 9074 631 9077
rect 0 9072 631 9074
rect 0 9016 570 9072
rect 626 9016 631 9072
rect 0 9014 631 9016
rect 0 8984 120 9014
rect 565 9011 631 9014
rect 14733 9074 14799 9077
rect 22645 9074 22711 9077
rect 14733 9072 22711 9074
rect 14733 9016 14738 9072
rect 14794 9016 22650 9072
rect 22706 9016 22711 9072
rect 14733 9014 22711 9016
rect 14733 9011 14799 9014
rect 22645 9011 22711 9014
rect 38469 9074 38535 9077
rect 39808 9074 39928 9104
rect 38469 9072 39928 9074
rect 38469 9016 38474 9072
rect 38530 9016 39928 9072
rect 38469 9014 39928 9016
rect 38469 9011 38535 9014
rect 39808 8984 39928 9014
rect 16389 8938 16455 8941
rect 25405 8938 25471 8941
rect 16389 8936 25471 8938
rect 16389 8880 16394 8936
rect 16450 8880 25410 8936
rect 25466 8880 25471 8936
rect 16389 8878 25471 8880
rect 16389 8875 16455 8878
rect 25405 8875 25471 8878
rect 0 8802 120 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 120 8742
rect 933 8739 999 8742
rect 36905 8802 36971 8805
rect 39808 8802 39928 8832
rect 36905 8800 39928 8802
rect 36905 8744 36910 8800
rect 36966 8744 39928 8800
rect 36905 8742 39928 8744
rect 36905 8739 36971 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 39808 8712 39928 8742
rect 33006 8671 33322 8672
rect 0 8530 120 8560
rect 1301 8530 1367 8533
rect 22185 8530 22251 8533
rect 0 8528 1367 8530
rect 0 8472 1306 8528
rect 1362 8472 1367 8528
rect 0 8470 1367 8472
rect 0 8440 120 8470
rect 1301 8467 1367 8470
rect 1534 8528 22251 8530
rect 1534 8472 22190 8528
rect 22246 8472 22251 8528
rect 1534 8470 22251 8472
rect 1301 8394 1367 8397
rect 1534 8394 1594 8470
rect 22185 8467 22251 8470
rect 38285 8530 38351 8533
rect 39808 8530 39928 8560
rect 38285 8528 39928 8530
rect 38285 8472 38290 8528
rect 38346 8472 39928 8528
rect 38285 8470 39928 8472
rect 38285 8467 38351 8470
rect 39808 8440 39928 8470
rect 1301 8392 1594 8394
rect 1301 8336 1306 8392
rect 1362 8336 1594 8392
rect 1301 8334 1594 8336
rect 1669 8394 1735 8397
rect 22737 8394 22803 8397
rect 1669 8392 22803 8394
rect 1669 8336 1674 8392
rect 1730 8336 22742 8392
rect 22798 8336 22803 8392
rect 1669 8334 22803 8336
rect 1301 8331 1367 8334
rect 1669 8331 1735 8334
rect 22737 8331 22803 8334
rect 0 8258 120 8288
rect 0 8198 1824 8258
rect 0 8168 120 8198
rect 0 7986 120 8016
rect 1117 7986 1183 7989
rect 0 7984 1183 7986
rect 0 7928 1122 7984
rect 1178 7928 1183 7984
rect 0 7926 1183 7928
rect 1764 7986 1824 8198
rect 19374 8196 19380 8260
rect 19444 8258 19450 8260
rect 19701 8258 19767 8261
rect 19444 8256 19767 8258
rect 19444 8200 19706 8256
rect 19762 8200 19767 8256
rect 19444 8198 19767 8200
rect 19444 8196 19450 8198
rect 19701 8195 19767 8198
rect 20713 8258 20779 8261
rect 25129 8258 25195 8261
rect 20713 8256 25195 8258
rect 20713 8200 20718 8256
rect 20774 8200 25134 8256
rect 25190 8200 25195 8256
rect 20713 8198 25195 8200
rect 20713 8195 20779 8198
rect 25129 8195 25195 8198
rect 38653 8258 38719 8261
rect 39808 8258 39928 8288
rect 38653 8256 39928 8258
rect 38653 8200 38658 8256
rect 38714 8200 39928 8256
rect 38653 8198 39928 8200
rect 38653 8195 38719 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 39808 8168 39928 8198
rect 37946 8127 38262 8128
rect 6269 7986 6335 7989
rect 1764 7984 6335 7986
rect 1764 7928 6274 7984
rect 6330 7928 6335 7984
rect 1764 7926 6335 7928
rect 0 7896 120 7926
rect 1117 7923 1183 7926
rect 6269 7923 6335 7926
rect 10133 7986 10199 7989
rect 19333 7986 19399 7989
rect 10133 7984 19399 7986
rect 10133 7928 10138 7984
rect 10194 7928 19338 7984
rect 19394 7928 19399 7984
rect 10133 7926 19399 7928
rect 10133 7923 10199 7926
rect 19333 7923 19399 7926
rect 38377 7986 38443 7989
rect 39808 7986 39928 8016
rect 38377 7984 39928 7986
rect 38377 7928 38382 7984
rect 38438 7928 39928 7984
rect 38377 7926 39928 7928
rect 38377 7923 38443 7926
rect 39808 7896 39928 7926
rect 9949 7850 10015 7853
rect 16205 7850 16271 7853
rect 9949 7848 16271 7850
rect 9949 7792 9954 7848
rect 10010 7792 16210 7848
rect 16266 7792 16271 7848
rect 9949 7790 16271 7792
rect 9949 7787 10015 7790
rect 16205 7787 16271 7790
rect 17217 7850 17283 7853
rect 26509 7850 26575 7853
rect 17217 7848 26575 7850
rect 17217 7792 17222 7848
rect 17278 7792 26514 7848
rect 26570 7792 26575 7848
rect 17217 7790 26575 7792
rect 17217 7787 17283 7790
rect 26509 7787 26575 7790
rect 0 7714 120 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 120 7654
rect 1301 7651 1367 7654
rect 38377 7714 38443 7717
rect 39808 7714 39928 7744
rect 38377 7712 39928 7714
rect 38377 7656 38382 7712
rect 38438 7656 39928 7712
rect 38377 7654 39928 7656
rect 38377 7651 38443 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 39808 7624 39928 7654
rect 33006 7583 33322 7584
rect 0 7442 120 7472
rect 19333 7442 19399 7445
rect 0 7440 19399 7442
rect 0 7384 19338 7440
rect 19394 7384 19399 7440
rect 0 7382 19399 7384
rect 0 7352 120 7382
rect 19333 7379 19399 7382
rect 19517 7442 19583 7445
rect 26693 7442 26759 7445
rect 19517 7440 26759 7442
rect 19517 7384 19522 7440
rect 19578 7384 26698 7440
rect 26754 7384 26759 7440
rect 19517 7382 26759 7384
rect 19517 7379 19583 7382
rect 26693 7379 26759 7382
rect 38009 7442 38075 7445
rect 39808 7442 39928 7472
rect 38009 7440 39928 7442
rect 38009 7384 38014 7440
rect 38070 7384 39928 7440
rect 38009 7382 39928 7384
rect 38009 7379 38075 7382
rect 39808 7352 39928 7382
rect 16205 7306 16271 7309
rect 19977 7306 20043 7309
rect 16205 7304 20043 7306
rect 16205 7248 16210 7304
rect 16266 7248 19982 7304
rect 20038 7248 20043 7304
rect 16205 7246 20043 7248
rect 16205 7243 16271 7246
rect 19977 7243 20043 7246
rect 23381 7306 23447 7309
rect 37733 7306 37799 7309
rect 23381 7304 37799 7306
rect 23381 7248 23386 7304
rect 23442 7248 37738 7304
rect 37794 7248 37799 7304
rect 23381 7246 37799 7248
rect 23381 7243 23447 7246
rect 37733 7243 37799 7246
rect 0 7170 120 7200
rect 1209 7170 1275 7173
rect 0 7168 1275 7170
rect 0 7112 1214 7168
rect 1270 7112 1275 7168
rect 0 7110 1275 7112
rect 0 7080 120 7110
rect 1209 7107 1275 7110
rect 27521 7170 27587 7173
rect 31753 7170 31819 7173
rect 27521 7168 31819 7170
rect 27521 7112 27526 7168
rect 27582 7112 31758 7168
rect 31814 7112 31819 7168
rect 27521 7110 31819 7112
rect 27521 7107 27587 7110
rect 31753 7107 31819 7110
rect 38377 7170 38443 7173
rect 39808 7170 39928 7200
rect 38377 7168 39928 7170
rect 38377 7112 38382 7168
rect 38438 7112 39928 7168
rect 38377 7110 39928 7112
rect 38377 7107 38443 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 39808 7080 39928 7110
rect 37946 7039 38262 7040
rect 0 6898 120 6928
rect 19241 6898 19307 6901
rect 0 6896 19307 6898
rect 0 6840 19246 6896
rect 19302 6840 19307 6896
rect 0 6838 19307 6840
rect 0 6808 120 6838
rect 19241 6835 19307 6838
rect 20989 6898 21055 6901
rect 34973 6898 35039 6901
rect 20989 6896 35039 6898
rect 20989 6840 20994 6896
rect 21050 6840 34978 6896
rect 35034 6840 35039 6896
rect 20989 6838 35039 6840
rect 20989 6835 21055 6838
rect 34973 6835 35039 6838
rect 36997 6898 37063 6901
rect 39808 6898 39928 6928
rect 36997 6896 39928 6898
rect 36997 6840 37002 6896
rect 37058 6840 39928 6896
rect 36997 6838 39928 6840
rect 36997 6835 37063 6838
rect 39808 6808 39928 6838
rect 1761 6762 1827 6765
rect 18689 6762 18755 6765
rect 28533 6762 28599 6765
rect 1761 6760 18755 6762
rect 1761 6704 1766 6760
rect 1822 6704 18694 6760
rect 18750 6704 18755 6760
rect 1761 6702 18755 6704
rect 1761 6699 1827 6702
rect 18689 6699 18755 6702
rect 18830 6760 28599 6762
rect 18830 6704 28538 6760
rect 28594 6704 28599 6760
rect 18830 6702 28599 6704
rect 0 6626 120 6656
rect 16297 6626 16363 6629
rect 18830 6626 18890 6702
rect 28533 6699 28599 6702
rect 0 6566 2790 6626
rect 0 6536 120 6566
rect 0 6354 120 6384
rect 2730 6354 2790 6566
rect 16297 6624 18890 6626
rect 16297 6568 16302 6624
rect 16358 6568 18890 6624
rect 16297 6566 18890 6568
rect 38377 6626 38443 6629
rect 39808 6626 39928 6656
rect 38377 6624 39928 6626
rect 38377 6568 38382 6624
rect 38438 6568 39928 6624
rect 38377 6566 39928 6568
rect 16297 6563 16363 6566
rect 38377 6563 38443 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 39808 6536 39928 6566
rect 33006 6495 33322 6496
rect 15653 6490 15719 6493
rect 22277 6490 22343 6493
rect 15653 6488 17602 6490
rect 15653 6432 15658 6488
rect 15714 6432 17602 6488
rect 15653 6430 17602 6432
rect 15653 6427 15719 6430
rect 16205 6354 16271 6357
rect 0 6294 2330 6354
rect 2730 6352 16271 6354
rect 2730 6296 16210 6352
rect 16266 6296 16271 6352
rect 2730 6294 16271 6296
rect 17542 6354 17602 6430
rect 22277 6488 26250 6490
rect 22277 6432 22282 6488
rect 22338 6432 26250 6488
rect 22277 6430 26250 6432
rect 22277 6427 22343 6430
rect 25957 6354 26023 6357
rect 17542 6352 26023 6354
rect 17542 6296 25962 6352
rect 26018 6296 26023 6352
rect 17542 6294 26023 6296
rect 26190 6354 26250 6430
rect 34789 6354 34855 6357
rect 26190 6352 34855 6354
rect 26190 6296 34794 6352
rect 34850 6296 34855 6352
rect 26190 6294 34855 6296
rect 0 6264 120 6294
rect 2270 6218 2330 6294
rect 16205 6291 16271 6294
rect 25957 6291 26023 6294
rect 34789 6291 34855 6294
rect 37641 6354 37707 6357
rect 39808 6354 39928 6384
rect 37641 6352 39928 6354
rect 37641 6296 37646 6352
rect 37702 6296 39928 6352
rect 37641 6294 39928 6296
rect 37641 6291 37707 6294
rect 39808 6264 39928 6294
rect 8385 6218 8451 6221
rect 2270 6216 8451 6218
rect 2270 6160 8390 6216
rect 8446 6160 8451 6216
rect 2270 6158 8451 6160
rect 8385 6155 8451 6158
rect 10041 6218 10107 6221
rect 10501 6218 10567 6221
rect 10041 6216 10567 6218
rect 10041 6160 10046 6216
rect 10102 6160 10506 6216
rect 10562 6160 10567 6216
rect 10041 6158 10567 6160
rect 10041 6155 10107 6158
rect 10501 6155 10567 6158
rect 13537 6218 13603 6221
rect 17217 6218 17283 6221
rect 13537 6216 17283 6218
rect 13537 6160 13542 6216
rect 13598 6160 17222 6216
rect 17278 6160 17283 6216
rect 13537 6158 17283 6160
rect 13537 6155 13603 6158
rect 17217 6155 17283 6158
rect 17861 6218 17927 6221
rect 24853 6218 24919 6221
rect 17861 6216 24919 6218
rect 17861 6160 17866 6216
rect 17922 6160 24858 6216
rect 24914 6160 24919 6216
rect 17861 6158 24919 6160
rect 17861 6155 17927 6158
rect 24853 6155 24919 6158
rect 0 6082 120 6112
rect 1761 6082 1827 6085
rect 0 6080 1827 6082
rect 0 6024 1766 6080
rect 1822 6024 1827 6080
rect 0 6022 1827 6024
rect 0 5992 120 6022
rect 1761 6019 1827 6022
rect 39573 6082 39639 6085
rect 39808 6082 39928 6112
rect 39573 6080 39928 6082
rect 39573 6024 39578 6080
rect 39634 6024 39928 6080
rect 39573 6022 39928 6024
rect 39573 6019 39639 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 39808 5992 39928 6022
rect 37946 5951 38262 5952
rect 27429 5946 27495 5949
rect 26374 5944 27495 5946
rect 26374 5888 27434 5944
rect 27490 5888 27495 5944
rect 26374 5886 27495 5888
rect 0 5810 120 5840
rect 7557 5810 7623 5813
rect 0 5808 7623 5810
rect 0 5752 7562 5808
rect 7618 5752 7623 5808
rect 0 5750 7623 5752
rect 0 5720 120 5750
rect 7557 5747 7623 5750
rect 16113 5810 16179 5813
rect 26374 5810 26434 5886
rect 27429 5883 27495 5886
rect 16113 5808 26434 5810
rect 16113 5752 16118 5808
rect 16174 5752 26434 5808
rect 16113 5750 26434 5752
rect 38377 5810 38443 5813
rect 39808 5810 39928 5840
rect 38377 5808 39928 5810
rect 38377 5752 38382 5808
rect 38438 5752 39928 5808
rect 38377 5750 39928 5752
rect 16113 5747 16179 5750
rect 38377 5747 38443 5750
rect 39808 5720 39928 5750
rect 11053 5674 11119 5677
rect 20805 5674 20871 5677
rect 11053 5672 20871 5674
rect 11053 5616 11058 5672
rect 11114 5616 20810 5672
rect 20866 5616 20871 5672
rect 11053 5614 20871 5616
rect 11053 5611 11119 5614
rect 20805 5611 20871 5614
rect 27245 5674 27311 5677
rect 29269 5674 29335 5677
rect 27245 5672 29335 5674
rect 27245 5616 27250 5672
rect 27306 5616 29274 5672
rect 29330 5616 29335 5672
rect 27245 5614 29335 5616
rect 27245 5611 27311 5614
rect 29269 5611 29335 5614
rect 0 5538 120 5568
rect 1117 5538 1183 5541
rect 0 5536 1183 5538
rect 0 5480 1122 5536
rect 1178 5480 1183 5536
rect 0 5478 1183 5480
rect 0 5448 120 5478
rect 1117 5475 1183 5478
rect 38009 5538 38075 5541
rect 39808 5538 39928 5568
rect 38009 5536 39928 5538
rect 38009 5480 38014 5536
rect 38070 5480 39928 5536
rect 38009 5478 39928 5480
rect 38009 5475 38075 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 39808 5448 39928 5478
rect 33006 5407 33322 5408
rect 0 5266 120 5296
rect 17769 5266 17835 5269
rect 0 5264 17835 5266
rect 0 5208 17774 5264
rect 17830 5208 17835 5264
rect 0 5206 17835 5208
rect 0 5176 120 5206
rect 17769 5203 17835 5206
rect 38377 5266 38443 5269
rect 39808 5266 39928 5296
rect 38377 5264 39928 5266
rect 38377 5208 38382 5264
rect 38438 5208 39928 5264
rect 38377 5206 39928 5208
rect 38377 5203 38443 5206
rect 39808 5176 39928 5206
rect 16757 5130 16823 5133
rect 1718 5128 16823 5130
rect 1718 5072 16762 5128
rect 16818 5072 16823 5128
rect 1718 5070 16823 5072
rect 0 4994 120 5024
rect 1718 4994 1778 5070
rect 16757 5067 16823 5070
rect 0 4934 1778 4994
rect 39113 4994 39179 4997
rect 39808 4994 39928 5024
rect 39113 4992 39928 4994
rect 39113 4936 39118 4992
rect 39174 4936 39928 4992
rect 39113 4934 39928 4936
rect 0 4904 120 4934
rect 39113 4931 39179 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 39808 4904 39928 4934
rect 37946 4863 38262 4864
rect 0 4722 120 4752
rect 19793 4722 19859 4725
rect 0 4720 19859 4722
rect 0 4664 19798 4720
rect 19854 4664 19859 4720
rect 0 4662 19859 4664
rect 0 4632 120 4662
rect 19793 4659 19859 4662
rect 38377 4722 38443 4725
rect 39808 4722 39928 4752
rect 38377 4720 39928 4722
rect 38377 4664 38382 4720
rect 38438 4664 39928 4720
rect 38377 4662 39928 4664
rect 38377 4659 38443 4662
rect 39808 4632 39928 4662
rect 21173 4586 21239 4589
rect 2730 4584 21239 4586
rect 2730 4528 21178 4584
rect 21234 4528 21239 4584
rect 2730 4526 21239 4528
rect 0 4450 120 4480
rect 2730 4450 2790 4526
rect 21173 4523 21239 4526
rect 0 4390 2790 4450
rect 38009 4450 38075 4453
rect 39808 4450 39928 4480
rect 38009 4448 39928 4450
rect 38009 4392 38014 4448
rect 38070 4392 39928 4448
rect 38009 4390 39928 4392
rect 0 4360 120 4390
rect 38009 4387 38075 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 39808 4360 39928 4390
rect 33006 4319 33322 4320
rect 0 4178 120 4208
rect 13721 4178 13787 4181
rect 0 4176 13787 4178
rect 0 4120 13726 4176
rect 13782 4120 13787 4176
rect 0 4118 13787 4120
rect 0 4088 120 4118
rect 13721 4115 13787 4118
rect 38377 4178 38443 4181
rect 39808 4178 39928 4208
rect 38377 4176 39928 4178
rect 38377 4120 38382 4176
rect 38438 4120 39928 4176
rect 38377 4118 39928 4120
rect 38377 4115 38443 4118
rect 39808 4088 39928 4118
rect 15377 4042 15443 4045
rect 32489 4042 32555 4045
rect 1718 3982 15210 4042
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 0 3846 1778 3906
rect 0 3816 120 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 15150 3770 15210 3982
rect 15377 4040 32555 4042
rect 15377 3984 15382 4040
rect 15438 3984 32494 4040
rect 32550 3984 32555 4040
rect 15377 3982 32555 3984
rect 15377 3979 15443 3982
rect 32489 3979 32555 3982
rect 39113 3906 39179 3909
rect 39808 3906 39928 3936
rect 39113 3904 39928 3906
rect 39113 3848 39118 3904
rect 39174 3848 39928 3904
rect 39113 3846 39928 3848
rect 39113 3843 39179 3846
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 39808 3816 39928 3846
rect 37946 3775 38262 3776
rect 22645 3770 22711 3773
rect 15150 3710 18706 3770
rect 0 3634 120 3664
rect 15101 3634 15167 3637
rect 0 3632 15167 3634
rect 0 3576 15106 3632
rect 15162 3576 15167 3632
rect 0 3574 15167 3576
rect 18646 3634 18706 3710
rect 20486 3768 22711 3770
rect 20486 3712 22650 3768
rect 22706 3712 22711 3768
rect 20486 3710 22711 3712
rect 20345 3634 20411 3637
rect 18646 3632 20411 3634
rect 18646 3576 20350 3632
rect 20406 3576 20411 3632
rect 18646 3574 20411 3576
rect 0 3544 120 3574
rect 15101 3571 15167 3574
rect 20345 3571 20411 3574
rect 20486 3498 20546 3710
rect 22645 3707 22711 3710
rect 26969 3634 27035 3637
rect 2730 3438 20546 3498
rect 20670 3632 27035 3634
rect 20670 3576 26974 3632
rect 27030 3576 27035 3632
rect 20670 3574 27035 3576
rect 0 3362 120 3392
rect 2730 3362 2790 3438
rect 0 3302 2790 3362
rect 16205 3362 16271 3365
rect 20670 3362 20730 3574
rect 26969 3571 27035 3574
rect 38377 3634 38443 3637
rect 39808 3634 39928 3664
rect 38377 3632 39928 3634
rect 38377 3576 38382 3632
rect 38438 3576 39928 3632
rect 38377 3574 39928 3576
rect 38377 3571 38443 3574
rect 39808 3544 39928 3574
rect 22093 3498 22159 3501
rect 33777 3498 33843 3501
rect 22093 3496 33843 3498
rect 22093 3440 22098 3496
rect 22154 3440 33782 3496
rect 33838 3440 33843 3496
rect 22093 3438 33843 3440
rect 22093 3435 22159 3438
rect 33777 3435 33843 3438
rect 16205 3360 20730 3362
rect 16205 3304 16210 3360
rect 16266 3304 20730 3360
rect 16205 3302 20730 3304
rect 38009 3362 38075 3365
rect 39808 3362 39928 3392
rect 38009 3360 39928 3362
rect 38009 3304 38014 3360
rect 38070 3304 39928 3360
rect 38009 3302 39928 3304
rect 0 3272 120 3302
rect 16205 3299 16271 3302
rect 38009 3299 38075 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 39808 3272 39928 3302
rect 33006 3231 33322 3232
rect 0 3090 120 3120
rect 20897 3090 20963 3093
rect 0 3088 20963 3090
rect 0 3032 20902 3088
rect 20958 3032 20963 3088
rect 0 3030 20963 3032
rect 0 3000 120 3030
rect 20897 3027 20963 3030
rect 38377 3090 38443 3093
rect 39808 3090 39928 3120
rect 38377 3088 39928 3090
rect 38377 3032 38382 3088
rect 38438 3032 39928 3088
rect 38377 3030 39928 3032
rect 38377 3027 38443 3030
rect 39808 3000 39928 3030
rect 21541 2954 21607 2957
rect 1718 2952 21607 2954
rect 1718 2896 21546 2952
rect 21602 2896 21607 2952
rect 1718 2894 21607 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 21541 2891 21607 2894
rect 0 2758 1778 2818
rect 39113 2818 39179 2821
rect 39808 2818 39928 2848
rect 39113 2816 39928 2818
rect 39113 2760 39118 2816
rect 39174 2760 39928 2816
rect 39113 2758 39928 2760
rect 0 2728 120 2758
rect 39113 2755 39179 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 39808 2728 39928 2758
rect 37946 2687 38262 2688
rect 0 2546 120 2576
rect 22185 2546 22251 2549
rect 0 2544 22251 2546
rect 0 2488 22190 2544
rect 22246 2488 22251 2544
rect 0 2486 22251 2488
rect 0 2456 120 2486
rect 22185 2483 22251 2486
rect 38377 2546 38443 2549
rect 39808 2546 39928 2576
rect 38377 2544 39928 2546
rect 38377 2488 38382 2544
rect 38438 2488 39928 2544
rect 38377 2486 39928 2488
rect 38377 2483 38443 2486
rect 39808 2456 39928 2486
rect 9489 2410 9555 2413
rect 2822 2408 9555 2410
rect 2822 2352 9494 2408
rect 9550 2352 9555 2408
rect 2822 2350 9555 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 9489 2347 9555 2350
rect 10685 2410 10751 2413
rect 25221 2410 25287 2413
rect 10685 2408 25287 2410
rect 10685 2352 10690 2408
rect 10746 2352 25226 2408
rect 25282 2352 25287 2408
rect 10685 2350 25287 2352
rect 10685 2347 10751 2350
rect 25221 2347 25287 2350
rect 0 2214 2882 2274
rect 38009 2274 38075 2277
rect 39808 2274 39928 2304
rect 38009 2272 39928 2274
rect 38009 2216 38014 2272
rect 38070 2216 39928 2272
rect 38009 2214 39928 2216
rect 0 2184 120 2214
rect 38009 2211 38075 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 39808 2184 39928 2214
rect 33006 2143 33322 2144
rect 0 2002 120 2032
rect 18689 2002 18755 2005
rect 0 2000 18755 2002
rect 0 1944 18694 2000
rect 18750 1944 18755 2000
rect 0 1942 18755 1944
rect 0 1912 120 1942
rect 18689 1939 18755 1942
rect 36629 2002 36695 2005
rect 39808 2002 39928 2032
rect 36629 2000 39928 2002
rect 36629 1944 36634 2000
rect 36690 1944 39928 2000
rect 36629 1942 39928 1944
rect 36629 1939 36695 1942
rect 39808 1912 39928 1942
rect 12525 1866 12591 1869
rect 26509 1866 26575 1869
rect 12525 1864 26575 1866
rect 12525 1808 12530 1864
rect 12586 1808 26514 1864
rect 26570 1808 26575 1864
rect 12525 1806 26575 1808
rect 12525 1803 12591 1806
rect 26509 1803 26575 1806
rect 0 1730 120 1760
rect 9581 1730 9647 1733
rect 0 1728 9647 1730
rect 0 1672 9586 1728
rect 9642 1672 9647 1728
rect 0 1670 9647 1672
rect 0 1640 120 1670
rect 9581 1667 9647 1670
rect 37825 1730 37891 1733
rect 39808 1730 39928 1760
rect 37825 1728 39928 1730
rect 37825 1672 37830 1728
rect 37886 1672 39928 1728
rect 37825 1670 39928 1672
rect 37825 1667 37891 1670
rect 39808 1640 39928 1670
rect 0 1458 120 1488
rect 8569 1458 8635 1461
rect 0 1456 8635 1458
rect 0 1400 8574 1456
rect 8630 1400 8635 1456
rect 0 1398 8635 1400
rect 0 1368 120 1398
rect 8569 1395 8635 1398
rect 36997 1458 37063 1461
rect 39808 1458 39928 1488
rect 36997 1456 39928 1458
rect 36997 1400 37002 1456
rect 37058 1400 39928 1456
rect 36997 1398 39928 1400
rect 36997 1395 37063 1398
rect 39808 1368 39928 1398
rect 0 1186 120 1216
rect 7833 1186 7899 1189
rect 0 1184 7899 1186
rect 0 1128 7838 1184
rect 7894 1128 7899 1184
rect 0 1126 7899 1128
rect 0 1096 120 1126
rect 7833 1123 7899 1126
rect 37641 1186 37707 1189
rect 39808 1186 39928 1216
rect 37641 1184 39928 1186
rect 37641 1128 37646 1184
rect 37702 1128 39928 1184
rect 37641 1126 39928 1128
rect 37641 1123 37707 1126
rect 39808 1096 39928 1126
<< via3 >>
rect 19380 9964 19444 10028
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 19380 8196 19444 8260
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
<< metal4 >>
rect 1944 8192 2264 11152
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11152
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11152
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11152
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11152
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11152
rect 19379 10028 19445 10029
rect 19379 9964 19380 10028
rect 19444 9964 19445 10028
rect 19379 9963 19445 9964
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 19382 8261 19442 9963
rect 19379 8260 19445 8261
rect 19379 8196 19380 8260
rect 19444 8196 19445 8260
rect 19379 8195 19445 8196
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11152
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11152
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11152
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11152
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11152
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11152
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11152
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
use sky130_fd_sc_hd__buf_1  _000_
timestamp -3599
transform 1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 17572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform 1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 18676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _004_
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _005_
timestamp -3599
transform 1 0 22356 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 21252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _009_
timestamp -3599
transform 1 0 17020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 22080 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 19688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _014_
timestamp -3599
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _015_
timestamp -3599
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _018_
timestamp -3599
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _021_
timestamp -3599
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 22908 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _023_
timestamp -3599
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 22356 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _025_
timestamp -3599
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _026_
timestamp -3599
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _029_
timestamp -3599
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_
timestamp -3599
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _032_
timestamp -3599
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _033_
timestamp -3599
transform 1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _034_
timestamp -3599
transform 1 0 20424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _035_
timestamp -3599
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp -3599
transform -1 0 25668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp -3599
transform -1 0 26956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp -3599
transform -1 0 27508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _039_
timestamp -3599
transform 1 0 26956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _040_
timestamp -3599
transform 1 0 26128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp -3599
transform -1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp -3599
transform -1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform -1 0 28428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp -3599
transform -1 0 28520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform -1 0 29532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform -1 0 31464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform -1 0 33396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform -1 0 34960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform -1 0 36156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 37444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 37168 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp -3599
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp -3599
transform 1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp -3599
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp -3599
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp -3599
transform 1 0 10212 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp -3599
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp -3599
transform 1 0 8096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp -3599
transform 1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp -3599
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp -3599
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp -3599
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp -3599
transform 1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp -3599
transform 1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp -3599
transform 1 0 10212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp -3599
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp -3599
transform 1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp -3599
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp -3599
transform 1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp -3599
transform 1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp -3599
transform -1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp -3599
transform 1 0 16744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp -3599
transform 1 0 17020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp -3599
transform 1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform 1 0 15364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp -3599
transform 1 0 14904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform 1 0 14168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp -3599
transform 1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp -3599
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp -3599
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp -3599
transform 1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp -3599
transform 1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp -3599
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform 1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform 1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp -3599
transform 1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _088_
timestamp -3599
transform -1 0 24472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _089_
timestamp -3599
transform -1 0 25668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _090_
timestamp -3599
transform -1 0 26220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _091_
timestamp -3599
transform -1 0 25944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _092_
timestamp -3599
transform -1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _093_
timestamp -3599
transform -1 0 27416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _094_
timestamp -3599
transform -1 0 28152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _095_
timestamp -3599
transform -1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp -3599
transform -1 0 30084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp -3599
transform -1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _098_
timestamp -3599
transform -1 0 29808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _099_
timestamp -3599
transform -1 0 29532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _100_
timestamp -3599
transform -1 0 29072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _101_
timestamp -3599
transform -1 0 28428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp -3599
transform -1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp -3599
transform 1 0 26220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 21712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 21344 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform 1 0 19504 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 17940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 19504 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform 1 0 18676 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 21160 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform 1 0 20148 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform 1 0 22724 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 20608 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 22632 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 21712 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform 1 0 18216 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 23368 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform -1 0 19136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform 1 0 22172 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform 1 0 21068 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform -1 0 23092 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 26680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform -1 0 10212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 13064 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform -1 0 22080 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform 1 0 22172 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6
timestamp -3599
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp -3599
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12
timestamp -3599
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18
timestamp -3599
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21
timestamp -3599
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp -3599
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35
timestamp -3599
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp -3599
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp -3599
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47
timestamp -3599
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50
timestamp -3599
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60
timestamp -3599
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp -3599
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp -3599
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp -3599
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78
timestamp -3599
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_88
timestamp -3599
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91
timestamp -3599
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp -3599
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp -3599
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100
timestamp -3599
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103
timestamp -3599
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106
timestamp -3599
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_116
timestamp -3599
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp -3599
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_122
timestamp -3599
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp -3599
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_128
timestamp -3599
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_131
timestamp -3599
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_134
timestamp -3599
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_144
timestamp -3599
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_147
timestamp -3599
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_150
timestamp -3599
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_153
timestamp -3599
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp -3599
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_159
timestamp -3599
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_162
timestamp -3599
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_172
timestamp -3599
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_175
timestamp -3599
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_178
timestamp -3599
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp -3599
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_184
timestamp -3599
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp -3599
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_190
timestamp -3599
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_200
timestamp -3599
transform 1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_203
timestamp -3599
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_206
timestamp -3599
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_209
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_212
timestamp -3599
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_215
timestamp -3599
transform 1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp -3599
transform 1 0 21160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_228
timestamp -3599
transform 1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_231
timestamp -3599
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_234
timestamp -3599
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_237
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_240
timestamp -3599
transform 1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_243
timestamp -3599
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_246
timestamp -3599
transform 1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_256
timestamp -3599
transform 1 0 24656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_259
timestamp -3599
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_262
timestamp -3599
transform 1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_265
timestamp -3599
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_268
timestamp -3599
transform 1 0 25760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_271
timestamp -3599
transform 1 0 26036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_274
timestamp -3599
transform 1 0 26312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_281
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_284
timestamp -3599
transform 1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_287
timestamp -3599
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_290
timestamp -3599
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_293
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp -3599
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_299
timestamp -3599
transform 1 0 28612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_302
timestamp -3599
transform 1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_312
timestamp -3599
transform 1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_315
timestamp -3599
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_318
timestamp -3599
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_321
timestamp -3599
transform 1 0 30636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_324
timestamp -3599
transform 1 0 30912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_327
timestamp -3599
transform 1 0 31188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_330
timestamp -3599
transform 1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_337
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_340
timestamp -3599
transform 1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_343
timestamp -3599
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_346
timestamp -3599
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_349
timestamp -3599
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_352
timestamp -3599
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_355
timestamp -3599
transform 1 0 33764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_358
timestamp -3599
transform 1 0 34040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_365
timestamp -3599
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_368
timestamp -3599
transform 1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_371
timestamp -3599
transform 1 0 35236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_374
timestamp -3599
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp -3599
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_380
timestamp -3599
transform 1 0 36064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_383
timestamp -3599
transform 1 0 36340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6
timestamp -3599
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_9
timestamp -3599
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_12
timestamp -3599
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_15
timestamp -3599
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_18
timestamp -3599
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_21
timestamp -3599
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_24
timestamp -3599
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp -3599
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_30
timestamp -3599
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_33
timestamp -3599
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_36
timestamp -3599
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_39
timestamp -3599
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_42
timestamp -3599
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_45
timestamp -3599
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_48
timestamp -3599
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -3599
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_60
timestamp -3599
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_63
timestamp -3599
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_66
timestamp -3599
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp -3599
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_72
timestamp -3599
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_75
timestamp -3599
transform 1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp -3599
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp -3599
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_84
timestamp -3599
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_87
timestamp -3599
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_90
timestamp -3599
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_93
timestamp -3599
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_96
timestamp -3599
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_99
timestamp -3599
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp -3599
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_108
timestamp -3599
transform 1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_116
timestamp -3599
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp -3599
transform 1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_122
timestamp -3599
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp -3599
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_128
timestamp -3599
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_131
timestamp -3599
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_134
timestamp -3599
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_137
timestamp -3599
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_140
timestamp -3599
transform 1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp -3599
transform 1 0 14260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_146
timestamp -3599
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_149
timestamp -3599
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp -3599
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_155
timestamp -3599
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_158
timestamp -3599
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_164
timestamp -3599
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_172
timestamp -3599
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_175
timestamp -3599
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_178
timestamp -3599
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_181
timestamp -3599
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp -3599
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_187
timestamp -3599
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_190
timestamp -3599
transform 1 0 18584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_193
timestamp -3599
transform 1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_196
timestamp -3599
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_199
timestamp -3599
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_202
timestamp -3599
transform 1 0 19688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_205
timestamp -3599
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp -3599
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_211
timestamp -3599
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_214
timestamp -3599
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_217
timestamp -3599
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp -3599
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -3599
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_228
timestamp -3599
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_231
timestamp -3599
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_234
timestamp -3599
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_237
timestamp -3599
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_240
timestamp -3599
transform 1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_243
timestamp -3599
transform 1 0 23460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_246
timestamp -3599
transform 1 0 23736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_249
timestamp -3599
transform 1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_252
timestamp -3599
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_255
timestamp -3599
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_258
timestamp -3599
transform 1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_261
timestamp -3599
transform 1 0 25116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_264
timestamp -3599
transform 1 0 25392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_267
timestamp -3599
transform 1 0 25668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_270
timestamp -3599
transform 1 0 25944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_273
timestamp -3599
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_276
timestamp -3599
transform 1 0 26496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_284
timestamp -3599
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_287
timestamp -3599
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_290
timestamp -3599
transform 1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_293
timestamp -3599
transform 1 0 28060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_296
timestamp -3599
transform 1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_299
timestamp -3599
transform 1 0 28612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_302
timestamp -3599
transform 1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_305
timestamp -3599
transform 1 0 29164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_308
timestamp -3599
transform 1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_311
timestamp -3599
transform 1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_314
timestamp -3599
transform 1 0 29992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_317
timestamp -3599
transform 1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_320
timestamp -3599
transform 1 0 30544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_323
timestamp -3599
transform 1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_326
timestamp -3599
transform 1 0 31096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_329
timestamp -3599
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_332
timestamp -3599
transform 1 0 31648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_340
timestamp -3599
transform 1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_343
timestamp -3599
transform 1 0 32660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_346
timestamp -3599
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_349
timestamp -3599
transform 1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_352
timestamp -3599
transform 1 0 33488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_355
timestamp -3599
transform 1 0 33764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_358
timestamp -3599
transform 1 0 34040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_361
timestamp -3599
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_364
timestamp -3599
transform 1 0 34592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_367
timestamp -3599
transform 1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_370
timestamp -3599
transform 1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_373
timestamp -3599
transform 1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_376
timestamp -3599
transform 1 0 35696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_379
timestamp -3599
transform 1 0 35972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_382
timestamp -3599
transform 1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_385
timestamp -3599
transform 1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_388
timestamp -3599
transform 1 0 36800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp -3599
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_6
timestamp -3599
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_9
timestamp -3599
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_12
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_18
timestamp -3599
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_21
timestamp -3599
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_24
timestamp -3599
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp -3599
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_35
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_38
timestamp -3599
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp -3599
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_44
timestamp -3599
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_47
timestamp -3599
transform 1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp -3599
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp -3599
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp -3599
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_59
timestamp -3599
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_62
timestamp -3599
transform 1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_65
timestamp -3599
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp -3599
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_71
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_74
timestamp -3599
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_80
timestamp -3599
transform 1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_88
timestamp -3599
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_91
timestamp -3599
transform 1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_94
timestamp -3599
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp -3599
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_100
timestamp -3599
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_103
timestamp -3599
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_106
timestamp -3599
transform 1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp -3599
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_112
timestamp -3599
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_115
timestamp -3599
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_118
timestamp -3599
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_121
timestamp -3599
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_124
timestamp -3599
transform 1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_127
timestamp -3599
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_130
timestamp -3599
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_136
timestamp -3599
transform 1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_144
timestamp -3599
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_147
timestamp -3599
transform 1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp -3599
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_153
timestamp -3599
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_156
timestamp -3599
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_159
timestamp -3599
transform 1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_162
timestamp -3599
transform 1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_165
timestamp -3599
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_168
timestamp -3599
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_171
timestamp -3599
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_174
timestamp -3599
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_177
timestamp -3599
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_180
timestamp -3599
transform 1 0 17664 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_186
timestamp -3599
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_189
timestamp -3599
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_192
timestamp -3599
transform 1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -3599
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_200
timestamp -3599
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_203
timestamp -3599
transform 1 0 19780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_206
timestamp -3599
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp -3599
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_212
timestamp -3599
transform 1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_215
timestamp -3599
transform 1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_218
timestamp -3599
transform 1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_221
timestamp -3599
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_229
timestamp -3599
transform 1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_232
timestamp -3599
transform 1 0 22448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_235
timestamp -3599
transform 1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_238
timestamp -3599
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_241
timestamp -3599
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_244
timestamp -3599
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_247
timestamp -3599
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp -3599
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_256
timestamp -3599
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_259
timestamp -3599
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_267
timestamp -3599
transform 1 0 25668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_270
timestamp -3599
transform 1 0 25944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_275
timestamp -3599
transform 1 0 26404 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_287
timestamp -3599
transform 1 0 27508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_290
timestamp -3599
transform 1 0 27784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_293
timestamp -3599
transform 1 0 28060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_296
timestamp -3599
transform 1 0 28336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_299
timestamp -3599
transform 1 0 28612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_302
timestamp -3599
transform 1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp -3599
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_312
timestamp -3599
transform 1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_315
timestamp -3599
transform 1 0 30084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_318
timestamp -3599
transform 1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_321
timestamp -3599
transform 1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_324
timestamp -3599
transform 1 0 30912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_327
timestamp -3599
transform 1 0 31188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_330
timestamp -3599
transform 1 0 31464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_333
timestamp -3599
transform 1 0 31740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_336
timestamp -3599
transform 1 0 32016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_339
timestamp -3599
transform 1 0 32292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_342
timestamp -3599
transform 1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_345
timestamp -3599
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_348
timestamp -3599
transform 1 0 33120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_351
timestamp -3599
transform 1 0 33396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_354
timestamp -3599
transform 1 0 33672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_357
timestamp -3599
transform 1 0 33948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_360
timestamp -3599
transform 1 0 34224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp -3599
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_365
timestamp -3599
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_368
timestamp -3599
transform 1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_371
timestamp -3599
transform 1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_374
timestamp -3599
transform 1 0 35512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_377
timestamp -3599
transform 1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_380
timestamp -3599
transform 1 0 36064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_383
timestamp -3599
transform 1 0 36340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_386
timestamp -3599
transform 1 0 36616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_389
timestamp -3599
transform 1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_392
timestamp -3599
transform 1 0 37168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_395
timestamp -3599
transform 1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_398
timestamp -3599
transform 1 0 37720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_6
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_9
timestamp -3599
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_12
timestamp -3599
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_18
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_21
timestamp -3599
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_24
timestamp -3599
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp -3599
transform 1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_30
timestamp -3599
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_33
timestamp -3599
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_36
timestamp -3599
transform 1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_39
timestamp -3599
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_42
timestamp -3599
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_45
timestamp -3599
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_48
timestamp -3599
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp -3599
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_60
timestamp -3599
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_63
timestamp -3599
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_66
timestamp -3599
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_69
timestamp -3599
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_72
timestamp -3599
transform 1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_75
timestamp -3599
transform 1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_78
timestamp -3599
transform 1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_81
timestamp -3599
transform 1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_84
timestamp -3599
transform 1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_87
timestamp -3599
transform 1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_90
timestamp -3599
transform 1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_93
timestamp -3599
transform 1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_96
timestamp -3599
transform 1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_99
timestamp -3599
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_102
timestamp -3599
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_108
timestamp -3599
transform 1 0 11040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_116
timestamp -3599
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp -3599
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_122
timestamp -3599
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_125
timestamp -3599
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_128
timestamp -3599
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_131
timestamp -3599
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_134
timestamp -3599
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_137
timestamp -3599
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_140
timestamp -3599
transform 1 0 13984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_143
timestamp -3599
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_146
timestamp -3599
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_149
timestamp -3599
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_152
timestamp -3599
transform 1 0 15088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_159
timestamp -3599
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_162
timestamp -3599
transform 1 0 16008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_172
timestamp -3599
transform 1 0 16928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_176
timestamp -3599
transform 1 0 17296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp -3599
transform 1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_196
timestamp -3599
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_202
timestamp -3599
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_205
timestamp -3599
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp -3599
transform 1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_213
timestamp -3599
transform 1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_216
timestamp -3599
transform 1 0 20976 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_228
timestamp -3599
transform 1 0 22080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_239
timestamp -3599
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_242
timestamp -3599
transform 1 0 23368 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_245
timestamp -3599
transform 1 0 23644 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_248
timestamp -3599
transform 1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_251
timestamp -3599
transform 1 0 24196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_254
timestamp -3599
transform 1 0 24472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_257
timestamp -3599
transform 1 0 24748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_260
timestamp -3599
transform 1 0 25024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp -3599
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_266
timestamp -3599
transform 1 0 25576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_269
timestamp -3599
transform 1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_272
timestamp -3599
transform 1 0 26128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_275
timestamp -3599
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp -3599
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_284
timestamp -3599
transform 1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_287
timestamp -3599
transform 1 0 27508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_290
timestamp -3599
transform 1 0 27784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_293
timestamp -3599
transform 1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_296
timestamp -3599
transform 1 0 28336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_299
timestamp -3599
transform 1 0 28612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_302
timestamp -3599
transform 1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_305
timestamp -3599
transform 1 0 29164 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_308
timestamp -3599
transform 1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_311
timestamp -3599
transform 1 0 29716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_314
timestamp -3599
transform 1 0 29992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_317
timestamp -3599
transform 1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_320
timestamp -3599
transform 1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_323
timestamp -3599
transform 1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_326
timestamp -3599
transform 1 0 31096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_329
timestamp -3599
transform 1 0 31372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_332
timestamp -3599
transform 1 0 31648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp -3599
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_340
timestamp -3599
transform 1 0 32384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_343
timestamp -3599
transform 1 0 32660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_346
timestamp -3599
transform 1 0 32936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_349
timestamp -3599
transform 1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_352
timestamp -3599
transform 1 0 33488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_355
timestamp -3599
transform 1 0 33764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_358
timestamp -3599
transform 1 0 34040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_361
timestamp -3599
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_364
timestamp -3599
transform 1 0 34592 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_367
timestamp -3599
transform 1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_370
timestamp -3599
transform 1 0 35144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_373
timestamp -3599
transform 1 0 35420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_376
timestamp -3599
transform 1 0 35696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_379
timestamp -3599
transform 1 0 35972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_382
timestamp -3599
transform 1 0 36248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_388
timestamp -3599
transform 1 0 36800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_393
timestamp -3599
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_396
timestamp -3599
transform 1 0 37536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_6
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp -3599
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_12
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_18
timestamp -3599
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_21
timestamp -3599
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_24
timestamp -3599
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp -3599
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_35
timestamp -3599
transform 1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp -3599
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_44
timestamp -3599
transform 1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_47
timestamp -3599
transform 1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_50
timestamp -3599
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp -3599
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_56
timestamp -3599
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_59
timestamp -3599
transform 1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_62
timestamp -3599
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp -3599
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_68
timestamp -3599
transform 1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_71
timestamp -3599
transform 1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_74
timestamp -3599
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_80
timestamp -3599
transform 1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_88
timestamp -3599
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_91
timestamp -3599
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_94
timestamp -3599
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_100
timestamp -3599
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_103
timestamp -3599
transform 1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_106
timestamp -3599
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp -3599
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_112
timestamp -3599
transform 1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_115
timestamp -3599
transform 1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_118
timestamp -3599
transform 1 0 11960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_121
timestamp -3599
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_124
timestamp -3599
transform 1 0 12512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_127
timestamp -3599
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_130
timestamp -3599
transform 1 0 13064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_133
timestamp -3599
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_136
timestamp -3599
transform 1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_144
timestamp -3599
transform 1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_147
timestamp -3599
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp -3599
transform 1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_153
timestamp -3599
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp -3599
transform 1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_159
timestamp -3599
transform 1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_162
timestamp -3599
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp -3599
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_168
timestamp -3599
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_171
timestamp -3599
transform 1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_174
timestamp -3599
transform 1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_177
timestamp -3599
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_180
timestamp -3599
transform 1 0 17664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_183
timestamp -3599
transform 1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_186
timestamp -3599
transform 1 0 18216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_189
timestamp -3599
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_192
timestamp -3599
transform 1 0 18768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_200
timestamp -3599
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_203
timestamp -3599
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_206
timestamp -3599
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp -3599
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_212
timestamp -3599
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_215
timestamp -3599
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_223
timestamp -3599
transform 1 0 21620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_231
timestamp -3599
transform 1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_234
timestamp -3599
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_237
timestamp -3599
transform 1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_240
timestamp -3599
transform 1 0 23184 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_243
timestamp -3599
transform 1 0 23460 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_246
timestamp -3599
transform 1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp -3599
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_256
timestamp -3599
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_259
timestamp -3599
transform 1 0 24932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_262
timestamp -3599
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_265
timestamp -3599
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_268
timestamp -3599
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_271
timestamp -3599
transform 1 0 26036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_274
timestamp -3599
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_277
timestamp -3599
transform 1 0 26588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_280
timestamp -3599
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_283
timestamp -3599
transform 1 0 27140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_286
timestamp -3599
transform 1 0 27416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_289
timestamp -3599
transform 1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_292
timestamp -3599
transform 1 0 27968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_295
timestamp -3599
transform 1 0 28244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_298
timestamp -3599
transform 1 0 28520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_301
timestamp -3599
transform 1 0 28796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_304
timestamp -3599
transform 1 0 29072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_312
timestamp -3599
transform 1 0 29808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_315
timestamp -3599
transform 1 0 30084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_318
timestamp -3599
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_324
timestamp -3599
transform 1 0 30912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_327
timestamp -3599
transform 1 0 31188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_330
timestamp -3599
transform 1 0 31464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp -3599
transform 1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_336
timestamp -3599
transform 1 0 32016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_339
timestamp -3599
transform 1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_342
timestamp -3599
transform 1 0 32568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_345
timestamp -3599
transform 1 0 32844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_348
timestamp -3599
transform 1 0 33120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_351
timestamp -3599
transform 1 0 33396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_354
timestamp -3599
transform 1 0 33672 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_357
timestamp -3599
transform 1 0 33948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_360
timestamp -3599
transform 1 0 34224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp -3599
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_365
timestamp -3599
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_368
timestamp -3599
transform 1 0 34960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_371
timestamp -3599
transform 1 0 35236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_374
timestamp -3599
transform 1 0 35512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_377
timestamp -3599
transform 1 0 35788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_380
timestamp -3599
transform 1 0 36064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_383
timestamp -3599
transform 1 0 36340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_386
timestamp -3599
transform 1 0 36616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_389
timestamp -3599
transform 1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_392
timestamp -3599
transform 1 0 37168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_395
timestamp -3599
transform 1 0 37444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_398
timestamp -3599
transform 1 0 37720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_6
timestamp -3599
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_9
timestamp -3599
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp -3599
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_18
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_21
timestamp -3599
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp -3599
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_33
timestamp -3599
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_36
timestamp -3599
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_42
timestamp -3599
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_45
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_48
timestamp -3599
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_60
timestamp -3599
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_63
timestamp -3599
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_66
timestamp -3599
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_72
timestamp -3599
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp -3599
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_84
timestamp -3599
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_87
timestamp -3599
transform 1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_90
timestamp -3599
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp -3599
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_96
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_99
timestamp -3599
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_102
timestamp -3599
transform 1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_108
timestamp -3599
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_116
timestamp -3599
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp -3599
transform 1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_122
timestamp -3599
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp -3599
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_128
timestamp -3599
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_131
timestamp -3599
transform 1 0 13156 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_134
timestamp -3599
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_137
timestamp -3599
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_140
timestamp -3599
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp -3599
transform 1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_146
timestamp -3599
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp -3599
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_152
timestamp -3599
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_155
timestamp -3599
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_158
timestamp -3599
transform 1 0 15640 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_164
timestamp -3599
transform 1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_172
timestamp -3599
transform 1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_175
timestamp -3599
transform 1 0 17204 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_178
timestamp -3599
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_181
timestamp -3599
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp -3599
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_187
timestamp -3599
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_190
timestamp -3599
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_193
timestamp -3599
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_196
timestamp -3599
transform 1 0 19136 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp -3599
transform 1 0 19412 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_205
timestamp -3599
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_208
timestamp -3599
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_211
timestamp -3599
transform 1 0 20516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_214
timestamp -3599
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp -3599
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_228
timestamp -3599
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_231
timestamp -3599
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_234
timestamp -3599
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_237
timestamp -3599
transform 1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_240
timestamp -3599
transform 1 0 23184 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_243
timestamp -3599
transform 1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_246
timestamp -3599
transform 1 0 23736 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_249
timestamp -3599
transform 1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_252
timestamp -3599
transform 1 0 24288 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_255
timestamp -3599
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_258
timestamp -3599
transform 1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_261
timestamp -3599
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_264
timestamp -3599
transform 1 0 25392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_267
timestamp -3599
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_270
timestamp -3599
transform 1 0 25944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_276
timestamp -3599
transform 1 0 26496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_284
timestamp -3599
transform 1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_287
timestamp -3599
transform 1 0 27508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_290
timestamp -3599
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_296
timestamp -3599
transform 1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_299
timestamp -3599
transform 1 0 28612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_302
timestamp -3599
transform 1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_305
timestamp -3599
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_308
timestamp -3599
transform 1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_311
timestamp -3599
transform 1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_314
timestamp -3599
transform 1 0 29992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_317
timestamp -3599
transform 1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_320
timestamp -3599
transform 1 0 30544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_323
timestamp -3599
transform 1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_326
timestamp -3599
transform 1 0 31096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_329
timestamp -3599
transform 1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_332
timestamp -3599
transform 1 0 31648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp -3599
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_337
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_340
timestamp -3599
transform 1 0 32384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_343
timestamp -3599
transform 1 0 32660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_346
timestamp -3599
transform 1 0 32936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_349
timestamp -3599
transform 1 0 33212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_352
timestamp -3599
transform 1 0 33488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_355
timestamp -3599
transform 1 0 33764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_358
timestamp -3599
transform 1 0 34040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_361
timestamp -3599
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_364
timestamp -3599
transform 1 0 34592 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_367
timestamp -3599
transform 1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_370
timestamp -3599
transform 1 0 35144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_373
timestamp -3599
transform 1 0 35420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_376
timestamp -3599
transform 1 0 35696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_379
timestamp -3599
transform 1 0 35972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_382
timestamp -3599
transform 1 0 36248 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_388
timestamp -3599
transform 1 0 36800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_393
timestamp -3599
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_396
timestamp -3599
transform 1 0 37536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_6
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_9
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_12
timestamp -3599
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_15
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_18
timestamp -3599
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_21
timestamp -3599
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_24
timestamp -3599
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_38
timestamp -3599
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_44
timestamp -3599
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_47
timestamp -3599
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_50
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp -3599
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp -3599
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_59
timestamp -3599
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_62
timestamp -3599
transform 1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_65
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_68
timestamp -3599
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_71
timestamp -3599
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_74
timestamp -3599
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_77
timestamp -3599
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_80
timestamp -3599
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_88
timestamp -3599
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_91
timestamp -3599
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_94
timestamp -3599
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_97
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_100
timestamp -3599
transform 1 0 10304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_103
timestamp -3599
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_106
timestamp -3599
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_109
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_112
timestamp -3599
transform 1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_115
timestamp -3599
transform 1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_118
timestamp -3599
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp -3599
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_124
timestamp -3599
transform 1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_127
timestamp -3599
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_130
timestamp -3599
transform 1 0 13064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_136
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_144
timestamp -3599
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_147
timestamp -3599
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp -3599
transform 1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_153
timestamp -3599
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp -3599
transform 1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_159
timestamp -3599
transform 1 0 15732 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_162
timestamp -3599
transform 1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp -3599
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_168
timestamp -3599
transform 1 0 16560 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_171
timestamp -3599
transform 1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_174
timestamp -3599
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_177
timestamp -3599
transform 1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_180
timestamp -3599
transform 1 0 17664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_183
timestamp -3599
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_186
timestamp -3599
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_189
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_192
timestamp -3599
transform 1 0 18768 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_200
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_203
timestamp -3599
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_206
timestamp -3599
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_212
timestamp -3599
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp -3599
transform 1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_218
timestamp -3599
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_221
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_224
timestamp -3599
transform 1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_227
timestamp -3599
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_230
timestamp -3599
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_233
timestamp -3599
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_236
timestamp -3599
transform 1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_239
timestamp -3599
transform 1 0 23092 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_242
timestamp -3599
transform 1 0 23368 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_245
timestamp -3599
transform 1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_248
timestamp -3599
transform 1 0 23920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -3599
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_256
timestamp -3599
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_259
timestamp -3599
transform 1 0 24932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_262
timestamp -3599
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_268
timestamp -3599
transform 1 0 25760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_271
timestamp -3599
transform 1 0 26036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_274
timestamp -3599
transform 1 0 26312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_277
timestamp -3599
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_280
timestamp -3599
transform 1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_283
timestamp -3599
transform 1 0 27140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_286
timestamp -3599
transform 1 0 27416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_289
timestamp -3599
transform 1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_292
timestamp -3599
transform 1 0 27968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_297
timestamp -3599
transform 1 0 28428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_300
timestamp -3599
transform 1 0 28704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_303
timestamp -3599
transform 1 0 28980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp -3599
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_312
timestamp -3599
transform 1 0 29808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_315
timestamp -3599
transform 1 0 30084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_318
timestamp -3599
transform 1 0 30360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_321
timestamp -3599
transform 1 0 30636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_324
timestamp -3599
transform 1 0 30912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_330
timestamp -3599
transform 1 0 31464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_333
timestamp -3599
transform 1 0 31740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_336
timestamp -3599
transform 1 0 32016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_339
timestamp -3599
transform 1 0 32292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_342
timestamp -3599
transform 1 0 32568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_345
timestamp -3599
transform 1 0 32844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_351
timestamp -3599
transform 1 0 33396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_354
timestamp -3599
transform 1 0 33672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_357
timestamp -3599
transform 1 0 33948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_360
timestamp -3599
transform 1 0 34224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_368
timestamp -3599
transform 1 0 34960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_371
timestamp -3599
transform 1 0 35236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_374
timestamp -3599
transform 1 0 35512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_377
timestamp -3599
transform 1 0 35788 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_381
timestamp -3599
transform 1 0 36156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_384
timestamp -3599
transform 1 0 36432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_387
timestamp -3599
transform 1 0 36708 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_395
timestamp -3599
transform 1 0 37444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_398
timestamp -3599
transform 1 0 37720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_6
timestamp -3599
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_9
timestamp -3599
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_12
timestamp -3599
transform 1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_18
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_21
timestamp -3599
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_30
timestamp -3599
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_33
timestamp -3599
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_36
timestamp -3599
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_39
timestamp -3599
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_42
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_45
timestamp -3599
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_48
timestamp -3599
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp -3599
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_60
timestamp -3599
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_63
timestamp -3599
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_66
timestamp -3599
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp -3599
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp -3599
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_79
timestamp -3599
transform 1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_82
timestamp -3599
transform 1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_85
timestamp -3599
transform 1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_88
timestamp -3599
transform 1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_91
timestamp -3599
transform 1 0 9476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_94
timestamp -3599
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp -3599
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_106
timestamp -3599
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp -3599
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_116
timestamp -3599
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp -3599
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp -3599
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_125
timestamp -3599
transform 1 0 12604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_128
timestamp -3599
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_134
timestamp -3599
transform 1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_137
timestamp -3599
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_140
timestamp -3599
transform 1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_143
timestamp -3599
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_146
timestamp -3599
transform 1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_149
timestamp -3599
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_152
timestamp -3599
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_155
timestamp -3599
transform 1 0 15364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_158
timestamp -3599
transform 1 0 15640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_164
timestamp -3599
transform 1 0 16192 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_174
timestamp -3599
transform 1 0 17112 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_177
timestamp -3599
transform 1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_180
timestamp -3599
transform 1 0 17664 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_183
timestamp -3599
transform 1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_186
timestamp -3599
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_189
timestamp -3599
transform 1 0 18492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_192
timestamp -3599
transform 1 0 18768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_195
timestamp -3599
transform 1 0 19044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_198
timestamp -3599
transform 1 0 19320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_201
timestamp -3599
transform 1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_204
timestamp -3599
transform 1 0 19872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_207
timestamp -3599
transform 1 0 20148 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_210
timestamp -3599
transform 1 0 20424 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_213
timestamp -3599
transform 1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_216
timestamp -3599
transform 1 0 20976 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_219
timestamp -3599
transform 1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp -3599
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_228
timestamp -3599
transform 1 0 22080 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_233
timestamp -3599
transform 1 0 22540 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_236
timestamp -3599
transform 1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_239
timestamp -3599
transform 1 0 23092 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_242
timestamp -3599
transform 1 0 23368 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_245
timestamp -3599
transform 1 0 23644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_248
timestamp -3599
transform 1 0 23920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_251
timestamp -3599
transform 1 0 24196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_254
timestamp -3599
transform 1 0 24472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_257
timestamp -3599
transform 1 0 24748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_260
timestamp -3599
transform 1 0 25024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_263
timestamp -3599
transform 1 0 25300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_266
timestamp -3599
transform 1 0 25576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_269
timestamp -3599
transform 1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_272
timestamp -3599
transform 1 0 26128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_275
timestamp -3599
transform 1 0 26404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp -3599
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_284
timestamp -3599
transform 1 0 27232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_287
timestamp -3599
transform 1 0 27508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_290
timestamp -3599
transform 1 0 27784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_298
timestamp -3599
transform 1 0 28520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_301
timestamp -3599
transform 1 0 28796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_304
timestamp -3599
transform 1 0 29072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_309
timestamp -3599
transform 1 0 29532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_312
timestamp -3599
transform 1 0 29808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_315
timestamp -3599
transform 1 0 30084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_318
timestamp -3599
transform 1 0 30360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_321
timestamp -3599
transform 1 0 30636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_324
timestamp -3599
transform 1 0 30912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_327
timestamp -3599
transform 1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_330
timestamp -3599
transform 1 0 31464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp -3599
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_340
timestamp -3599
transform 1 0 32384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_343
timestamp -3599
transform 1 0 32660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_346
timestamp -3599
transform 1 0 32936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_349
timestamp -3599
transform 1 0 33212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_352
timestamp -3599
transform 1 0 33488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_355
timestamp -3599
transform 1 0 33764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_358
timestamp -3599
transform 1 0 34040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_361
timestamp -3599
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_364
timestamp -3599
transform 1 0 34592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_367
timestamp -3599
transform 1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_370
timestamp -3599
transform 1 0 35144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_373
timestamp -3599
transform 1 0 35420 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_376
timestamp -3599
transform 1 0 35696 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_379
timestamp -3599
transform 1 0 35972 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_382
timestamp -3599
transform 1 0 36248 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_385
timestamp -3599
transform 1 0 36524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_388
timestamp -3599
transform 1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_393
timestamp -3599
transform 1 0 37260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_396
timestamp -3599
transform 1 0 37536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_6
timestamp -3599
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_9
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_12
timestamp -3599
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp -3599
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_18
timestamp -3599
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_21
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp -3599
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_35
timestamp -3599
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp -3599
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp -3599
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_47
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_50
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp -3599
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_59
timestamp -3599
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_76
timestamp -3599
transform 1 0 8096 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_95
timestamp -3599
transform 1 0 9844 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_102
timestamp -3599
transform 1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_105
timestamp -3599
transform 1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_108
timestamp -3599
transform 1 0 11040 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_111
timestamp -3599
transform 1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_114
timestamp -3599
transform 1 0 11592 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_117
timestamp -3599
transform 1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_120
timestamp -3599
transform 1 0 12144 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_123
timestamp -3599
transform 1 0 12420 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_126
timestamp -3599
transform 1 0 12696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_147
timestamp -3599
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp -3599
transform 1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp -3599
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_159
timestamp -3599
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_162
timestamp -3599
transform 1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp -3599
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp -3599
transform 1 0 16560 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_171
timestamp -3599
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_174
timestamp -3599
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_180
timestamp -3599
transform 1 0 17664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_186
timestamp -3599
transform 1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_192
timestamp -3599
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_203
timestamp -3599
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_206
timestamp -3599
transform 1 0 20056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_212
timestamp -3599
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_215
timestamp -3599
transform 1 0 20884 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_221
timestamp -3599
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_224
timestamp -3599
transform 1 0 21712 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_227
timestamp -3599
transform 1 0 21988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_234
timestamp -3599
transform 1 0 22632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_240
timestamp -3599
transform 1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_243
timestamp -3599
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_246
timestamp -3599
transform 1 0 23736 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp -3599
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_256
timestamp -3599
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_259
timestamp -3599
transform 1 0 24932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_262
timestamp -3599
transform 1 0 25208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_276
timestamp -3599
transform 1 0 26496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_279
timestamp -3599
transform 1 0 26772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_289
timestamp -3599
transform 1 0 27692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_297
timestamp -3599
transform 1 0 28428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_301
timestamp -3599
transform 1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_304
timestamp -3599
transform 1 0 29072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_312
timestamp -3599
transform 1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_315
timestamp -3599
transform 1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_318
timestamp -3599
transform 1 0 30360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_321
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_324
timestamp -3599
transform 1 0 30912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_327
timestamp -3599
transform 1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_330
timestamp -3599
transform 1 0 31464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_333
timestamp -3599
transform 1 0 31740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_336
timestamp -3599
transform 1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_339
timestamp -3599
transform 1 0 32292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_342
timestamp -3599
transform 1 0 32568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_345
timestamp -3599
transform 1 0 32844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_348
timestamp -3599
transform 1 0 33120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_351
timestamp -3599
transform 1 0 33396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_354
timestamp -3599
transform 1 0 33672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_357
timestamp -3599
transform 1 0 33948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_360
timestamp -3599
transform 1 0 34224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp -3599
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_365
timestamp -3599
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_368
timestamp -3599
transform 1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_371
timestamp -3599
transform 1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_374
timestamp -3599
transform 1 0 35512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_377
timestamp -3599
transform 1 0 35788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_380
timestamp -3599
transform 1 0 36064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_383
timestamp -3599
transform 1 0 36340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_386
timestamp -3599
transform 1 0 36616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_389
timestamp -3599
transform 1 0 36892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_392
timestamp -3599
transform 1 0 37168 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6
timestamp -3599
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_9
timestamp -3599
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_12
timestamp -3599
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp -3599
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_18
timestamp -3599
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_21
timestamp -3599
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_24
timestamp -3599
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp -3599
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_30
timestamp -3599
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_33
timestamp -3599
transform 1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_36
timestamp -3599
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_39
timestamp -3599
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_42
timestamp -3599
transform 1 0 4968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_68
timestamp -3599
transform 1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_74
timestamp -3599
transform 1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_77
timestamp -3599
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_80
timestamp -3599
transform 1 0 8464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_83
timestamp -3599
transform 1 0 8740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_86
timestamp -3599
transform 1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_89
timestamp -3599
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_92
timestamp -3599
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_95
timestamp -3599
transform 1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_98
timestamp -3599
transform 1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_101
timestamp -3599
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_104
timestamp -3599
transform 1 0 10672 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_107
timestamp -3599
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp -3599
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_116
timestamp -3599
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp -3599
transform 1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_122
timestamp -3599
transform 1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_125
timestamp -3599
transform 1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_133
timestamp -3599
transform 1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_136
timestamp -3599
transform 1 0 13616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_148
timestamp -3599
transform 1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_153
timestamp -3599
transform 1 0 15180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_158
timestamp -3599
transform 1 0 15640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_162
timestamp -3599
transform 1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp -3599
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_176
timestamp -3599
transform 1 0 17296 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_179
timestamp -3599
transform 1 0 17572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_182
timestamp -3599
transform 1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_185
timestamp -3599
transform 1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_188
timestamp -3599
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_196
timestamp -3599
transform 1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_199
timestamp -3599
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_218
timestamp -3599
transform 1 0 21160 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_231
timestamp -3599
transform 1 0 22356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_242
timestamp -3599
transform 1 0 23368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_245
timestamp -3599
transform 1 0 23644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_248
timestamp -3599
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_254
timestamp -3599
transform 1 0 24472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_257
timestamp -3599
transform 1 0 24748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_260
timestamp -3599
transform 1 0 25024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_263
timestamp -3599
transform 1 0 25300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_266
timestamp -3599
transform 1 0 25576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_269
timestamp -3599
transform 1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_272
timestamp -3599
transform 1 0 26128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_275
timestamp -3599
transform 1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp -3599
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_284
timestamp -3599
transform 1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_287
timestamp -3599
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_290
timestamp -3599
transform 1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_293
timestamp -3599
transform 1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_296
timestamp -3599
transform 1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_299
timestamp -3599
transform 1 0 28612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_304
timestamp -3599
transform 1 0 29072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_318
timestamp -3599
transform 1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_321
timestamp -3599
transform 1 0 30636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_324
timestamp -3599
transform 1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_327
timestamp -3599
transform 1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_330
timestamp -3599
transform 1 0 31464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp -3599
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_340
timestamp -3599
transform 1 0 32384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_343
timestamp -3599
transform 1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_346
timestamp -3599
transform 1 0 32936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_349
timestamp -3599
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_352
timestamp -3599
transform 1 0 33488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_355
timestamp -3599
transform 1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_358
timestamp -3599
transform 1 0 34040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp -3599
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_364
timestamp -3599
transform 1 0 34592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_367
timestamp -3599
transform 1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_370
timestamp -3599
transform 1 0 35144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_373
timestamp -3599
transform 1 0 35420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_376
timestamp -3599
transform 1 0 35696 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_379
timestamp -3599
transform 1 0 35972 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_382
timestamp -3599
transform 1 0 36248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_385
timestamp -3599
transform 1 0 36524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_6
timestamp -3599
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_9
timestamp -3599
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_12
timestamp -3599
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_18
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_21
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp -3599
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp -3599
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_38
timestamp -3599
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_44
timestamp -3599
transform 1 0 5152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_50
timestamp -3599
transform 1 0 5704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp -3599
transform 1 0 5980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp -3599
transform 1 0 6532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_65
timestamp -3599
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp -3599
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_74
timestamp -3599
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -3599
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_92
timestamp -3599
transform 1 0 9568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_98
timestamp -3599
transform 1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_101
timestamp -3599
transform 1 0 10396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp -3599
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_110
timestamp -3599
transform 1 0 11224 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_116
timestamp -3599
transform 1 0 11776 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_122
timestamp -3599
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_125
timestamp -3599
transform 1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp -3599
transform 1 0 12880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_134
timestamp -3599
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_144
timestamp -3599
transform 1 0 14352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_149
timestamp -3599
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp -3599
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_158
timestamp -3599
transform 1 0 15640 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_161
timestamp -3599
transform 1 0 15916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_164
timestamp -3599
transform 1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_167
timestamp -3599
transform 1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_170
timestamp -3599
transform 1 0 16744 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_173
timestamp -3599
transform 1 0 17020 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_176
timestamp -3599
transform 1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_179
timestamp -3599
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_182
timestamp -3599
transform 1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_185
timestamp -3599
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_188
timestamp -3599
transform 1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_191
timestamp -3599
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp -3599
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_200
timestamp -3599
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_203
timestamp -3599
transform 1 0 19780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_206
timestamp -3599
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp -3599
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_212
timestamp -3599
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp -3599
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_218
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_221
timestamp -3599
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_224
timestamp -3599
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_227
timestamp -3599
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp -3599
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_233
timestamp -3599
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_236
timestamp -3599
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_239
timestamp -3599
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_242
timestamp -3599
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_248
timestamp -3599
transform 1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_256
timestamp -3599
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_259
timestamp -3599
transform 1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_262
timestamp -3599
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_265
timestamp -3599
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_268
timestamp -3599
transform 1 0 25760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_271
timestamp -3599
transform 1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_274
timestamp -3599
transform 1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_277
timestamp -3599
transform 1 0 26588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_280
timestamp -3599
transform 1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_283
timestamp -3599
transform 1 0 27140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_286
timestamp -3599
transform 1 0 27416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_289
timestamp -3599
transform 1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_292
timestamp -3599
transform 1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_295
timestamp -3599
transform 1 0 28244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_298
timestamp -3599
transform 1 0 28520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_301
timestamp -3599
transform 1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_304
timestamp -3599
transform 1 0 29072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_312
timestamp -3599
transform 1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_315
timestamp -3599
transform 1 0 30084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_318
timestamp -3599
transform 1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_321
timestamp -3599
transform 1 0 30636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_324
timestamp -3599
transform 1 0 30912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_327
timestamp -3599
transform 1 0 31188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_330
timestamp -3599
transform 1 0 31464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_333
timestamp -3599
transform 1 0 31740 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_336
timestamp -3599
transform 1 0 32016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_339
timestamp -3599
transform 1 0 32292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_342
timestamp -3599
transform 1 0 32568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_345
timestamp -3599
transform 1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_348
timestamp -3599
transform 1 0 33120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_351
timestamp -3599
transform 1 0 33396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_360
timestamp -3599
transform 1 0 34224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp -3599
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp -3599
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_371
timestamp -3599
transform 1 0 35236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_374
timestamp -3599
transform 1 0 35512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_377
timestamp -3599
transform 1 0 35788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_6
timestamp -3599
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_9
timestamp -3599
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_12
timestamp -3599
transform 1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp -3599
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp -3599
transform 1 0 17664 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_183
timestamp -3599
transform 1 0 17940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_186
timestamp -3599
transform 1 0 18216 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_189
timestamp -3599
transform 1 0 18492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_192
timestamp -3599
transform 1 0 18768 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_195
timestamp -3599
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_200
timestamp -3599
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_203
timestamp -3599
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_206
timestamp -3599
transform 1 0 20056 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_209
timestamp -3599
transform 1 0 20332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_212
timestamp -3599
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_215
timestamp -3599
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_218
timestamp -3599
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp -3599
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_228
timestamp -3599
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_231
timestamp -3599
transform 1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_234
timestamp -3599
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_237
timestamp -3599
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_240
timestamp -3599
transform 1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_243
timestamp -3599
transform 1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_246
timestamp -3599
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_249
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_253
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_256
timestamp -3599
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_259
timestamp -3599
transform 1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_262
timestamp -3599
transform 1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_265
timestamp -3599
transform 1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_268
timestamp -3599
transform 1 0 25760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_271
timestamp -3599
transform 1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_274
timestamp -3599
transform 1 0 26312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp -3599
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_284
timestamp -3599
transform 1 0 27232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_287
timestamp -3599
transform 1 0 27508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_290
timestamp -3599
transform 1 0 27784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_293
timestamp -3599
transform 1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_296
timestamp -3599
transform 1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_299
timestamp -3599
transform 1 0 28612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_302
timestamp -3599
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp -3599
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_309
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_312
timestamp -3599
transform 1 0 29808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_315
timestamp -3599
transform 1 0 30084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_318
timestamp -3599
transform 1 0 30360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_321
timestamp -3599
transform 1 0 30636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_324
timestamp -3599
transform 1 0 30912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_327
timestamp -3599
transform 1 0 31188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_330
timestamp -3599
transform 1 0 31464 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp -3599
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_361
timestamp -3599
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_401
timestamp -3599
transform 1 0 37996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 37812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 37444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 37812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 37444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 37444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 36432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 37812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 37812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform 1 0 35420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform 1 0 34868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform 1 0 36156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 35972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 36340 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform 1 0 32476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 32844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 33580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 33948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform 1 0 33488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform 1 0 33856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform 1 0 34684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform -1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform -1 0 3496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform -1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform -1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform -1 0 4600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform -1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform -1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform -1 0 6532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform -1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform -1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform -1 0 7912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform -1 0 8740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform -1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform -1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform -1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform -1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform -1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform -1 0 10120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform -1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 16560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform -1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform -1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 13432 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 13984 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 14812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform -1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 31832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1096 120 1216 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 39808 1096 39928 1216 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 39808 3816 39928 3936 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 39808 4088 39928 4208 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 39808 4360 39928 4480 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 39808 4632 39928 4752 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 39808 4904 39928 5024 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 39808 5176 39928 5296 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 39808 5448 39928 5568 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 39808 5720 39928 5840 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 39808 5992 39928 6112 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 39808 6264 39928 6384 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 39808 1368 39928 1488 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 39808 6536 39928 6656 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 39808 6808 39928 6928 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 39808 7080 39928 7200 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 39808 7352 39928 7472 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 39808 7624 39928 7744 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 39808 7896 39928 8016 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 39808 8168 39928 8288 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 39808 8440 39928 8560 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 39808 8712 39928 8832 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 39808 8984 39928 9104 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 39808 1640 39928 1760 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 39808 9256 39928 9376 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 39808 9528 39928 9648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 39808 1912 39928 2032 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 39808 2184 39928 2304 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 39808 2456 39928 2576 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 39808 2728 39928 2848 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 39808 3000 39928 3120 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 39808 3272 39928 3392 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 39808 3544 39928 3664 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 3330 0 3386 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 21730 0 21786 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 23570 0 23626 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 25410 0 25466 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 27250 0 27306 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 29090 0 29146 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 30930 0 30986 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 32770 0 32826 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 34610 0 34666 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 36450 0 36506 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 38290 0 38346 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 5170 0 5226 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 7010 0 7066 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 8850 0 8906 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 10690 0 10746 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 12530 0 12586 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 14370 0 14426 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 16210 0 16266 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 18050 0 18106 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 19890 0 19946 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 31758 11096 31814 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 34518 11096 34574 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 34794 11096 34850 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 35070 11096 35126 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 35346 11096 35402 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 35622 11096 35678 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 35898 11096 35954 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 36174 11096 36230 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 36450 11096 36506 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 36726 11096 36782 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 37002 11096 37058 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 32034 11096 32090 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 32310 11096 32366 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 32586 11096 32642 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 32862 11096 32918 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 33138 11096 33194 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 33414 11096 33470 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 33690 11096 33746 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 33966 11096 34022 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 34242 11096 34298 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 2778 11096 2834 11152 0 FreeSans 224 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 3054 11096 3110 11152 0 FreeSans 224 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 3330 11096 3386 11152 0 FreeSans 224 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 3606 11096 3662 11152 0 FreeSans 224 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 3882 11096 3938 11152 0 FreeSans 224 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 4158 11096 4214 11152 0 FreeSans 224 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 4434 11096 4490 11152 0 FreeSans 224 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 4710 11096 4766 11152 0 FreeSans 224 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 4986 11096 5042 11152 0 FreeSans 224 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 5262 11096 5318 11152 0 FreeSans 224 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 5538 11096 5594 11152 0 FreeSans 224 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 5814 11096 5870 11152 0 FreeSans 224 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 6090 11096 6146 11152 0 FreeSans 224 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 6366 11096 6422 11152 0 FreeSans 224 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 6642 11096 6698 11152 0 FreeSans 224 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 6918 11096 6974 11152 0 FreeSans 224 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 7194 11096 7250 11152 0 FreeSans 224 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 7470 11096 7526 11152 0 FreeSans 224 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 7746 11096 7802 11152 0 FreeSans 224 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 8022 11096 8078 11152 0 FreeSans 224 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 8298 11096 8354 11152 0 FreeSans 224 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 11058 11096 11114 11152 0 FreeSans 224 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 11334 11096 11390 11152 0 FreeSans 224 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 11610 11096 11666 11152 0 FreeSans 224 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 11886 11096 11942 11152 0 FreeSans 224 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 12162 11096 12218 11152 0 FreeSans 224 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 12438 11096 12494 11152 0 FreeSans 224 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 8574 11096 8630 11152 0 FreeSans 224 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 8850 11096 8906 11152 0 FreeSans 224 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 9126 11096 9182 11152 0 FreeSans 224 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 9402 11096 9458 11152 0 FreeSans 224 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 9678 11096 9734 11152 0 FreeSans 224 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 9954 11096 10010 11152 0 FreeSans 224 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 10230 11096 10286 11152 0 FreeSans 224 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 10506 11096 10562 11152 0 FreeSans 224 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 10782 11096 10838 11152 0 FreeSans 224 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 12714 11096 12770 11152 0 FreeSans 224 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal2 s 15474 11096 15530 11152 0 FreeSans 224 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal2 s 15750 11096 15806 11152 0 FreeSans 224 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal2 s 16026 11096 16082 11152 0 FreeSans 224 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal2 s 16302 11096 16358 11152 0 FreeSans 224 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal2 s 16578 11096 16634 11152 0 FreeSans 224 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal2 s 16854 11096 16910 11152 0 FreeSans 224 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal2 s 12990 11096 13046 11152 0 FreeSans 224 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal2 s 13266 11096 13322 11152 0 FreeSans 224 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal2 s 13542 11096 13598 11152 0 FreeSans 224 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal2 s 13818 11096 13874 11152 0 FreeSans 224 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal2 s 14094 11096 14150 11152 0 FreeSans 224 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal2 s 14370 11096 14426 11152 0 FreeSans 224 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal2 s 14646 11096 14702 11152 0 FreeSans 224 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal2 s 14922 11096 14978 11152 0 FreeSans 224 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal2 s 15198 11096 15254 11152 0 FreeSans 224 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal2 s 17130 11096 17186 11152 0 FreeSans 224 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal2 s 17406 11096 17462 11152 0 FreeSans 224 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal2 s 17682 11096 17738 11152 0 FreeSans 224 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal2 s 17958 11096 18014 11152 0 FreeSans 224 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal2 s 20442 11096 20498 11152 0 FreeSans 224 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal2 s 20718 11096 20774 11152 0 FreeSans 224 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal2 s 20994 11096 21050 11152 0 FreeSans 224 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal2 s 21270 11096 21326 11152 0 FreeSans 224 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal2 s 21546 11096 21602 11152 0 FreeSans 224 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal2 s 21822 11096 21878 11152 0 FreeSans 224 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal2 s 22098 11096 22154 11152 0 FreeSans 224 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal2 s 22374 11096 22430 11152 0 FreeSans 224 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal2 s 18234 11096 18290 11152 0 FreeSans 224 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal2 s 18510 11096 18566 11152 0 FreeSans 224 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal2 s 18786 11096 18842 11152 0 FreeSans 224 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal2 s 19062 11096 19118 11152 0 FreeSans 224 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal2 s 19338 11096 19394 11152 0 FreeSans 224 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal2 s 19614 11096 19670 11152 0 FreeSans 224 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal2 s 19890 11096 19946 11152 0 FreeSans 224 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal2 s 20166 11096 20222 11152 0 FreeSans 224 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal2 s 22650 11096 22706 11152 0 FreeSans 224 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal2 s 25410 11096 25466 11152 0 FreeSans 224 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal2 s 25686 11096 25742 11152 0 FreeSans 224 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal2 s 25962 11096 26018 11152 0 FreeSans 224 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal2 s 26238 11096 26294 11152 0 FreeSans 224 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal2 s 26514 11096 26570 11152 0 FreeSans 224 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal2 s 26790 11096 26846 11152 0 FreeSans 224 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal2 s 22926 11096 22982 11152 0 FreeSans 224 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal2 s 23202 11096 23258 11152 0 FreeSans 224 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal2 s 23478 11096 23534 11152 0 FreeSans 224 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal2 s 23754 11096 23810 11152 0 FreeSans 224 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal2 s 24030 11096 24086 11152 0 FreeSans 224 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal2 s 24306 11096 24362 11152 0 FreeSans 224 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal2 s 24582 11096 24638 11152 0 FreeSans 224 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal2 s 24858 11096 24914 11152 0 FreeSans 224 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal2 s 25134 11096 25190 11152 0 FreeSans 224 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal2 s 27066 11096 27122 11152 0 FreeSans 224 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal2 s 29826 11096 29882 11152 0 FreeSans 224 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal2 s 30102 11096 30158 11152 0 FreeSans 224 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal2 s 30378 11096 30434 11152 0 FreeSans 224 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal2 s 30654 11096 30710 11152 0 FreeSans 224 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal2 s 30930 11096 30986 11152 0 FreeSans 224 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal2 s 31206 11096 31262 11152 0 FreeSans 224 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal2 s 27342 11096 27398 11152 0 FreeSans 224 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal2 s 27618 11096 27674 11152 0 FreeSans 224 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal2 s 27894 11096 27950 11152 0 FreeSans 224 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal2 s 28170 11096 28226 11152 0 FreeSans 224 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal2 s 28446 11096 28502 11152 0 FreeSans 224 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal2 s 28722 11096 28778 11152 0 FreeSans 224 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal2 s 28998 11096 29054 11152 0 FreeSans 224 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal2 s 29274 11096 29330 11152 0 FreeSans 224 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal2 s 29550 11096 29606 11152 0 FreeSans 224 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal2 s 1490 0 1546 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 31482 11096 31538 11152 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3004 0 3324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 11092 3324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 11092 9324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 11092 15324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 11092 21324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 11092 27324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 11092 33324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 11092 2264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 11092 8264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 11092 14264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 11092 20264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 11092 26264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 11092 32264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 11092 38264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 19964 8704 19964 8704 0 VGND
rlabel via1 19964 8160 19964 8160 0 VPWR
rlabel metal3 3978 1156 3978 1156 0 FrameData[0]
rlabel metal3 919 3876 919 3876 0 FrameData[10]
rlabel metal1 17848 4658 17848 4658 0 FrameData[11]
rlabel via2 21206 4539 21206 4539 0 FrameData[12]
rlabel metal2 19780 5202 19780 5202 0 FrameData[13]
rlabel metal3 919 4964 919 4964 0 FrameData[14]
rlabel metal2 17802 5933 17802 5933 0 FrameData[15]
rlabel metal3 620 5508 620 5508 0 FrameData[16]
rlabel metal2 7590 5423 7590 5423 0 FrameData[17]
rlabel metal3 942 6052 942 6052 0 FrameData[18]
rlabel metal3 1195 6324 1195 6324 0 FrameData[19]
rlabel metal3 4346 1428 4346 1428 0 FrameData[1]
rlabel metal2 16238 6800 16238 6800 0 FrameData[20]
rlabel metal1 19734 6698 19734 6698 0 FrameData[21]
rlabel metal3 666 7140 666 7140 0 FrameData[22]
rlabel metal1 19918 7242 19918 7242 0 FrameData[23]
rlabel metal3 712 7684 712 7684 0 FrameData[24]
rlabel metal3 620 7956 620 7956 0 FrameData[25]
rlabel metal3 942 8228 942 8228 0 FrameData[26]
rlabel metal3 712 8500 712 8500 0 FrameData[27]
rlabel metal3 528 8772 528 8772 0 FrameData[28]
rlabel metal3 344 9044 344 9044 0 FrameData[29]
rlabel metal3 4852 1700 4852 1700 0 FrameData[2]
rlabel metal2 20378 8347 20378 8347 0 FrameData[30]
rlabel metal3 735 9588 735 9588 0 FrameData[31]
rlabel metal3 9406 1972 9406 1972 0 FrameData[3]
rlabel metal3 1471 2244 1471 2244 0 FrameData[4]
rlabel metal3 11154 2516 11154 2516 0 FrameData[5]
rlabel metal3 919 2788 919 2788 0 FrameData[6]
rlabel metal1 21022 3910 21022 3910 0 FrameData[7]
rlabel metal3 20516 3604 20516 3604 0 FrameData[8]
rlabel metal1 17066 4046 17066 4046 0 FrameData[9]
rlabel metal3 38756 1156 38756 1156 0 FrameData_O[0]
rlabel metal3 39492 3876 39492 3876 0 FrameData_O[10]
rlabel metal3 39124 4148 39124 4148 0 FrameData_O[11]
rlabel metal3 38940 4420 38940 4420 0 FrameData_O[12]
rlabel metal3 39124 4692 39124 4692 0 FrameData_O[13]
rlabel metal3 39492 4964 39492 4964 0 FrameData_O[14]
rlabel metal3 39124 5236 39124 5236 0 FrameData_O[15]
rlabel metal3 38940 5508 38940 5508 0 FrameData_O[16]
rlabel metal3 39124 5780 39124 5780 0 FrameData_O[17]
rlabel metal3 39722 6052 39722 6052 0 FrameData_O[18]
rlabel metal3 38756 6324 38756 6324 0 FrameData_O[19]
rlabel metal3 38434 1428 38434 1428 0 FrameData_O[1]
rlabel metal2 38410 6511 38410 6511 0 FrameData_O[20]
rlabel metal3 38434 6868 38434 6868 0 FrameData_O[21]
rlabel metal3 39124 7140 39124 7140 0 FrameData_O[22]
rlabel metal3 38940 7412 38940 7412 0 FrameData_O[23]
rlabel metal3 39124 7684 39124 7684 0 FrameData_O[24]
rlabel metal3 39124 7956 39124 7956 0 FrameData_O[25]
rlabel metal1 38180 8058 38180 8058 0 FrameData_O[26]
rlabel metal1 38180 7514 38180 7514 0 FrameData_O[27]
rlabel metal2 36938 8415 36938 8415 0 FrameData_O[28]
rlabel metal1 38456 6630 38456 6630 0 FrameData_O[29]
rlabel metal3 38848 1700 38848 1700 0 FrameData_O[2]
rlabel metal2 37674 8415 37674 8415 0 FrameData_O[30]
rlabel metal1 38042 6664 38042 6664 0 FrameData_O[31]
rlabel metal3 38250 1972 38250 1972 0 FrameData_O[3]
rlabel metal3 38940 2244 38940 2244 0 FrameData_O[4]
rlabel metal3 39124 2516 39124 2516 0 FrameData_O[5]
rlabel metal3 39492 2788 39492 2788 0 FrameData_O[6]
rlabel metal3 39124 3060 39124 3060 0 FrameData_O[7]
rlabel metal3 38940 3332 38940 3332 0 FrameData_O[8]
rlabel metal3 39124 3604 39124 3604 0 FrameData_O[9]
rlabel metal2 3358 1007 3358 1007 0 FrameStrobe[0]
rlabel metal2 21758 55 21758 55 0 FrameStrobe[10]
rlabel metal1 25898 5678 25898 5678 0 FrameStrobe[11]
rlabel metal2 25438 1401 25438 1401 0 FrameStrobe[12]
rlabel metal2 27278 735 27278 735 0 FrameStrobe[13]
rlabel metal1 30176 5678 30176 5678 0 FrameStrobe[14]
rlabel metal1 32453 5678 32453 5678 0 FrameStrobe[15]
rlabel metal1 33028 5610 33028 5610 0 FrameStrobe[16]
rlabel metal1 35282 5610 35282 5610 0 FrameStrobe[17]
rlabel metal1 36754 5610 36754 5610 0 FrameStrobe[18]
rlabel metal1 37628 6086 37628 6086 0 FrameStrobe[19]
rlabel metal2 5198 2078 5198 2078 0 FrameStrobe[1]
rlabel metal2 20470 3604 20470 3604 0 FrameStrobe[2]
rlabel metal2 17158 3876 17158 3876 0 FrameStrobe[3]
rlabel metal2 10718 1211 10718 1211 0 FrameStrobe[4]
rlabel metal2 12558 939 12558 939 0 FrameStrobe[5]
rlabel metal2 14398 1058 14398 1058 0 FrameStrobe[6]
rlabel metal3 18469 3332 18469 3332 0 FrameStrobe[7]
rlabel metal2 18078 1806 18078 1806 0 FrameStrobe[8]
rlabel metal2 19918 786 19918 786 0 FrameStrobe[9]
rlabel metal1 32062 8602 32062 8602 0 FrameStrobe_O[0]
rlabel metal1 35650 8364 35650 8364 0 FrameStrobe_O[10]
rlabel metal1 34960 8058 34960 8058 0 FrameStrobe_O[11]
rlabel metal1 35558 8602 35558 8602 0 FrameStrobe_O[12]
rlabel metal1 36064 8330 36064 8330 0 FrameStrobe_O[13]
rlabel metal1 36754 8364 36754 8364 0 FrameStrobe_O[14]
rlabel metal1 36064 8058 36064 8058 0 FrameStrobe_O[15]
rlabel metal1 36432 8058 36432 8058 0 FrameStrobe_O[16]
rlabel metal1 36984 8602 36984 8602 0 FrameStrobe_O[17]
rlabel metal1 37858 8568 37858 8568 0 FrameStrobe_O[18]
rlabel metal1 37168 8058 37168 8058 0 FrameStrobe_O[19]
rlabel metal1 32384 8330 32384 8330 0 FrameStrobe_O[1]
rlabel metal1 32752 8602 32752 8602 0 FrameStrobe_O[2]
rlabel metal1 33442 8568 33442 8568 0 FrameStrobe_O[3]
rlabel metal1 33350 8330 33350 8330 0 FrameStrobe_O[4]
rlabel metal2 34178 8568 34178 8568 0 FrameStrobe_O[5]
rlabel metal1 33580 8058 33580 8058 0 FrameStrobe_O[6]
rlabel metal1 33948 8058 33948 8058 0 FrameStrobe_O[7]
rlabel metal1 34454 8602 34454 8602 0 FrameStrobe_O[8]
rlabel metal1 34776 8330 34776 8330 0 FrameStrobe_O[9]
rlabel metal2 2806 9856 2806 9856 0 N1BEG[0]
rlabel metal1 3082 8058 3082 8058 0 N1BEG[1]
rlabel metal1 3266 8602 3266 8602 0 N1BEG[2]
rlabel metal1 3772 8058 3772 8058 0 N1BEG[3]
rlabel metal1 3680 8330 3680 8330 0 N2BEG[0]
rlabel metal1 4278 8058 4278 8058 0 N2BEG[1]
rlabel metal1 4324 8602 4324 8602 0 N2BEG[2]
rlabel metal1 4646 8602 4646 8602 0 N2BEG[3]
rlabel metal1 4968 8602 4968 8602 0 N2BEG[4]
rlabel metal1 5382 8058 5382 8058 0 N2BEG[5]
rlabel metal1 5428 8602 5428 8602 0 N2BEG[6]
rlabel metal1 5796 8602 5796 8602 0 N2BEG[7]
rlabel metal1 6210 8058 6210 8058 0 N2BEGb[0]
rlabel metal1 6210 8602 6210 8602 0 N2BEGb[1]
rlabel metal1 6762 8058 6762 8058 0 N2BEGb[2]
rlabel metal1 6854 8602 6854 8602 0 N2BEGb[3]
rlabel metal1 7176 8602 7176 8602 0 N2BEGb[4]
rlabel metal1 7590 8058 7590 8058 0 N2BEGb[5]
rlabel metal1 7636 8602 7636 8602 0 N2BEGb[6]
rlabel metal1 8004 8602 8004 8602 0 N2BEGb[7]
rlabel metal1 8418 8058 8418 8058 0 N4BEG[0]
rlabel metal1 10948 8602 10948 8602 0 N4BEG[10]
rlabel metal1 11454 8058 11454 8058 0 N4BEG[11]
rlabel metal1 11408 8602 11408 8602 0 N4BEG[12]
rlabel metal1 12006 8058 12006 8058 0 N4BEG[13]
rlabel metal1 12052 8602 12052 8602 0 N4BEG[14]
rlabel metal2 12466 9856 12466 9856 0 N4BEG[15]
rlabel metal1 8372 8602 8372 8602 0 N4BEG[1]
rlabel metal1 8694 8602 8694 8602 0 N4BEG[2]
rlabel metal1 9108 8058 9108 8058 0 N4BEG[3]
rlabel metal1 9384 8602 9384 8602 0 N4BEG[4]
rlabel metal1 9798 8058 9798 8058 0 N4BEG[5]
rlabel metal1 9844 8602 9844 8602 0 N4BEG[6]
rlabel metal1 10166 8602 10166 8602 0 N4BEG[7]
rlabel metal1 10488 8602 10488 8602 0 N4BEG[8]
rlabel metal1 10902 8058 10902 8058 0 N4BEG[9]
rlabel metal1 12696 8602 12696 8602 0 NN4BEG[0]
rlabel metal1 15364 8602 15364 8602 0 NN4BEG[10]
rlabel metal1 15686 8602 15686 8602 0 NN4BEG[11]
rlabel metal1 16008 8602 16008 8602 0 NN4BEG[12]
rlabel metal2 16330 9856 16330 9856 0 NN4BEG[13]
rlabel metal1 17020 8330 17020 8330 0 NN4BEG[14]
rlabel metal1 16974 8602 16974 8602 0 NN4BEG[15]
rlabel metal1 13110 8058 13110 8058 0 NN4BEG[1]
rlabel metal1 13156 8602 13156 8602 0 NN4BEG[2]
rlabel metal1 13662 8058 13662 8058 0 NN4BEG[3]
rlabel metal1 13616 8330 13616 8330 0 NN4BEG[4]
rlabel metal1 13938 8602 13938 8602 0 NN4BEG[5]
rlabel metal1 14490 8058 14490 8058 0 NN4BEG[6]
rlabel metal1 14582 8602 14582 8602 0 NN4BEG[7]
rlabel metal1 14904 8602 14904 8602 0 NN4BEG[8]
rlabel metal2 15410 8755 15410 8755 0 NN4BEG[9]
rlabel metal2 17158 10621 17158 10621 0 S1END[0]
rlabel metal2 17434 10332 17434 10332 0 S1END[1]
rlabel metal2 17710 10502 17710 10502 0 S1END[2]
rlabel metal2 17986 11046 17986 11046 0 S1END[3]
rlabel metal2 20470 8598 20470 8598 0 S2END[0]
rlabel metal2 20746 10944 20746 10944 0 S2END[1]
rlabel metal2 21022 11097 21022 11097 0 S2END[2]
rlabel metal2 21298 11029 21298 11029 0 S2END[3]
rlabel metal2 21574 11012 21574 11012 0 S2END[4]
rlabel via2 21850 11097 21850 11097 0 S2END[5]
rlabel metal1 10442 11084 10442 11084 0 S2END[6]
rlabel metal2 10994 8670 10994 8670 0 S2END[7]
rlabel metal2 18262 10026 18262 10026 0 S2MID[0]
rlabel metal2 18538 10536 18538 10536 0 S2MID[1]
rlabel metal2 18814 10434 18814 10434 0 S2MID[2]
rlabel metal2 19090 9584 19090 9584 0 S2MID[3]
rlabel metal2 19366 9533 19366 9533 0 S2MID[4]
rlabel metal2 19642 9958 19642 9958 0 S2MID[5]
rlabel metal2 19918 10060 19918 10060 0 S2MID[6]
rlabel metal2 20194 10009 20194 10009 0 S2MID[7]
rlabel metal2 14766 8211 14766 8211 0 S4END[0]
rlabel metal2 16422 8075 16422 8075 0 S4END[10]
rlabel metal2 16698 8636 16698 8636 0 S4END[11]
rlabel metal2 15594 7548 15594 7548 0 S4END[12]
rlabel metal2 16514 9095 16514 9095 0 S4END[13]
rlabel metal2 17250 7599 17250 7599 0 S4END[14]
rlabel via2 19550 7429 19550 7429 0 S4END[15]
rlabel metal2 14306 6154 14306 6154 0 S4END[1]
rlabel metal2 14490 9622 14490 9622 0 S4END[2]
rlabel metal2 13018 6256 13018 6256 0 S4END[3]
rlabel metal2 23782 8700 23782 8700 0 S4END[4]
rlabel metal1 13524 7378 13524 7378 0 S4END[5]
rlabel metal2 13294 6222 13294 6222 0 S4END[6]
rlabel metal2 21574 8194 21574 8194 0 S4END[7]
rlabel metal2 17894 6477 17894 6477 0 S4END[8]
rlabel metal2 20746 7769 20746 7769 0 S4END[9]
rlabel metal2 27094 11097 27094 11097 0 SS4END[0]
rlabel metal2 29854 8972 29854 8972 0 SS4END[10]
rlabel metal2 30130 8632 30130 8632 0 SS4END[11]
rlabel metal2 30406 10434 30406 10434 0 SS4END[12]
rlabel metal2 30682 10400 30682 10400 0 SS4END[13]
rlabel metal2 30958 10502 30958 10502 0 SS4END[14]
rlabel metal2 31234 10570 31234 10570 0 SS4END[15]
rlabel metal2 27370 9261 27370 9261 0 SS4END[1]
rlabel metal2 27646 11097 27646 11097 0 SS4END[2]
rlabel metal2 27922 9244 27922 9244 0 SS4END[3]
rlabel metal2 28198 10213 28198 10213 0 SS4END[4]
rlabel metal2 28474 10145 28474 10145 0 SS4END[5]
rlabel metal2 28750 10281 28750 10281 0 SS4END[6]
rlabel metal2 29026 9584 29026 9584 0 SS4END[7]
rlabel metal2 29302 8938 29302 8938 0 SS4END[8]
rlabel metal2 29578 8904 29578 8904 0 SS4END[9]
rlabel metal2 1518 1772 1518 1772 0 UserCLK
rlabel metal1 31556 8602 31556 8602 0 UserCLKo
rlabel metal1 36202 2312 36202 2312 0 net1
rlabel metal2 19090 6256 19090 6256 0 net10
rlabel metal2 14214 8908 14214 8908 0 net100
rlabel metal2 18446 7072 18446 7072 0 net101
rlabel metal3 18860 6664 18860 6664 0 net102
rlabel metal1 17894 8330 17894 8330 0 net103
rlabel metal1 30084 7174 30084 7174 0 net104
rlabel metal2 23046 6086 23046 6086 0 net105
rlabel metal2 37490 6562 37490 6562 0 net11
rlabel metal1 36294 2380 36294 2380 0 net12
rlabel metal1 21206 7208 21206 7208 0 net13
rlabel metal1 20562 6664 20562 6664 0 net14
rlabel metal2 34730 6358 34730 6358 0 net15
rlabel metal1 20838 7276 20838 7276 0 net16
rlabel metal2 35190 7038 35190 7038 0 net17
rlabel metal2 38226 8704 38226 8704 0 net18
rlabel metal2 37490 7684 37490 7684 0 net19
rlabel metal2 33810 3791 33810 3791 0 net2
rlabel metal2 22034 7480 22034 7480 0 net20
rlabel metal2 21482 7038 21482 7038 0 net21
rlabel metal2 21022 7191 21022 7191 0 net22
rlabel metal1 21758 4148 21758 4148 0 net23
rlabel metal1 21114 7276 21114 7276 0 net24
rlabel metal2 37582 6494 37582 6494 0 net25
rlabel metal2 18906 3264 18906 3264 0 net26
rlabel metal2 16882 3196 16882 3196 0 net27
rlabel metal2 35006 2176 35006 2176 0 net28
rlabel metal2 37858 3366 37858 3366 0 net29
rlabel metal1 38226 4080 38226 4080 0 net3
rlabel metal1 21482 4012 21482 4012 0 net30
rlabel metal1 34799 3502 34799 3502 0 net31
rlabel metal2 17250 3536 17250 3536 0 net32
rlabel metal2 16330 3468 16330 3468 0 net33
rlabel metal2 35466 6732 35466 6732 0 net34
rlabel metal2 32798 6868 32798 6868 0 net35
rlabel metal2 35834 8738 35834 8738 0 net36
rlabel metal2 36018 7446 36018 7446 0 net37
rlabel metal2 32890 6851 32890 6851 0 net38
rlabel metal1 34224 5814 34224 5814 0 net39
rlabel metal1 21574 4488 21574 4488 0 net4
rlabel metal1 35650 5882 35650 5882 0 net40
rlabel metal1 36708 5814 36708 5814 0 net41
rlabel metal2 37398 7174 37398 7174 0 net42
rlabel metal2 37122 6868 37122 6868 0 net43
rlabel metal2 15410 4063 15410 4063 0 net44
rlabel metal2 20654 3400 20654 3400 0 net45
rlabel metal2 19642 3434 19642 3434 0 net46
rlabel metal2 31878 5916 31878 5916 0 net47
rlabel metal1 33994 8432 33994 8432 0 net48
rlabel metal2 32430 5746 32430 5746 0 net49
rlabel metal1 38226 4624 38226 4624 0 net5
rlabel metal2 31786 7429 31786 7429 0 net50
rlabel metal2 34546 4403 34546 4403 0 net51
rlabel metal2 34914 8806 34914 8806 0 net52
rlabel metal1 6486 7242 6486 7242 0 net53
rlabel metal1 6486 7514 6486 7514 0 net54
rlabel metal1 5428 7514 5428 7514 0 net55
rlabel metal1 4646 7514 4646 7514 0 net56
rlabel metal2 10258 7361 10258 7361 0 net57
rlabel metal1 8280 6630 8280 6630 0 net58
rlabel metal1 6256 6086 6256 6086 0 net59
rlabel metal1 34799 5202 34799 5202 0 net6
rlabel metal1 7682 7480 7682 7480 0 net60
rlabel metal1 7038 7514 7038 7514 0 net61
rlabel metal2 6026 7684 6026 7684 0 net62
rlabel metal1 5888 6630 5888 6630 0 net63
rlabel metal1 5658 7514 5658 7514 0 net64
rlabel metal2 7130 7021 7130 7021 0 net65
rlabel metal2 9614 7378 9614 7378 0 net66
rlabel metal1 9246 6970 9246 6970 0 net67
rlabel metal1 9384 6630 9384 6630 0 net68
rlabel metal1 9016 6902 9016 6902 0 net69
rlabel metal2 18170 5950 18170 5950 0 net7
rlabel metal2 8326 7412 8326 7412 0 net70
rlabel metal1 7820 6630 7820 6630 0 net71
rlabel metal2 7590 7514 7590 7514 0 net72
rlabel metal2 16790 7718 16790 7718 0 net73
rlabel metal2 11270 7854 11270 7854 0 net74
rlabel metal2 11730 7140 11730 7140 0 net75
rlabel metal2 11822 7548 11822 7548 0 net76
rlabel metal2 12282 7412 12282 7412 0 net77
rlabel metal1 14168 6630 14168 6630 0 net78
rlabel metal1 13984 7242 13984 7242 0 net79
rlabel metal1 19734 6868 19734 6868 0 net8
rlabel metal2 17066 8296 17066 8296 0 net80
rlabel metal1 15824 7514 15824 7514 0 net81
rlabel metal1 15410 7480 15410 7480 0 net82
rlabel metal1 14904 7514 14904 7514 0 net83
rlabel metal2 10074 7684 10074 7684 0 net84
rlabel metal2 11086 7718 11086 7718 0 net85
rlabel metal1 14398 6868 14398 6868 0 net86
rlabel metal1 12926 6732 12926 6732 0 net87
rlabel metal1 13110 6868 13110 6868 0 net88
rlabel metal2 12834 8670 12834 8670 0 net89
rlabel metal1 38226 5712 38226 5712 0 net9
rlabel metal2 15686 8840 15686 8840 0 net90
rlabel metal2 15962 8874 15962 8874 0 net91
rlabel metal2 16146 8908 16146 8908 0 net92
rlabel metal1 28290 6630 28290 6630 0 net93
rlabel metal1 19849 8466 19849 8466 0 net94
rlabel metal1 25898 6630 25898 6630 0 net95
rlabel metal2 25438 6392 25438 6392 0 net96
rlabel metal3 17572 6392 17572 6392 0 net97
rlabel metal2 17710 6528 17710 6528 0 net98
rlabel metal2 16146 7055 16146 7055 0 net99
<< properties >>
string FIXED_BBOX 0 0 39928 11152
<< end >>
