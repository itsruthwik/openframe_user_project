* NGSPICE file created from W_term_single.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

.subckt W_term_single E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E2BEG[0] E2BEG[1] E2BEG[2]
+ E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3]
+ E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1] E6BEG[2]
+ E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] EE4BEG[0] EE4BEG[10]
+ EE4BEG[11] EE4BEG[12] EE4BEG[13] EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3]
+ EE4BEG[4] EE4BEG[5] EE4BEG[6] EE4BEG[7] EE4BEG[8] EE4BEG[9] FrameData[0] FrameData[10]
+ FrameData[11] FrameData[12] FrameData[13] FrameData[14] FrameData[15] FrameData[16]
+ FrameData[17] FrameData[18] FrameData[19] FrameData[1] FrameData[20] FrameData[21]
+ FrameData[22] FrameData[23] FrameData[24] FrameData[25] FrameData[26] FrameData[27]
+ FrameData[28] FrameData[29] FrameData[2] FrameData[30] FrameData[31] FrameData[3]
+ FrameData[4] FrameData[5] FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0]
+ FrameData_O[10] FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14]
+ FrameData_O[15] FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19]
+ FrameData_O[1] FrameData_O[20] FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24]
+ FrameData_O[25] FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29]
+ FrameData_O[2] FrameData_O[30] FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5]
+ FrameData_O[6] FrameData_O[7] FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10]
+ FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14] FrameStrobe[15]
+ FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2]
+ FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8]
+ FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12]
+ FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17]
+ FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3]
+ FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8]
+ FrameStrobe_O[9] UserCLK UserCLKo VGND VPWR W1END[0] W1END[1] W1END[2] W1END[3]
+ W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0]
+ W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6] W2MID[7] W6END[0] W6END[10]
+ W6END[11] W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8]
+ W6END[9] WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15]
+ WW4END[1] WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8]
+ WW4END[9]
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_062_ FrameData[14] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_1
XFILLER_48_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_045_ WW4END[2] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_028_ W6END[3] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XANTENNA_5 FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput64 net64 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput53 net53 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
Xoutput31 net31 VGND VGND VPWR VPWR E6BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_31_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput7 net7 VGND VGND VPWR VPWR E2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput20 net20 VGND VGND VPWR VPWR E2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput42 net42 VGND VGND VPWR VPWR EE4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput86 net86 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput97 net97 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
XFILLER_56_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_061_ FrameData[13] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
XFILLER_48_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_044_ WW4END[3] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_6 FrameStrobe[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_027_ W6END[4] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_44_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput87 net87 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput98 net98 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
Xoutput65 net65 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput54 net54 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput76 net76 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
Xoutput32 net32 VGND VGND VPWR VPWR E6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput10 net10 VGND VGND VPWR VPWR E2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput8 net8 VGND VGND VPWR VPWR E2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput43 net43 VGND VGND VPWR VPWR EE4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VPWR VPWR E6BEG[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_73_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_060_ FrameData[12] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_043_ WW4END[4] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_026_ W6END[5] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 W2END[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput88 net88 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput99 net99 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput66 net66 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput55 net55 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput77 net77 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VPWR VPWR E6BEG[10] sky130_fd_sc_hd__buf_2
Xoutput9 net9 VGND VGND VPWR VPWR E2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR E2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput33 net33 VGND VGND VPWR VPWR EE4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput44 net44 VGND VGND VPWR VPWR EE4BEG[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_73_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_009_ W2MID[2] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_042_ WW4END[5] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 WW4END[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_025_ W6END[6] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput23 net23 VGND VGND VPWR VPWR E6BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput12 net12 VGND VGND VPWR VPWR E2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput34 net34 VGND VGND VPWR VPWR EE4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput89 net89 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput56 net56 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput78 net78 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
XFILLER_56_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput45 net45 VGND VGND VPWR VPWR EE4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_008_ W2MID[3] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_64_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_041_ WW4END[6] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 FrameStrobe[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_024_ W6END[7] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput57 net57 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput13 net13 VGND VGND VPWR VPWR E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR EE4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput35 net35 VGND VGND VPWR VPWR EE4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput24 net24 VGND VGND VPWR VPWR E6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput68 net68 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput79 net79 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_007_ W2MID[4] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_040_ WW4END[7] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_023_ W6END[8] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput69 net69 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput58 net58 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR E2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VGND VGND VPWR VPWR EE4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput36 net36 VGND VGND VPWR VPWR EE4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput25 net25 VGND VGND VPWR VPWR E6BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_006_ W2MID[5] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_099_ FrameStrobe[19] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_022_ W6END[9] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput59 net59 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR E2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput48 net48 VGND VGND VPWR VPWR EE4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput37 net37 VGND VGND VPWR VPWR EE4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput26 net26 VGND VGND VPWR VPWR E6BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_005_ W2MID[6] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_098_ FrameStrobe[18] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_1
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_021_ W6END[10] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput49 net49 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VPWR VPWR E2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput38 net38 VGND VGND VPWR VPWR EE4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR E6BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_004_ W2MID[7] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_097_ FrameStrobe[17] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_1
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_020_ W6END[11] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput17 net17 VGND VGND VPWR VPWR E2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput39 net39 VGND VGND VPWR VPWR EE4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput28 net28 VGND VGND VPWR VPWR E6BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_003_ W1END[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_096_ FrameStrobe[16] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_1
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_079_ FrameData[31] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput18 net18 VGND VGND VPWR VPWR E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput29 net29 VGND VGND VPWR VPWR E6BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_56_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_002_ W1END[1] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_095_ FrameStrobe[15] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
XFILLER_40_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_078_ FrameData[30] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR E2BEGb[6] sky130_fd_sc_hd__buf_2
XFILLER_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_001_ W1END[2] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_094_ FrameStrobe[14] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_1
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_077_ FrameData[29] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_32_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_000_ W1END[3] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_093_ FrameStrobe[13] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_076_ FrameData[28] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_29_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ FrameData[11] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_1
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_092_ FrameStrobe[12] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_1
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_075_ FrameData[27] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ FrameData[10] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_091_ FrameStrobe[11] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
XFILLER_40_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_074_ FrameData[26] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_057_ FrameData[9] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_090_ FrameStrobe[10] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_1
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_073_ FrameData[25] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_056_ FrameData[8] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_1
XFILLER_23_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_039_ WW4END[8] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
XFILLER_27_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_072_ FrameData[24] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_055_ FrameData[7] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_038_ WW4END[9] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_44_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_071_ FrameData[23] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_054_ FrameData[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_037_ WW4END[10] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_070_ FrameData[22] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_053_ FrameData[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_036_ WW4END[11] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_019_ W2END[0] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_052_ FrameData[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_035_ WW4END[12] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_018_ W2END[1] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_051_ FrameData[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_034_ WW4END[13] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_017_ W2END[2] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput100 net100 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_050_ FrameData[2] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_033_ WW4END[14] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_016_ W2END[3] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
XFILLER_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput101 net101 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
XFILLER_46_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_032_ WW4END[15] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_015_ W2END[4] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_031_ W6END[0] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
X_100_ UserCLK VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
XFILLER_63_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_014_ W2END[5] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_030_ W6END[1] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_013_ W2END[6] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_089_ FrameStrobe[9] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_012_ W2END[7] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ FrameStrobe[8] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_1
XFILLER_40_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_011_ W2MID[0] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_33_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ FrameStrobe[7] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_1
XFILLER_33_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_010_ W2MID[1] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ FrameStrobe[6] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_1
XFILLER_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_069_ FrameData[21] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput90 net90 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_65_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_085_ FrameStrobe[5] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_1
XFILLER_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_068_ FrameData[20] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput1 net1 VGND VGND VPWR VPWR E1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_49_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput91 net91 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput80 net80 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_084_ FrameStrobe[4] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_1
XFILLER_33_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_067_ FrameData[19] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput70 net70 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
XFILLER_63_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput2 net2 VGND VGND VPWR VPWR E1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput92 net92 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput81 net81 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
XFILLER_11_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_083_ FrameStrobe[3] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_066_ FrameData[18] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_1
XFILLER_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_049_ FrameData[1] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 FrameData[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput82 net82 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput93 net93 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput71 net71 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput60 net60 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput3 net3 VGND VGND VPWR VPWR E1BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_082_ FrameStrobe[2] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_1
XFILLER_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_065_ FrameData[17] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_048_ FrameData[0] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_2 FrameStrobe[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput83 net83 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput94 net94 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput61 net61 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput50 net50 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
Xoutput4 net4 VGND VGND VPWR VPWR E1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_081_ FrameStrobe[1] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_064_ FrameData[16] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_047_ WW4END[0] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_3 FrameStrobe[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput5 net5 VGND VGND VPWR VPWR E2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput84 net84 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput95 net95 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput73 net73 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput62 net62 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
Xoutput51 net51 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput40 net40 VGND VGND VPWR VPWR EE4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_080_ FrameStrobe[0] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_063_ FrameData[15] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_046_ WW4END[1] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_029_ W6END[2] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
XANTENNA_4 FrameStrobe[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput52 net52 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
XFILLER_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput6 net6 VGND VGND VPWR VPWR E2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput41 net41 VGND VGND VPWR VPWR EE4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput30 net30 VGND VGND VPWR VPWR E6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput85 net85 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput96 net96 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput63 net63 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput74 net74 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
.ends

