module eFPGA_Config (CLK,
    ComActive,
    ConfigWriteStrobe,
    LongFrameStrobe,
    ReceiveLED,
    Rx,
    SelfWriteStrobe,
    resetn,
    s_clk,
    s_data,
    vccd1,
    vssd1,
    ConfigWriteData,
    FrameAddressRegister,
    RowSelect,
    SelfWriteData);
 input CLK;
 output ComActive;
 output ConfigWriteStrobe;
 output LongFrameStrobe;
 output ReceiveLED;
 input Rx;
 input SelfWriteStrobe;
 input resetn;
 input s_clk;
 input s_data;
 input vccd1;
 input vssd1;
 output [31:0] ConfigWriteData;
 output [31:0] FrameAddressRegister;
 output [4:0] RowSelect;
 input [31:0] SelfWriteData;

 wire \ConfigFSM_inst.FSM_Reset ;
 wire \ConfigFSM_inst.FrameAddressRegister[0] ;
 wire \ConfigFSM_inst.FrameAddressRegister[10] ;
 wire \ConfigFSM_inst.FrameAddressRegister[11] ;
 wire \ConfigFSM_inst.FrameAddressRegister[12] ;
 wire \ConfigFSM_inst.FrameAddressRegister[13] ;
 wire \ConfigFSM_inst.FrameAddressRegister[14] ;
 wire \ConfigFSM_inst.FrameAddressRegister[15] ;
 wire \ConfigFSM_inst.FrameAddressRegister[16] ;
 wire \ConfigFSM_inst.FrameAddressRegister[17] ;
 wire \ConfigFSM_inst.FrameAddressRegister[18] ;
 wire \ConfigFSM_inst.FrameAddressRegister[19] ;
 wire \ConfigFSM_inst.FrameAddressRegister[1] ;
 wire \ConfigFSM_inst.FrameAddressRegister[21] ;
 wire \ConfigFSM_inst.FrameAddressRegister[22] ;
 wire \ConfigFSM_inst.FrameAddressRegister[23] ;
 wire \ConfigFSM_inst.FrameAddressRegister[24] ;
 wire \ConfigFSM_inst.FrameAddressRegister[25] ;
 wire \ConfigFSM_inst.FrameAddressRegister[26] ;
 wire \ConfigFSM_inst.FrameAddressRegister[27] ;
 wire \ConfigFSM_inst.FrameAddressRegister[28] ;
 wire \ConfigFSM_inst.FrameAddressRegister[29] ;
 wire \ConfigFSM_inst.FrameAddressRegister[2] ;
 wire \ConfigFSM_inst.FrameAddressRegister[30] ;
 wire \ConfigFSM_inst.FrameAddressRegister[31] ;
 wire \ConfigFSM_inst.FrameAddressRegister[3] ;
 wire \ConfigFSM_inst.FrameAddressRegister[4] ;
 wire \ConfigFSM_inst.FrameAddressRegister[5] ;
 wire \ConfigFSM_inst.FrameAddressRegister[6] ;
 wire \ConfigFSM_inst.FrameAddressRegister[7] ;
 wire \ConfigFSM_inst.FrameAddressRegister[8] ;
 wire \ConfigFSM_inst.FrameAddressRegister[9] ;
 wire \ConfigFSM_inst.FrameShiftState[0] ;
 wire \ConfigFSM_inst.FrameShiftState[1] ;
 wire \ConfigFSM_inst.FrameShiftState[2] ;
 wire \ConfigFSM_inst.FrameShiftState[3] ;
 wire \ConfigFSM_inst.FrameShiftState[4] ;
 wire \ConfigFSM_inst.FrameStrobe ;
 wire \ConfigFSM_inst.RowSelect[0] ;
 wire \ConfigFSM_inst.RowSelect[1] ;
 wire \ConfigFSM_inst.RowSelect[2] ;
 wire \ConfigFSM_inst.RowSelect[3] ;
 wire \ConfigFSM_inst.RowSelect[4] ;
 wire \ConfigFSM_inst.WriteData[0] ;
 wire \ConfigFSM_inst.WriteData[10] ;
 wire \ConfigFSM_inst.WriteData[11] ;
 wire \ConfigFSM_inst.WriteData[12] ;
 wire \ConfigFSM_inst.WriteData[13] ;
 wire \ConfigFSM_inst.WriteData[14] ;
 wire \ConfigFSM_inst.WriteData[15] ;
 wire \ConfigFSM_inst.WriteData[16] ;
 wire \ConfigFSM_inst.WriteData[17] ;
 wire \ConfigFSM_inst.WriteData[18] ;
 wire \ConfigFSM_inst.WriteData[19] ;
 wire \ConfigFSM_inst.WriteData[1] ;
 wire \ConfigFSM_inst.WriteData[20] ;
 wire \ConfigFSM_inst.WriteData[21] ;
 wire \ConfigFSM_inst.WriteData[22] ;
 wire \ConfigFSM_inst.WriteData[23] ;
 wire \ConfigFSM_inst.WriteData[24] ;
 wire \ConfigFSM_inst.WriteData[25] ;
 wire \ConfigFSM_inst.WriteData[26] ;
 wire \ConfigFSM_inst.WriteData[27] ;
 wire \ConfigFSM_inst.WriteData[28] ;
 wire \ConfigFSM_inst.WriteData[29] ;
 wire \ConfigFSM_inst.WriteData[2] ;
 wire \ConfigFSM_inst.WriteData[30] ;
 wire \ConfigFSM_inst.WriteData[31] ;
 wire \ConfigFSM_inst.WriteData[3] ;
 wire \ConfigFSM_inst.WriteData[4] ;
 wire \ConfigFSM_inst.WriteData[5] ;
 wire \ConfigFSM_inst.WriteData[6] ;
 wire \ConfigFSM_inst.WriteData[7] ;
 wire \ConfigFSM_inst.WriteData[8] ;
 wire \ConfigFSM_inst.WriteData[9] ;
 wire \ConfigFSM_inst._000_ ;
 wire \ConfigFSM_inst._001_ ;
 wire \ConfigFSM_inst._002_ ;
 wire \ConfigFSM_inst._003_ ;
 wire \ConfigFSM_inst._004_ ;
 wire \ConfigFSM_inst._005_ ;
 wire \ConfigFSM_inst._006_ ;
 wire \ConfigFSM_inst._007_ ;
 wire \ConfigFSM_inst._008_ ;
 wire \ConfigFSM_inst._009_ ;
 wire \ConfigFSM_inst._010_ ;
 wire \ConfigFSM_inst._011_ ;
 wire \ConfigFSM_inst._012_ ;
 wire \ConfigFSM_inst._013_ ;
 wire \ConfigFSM_inst._014_ ;
 wire \ConfigFSM_inst._015_ ;
 wire \ConfigFSM_inst._016_ ;
 wire \ConfigFSM_inst._017_ ;
 wire \ConfigFSM_inst._018_ ;
 wire \ConfigFSM_inst._019_ ;
 wire \ConfigFSM_inst._020_ ;
 wire \ConfigFSM_inst._021_ ;
 wire \ConfigFSM_inst._022_ ;
 wire \ConfigFSM_inst._023_ ;
 wire \ConfigFSM_inst._024_ ;
 wire \ConfigFSM_inst._025_ ;
 wire \ConfigFSM_inst._026_ ;
 wire \ConfigFSM_inst._027_ ;
 wire \ConfigFSM_inst._028_ ;
 wire \ConfigFSM_inst._029_ ;
 wire \ConfigFSM_inst._030_ ;
 wire \ConfigFSM_inst._031_ ;
 wire \ConfigFSM_inst._032_ ;
 wire \ConfigFSM_inst._033_ ;
 wire \ConfigFSM_inst._034_ ;
 wire \ConfigFSM_inst._035_ ;
 wire \ConfigFSM_inst._036_ ;
 wire \ConfigFSM_inst._037_ ;
 wire \ConfigFSM_inst._038_ ;
 wire \ConfigFSM_inst._039_ ;
 wire \ConfigFSM_inst._040_ ;
 wire \ConfigFSM_inst._041_ ;
 wire \ConfigFSM_inst._042_ ;
 wire \ConfigFSM_inst._043_ ;
 wire \ConfigFSM_inst._044_ ;
 wire \ConfigFSM_inst._045_ ;
 wire \ConfigFSM_inst._046_ ;
 wire \ConfigFSM_inst._047_ ;
 wire \ConfigFSM_inst._048_ ;
 wire \ConfigFSM_inst._049_ ;
 wire \ConfigFSM_inst._050_ ;
 wire \ConfigFSM_inst._051_ ;
 wire \ConfigFSM_inst._052_ ;
 wire \ConfigFSM_inst._053_ ;
 wire \ConfigFSM_inst._054_ ;
 wire \ConfigFSM_inst._055_ ;
 wire \ConfigFSM_inst._056_ ;
 wire \ConfigFSM_inst._057_ ;
 wire \ConfigFSM_inst._058_ ;
 wire \ConfigFSM_inst._059_ ;
 wire \ConfigFSM_inst._060_ ;
 wire \ConfigFSM_inst._061_ ;
 wire \ConfigFSM_inst._062_ ;
 wire \ConfigFSM_inst._063_ ;
 wire \ConfigFSM_inst._064_ ;
 wire \ConfigFSM_inst._065_ ;
 wire \ConfigFSM_inst._066_ ;
 wire \ConfigFSM_inst._067_ ;
 wire \ConfigFSM_inst._068_ ;
 wire \ConfigFSM_inst._069_ ;
 wire \ConfigFSM_inst._070_ ;
 wire \ConfigFSM_inst._071_ ;
 wire \ConfigFSM_inst._072_ ;
 wire \ConfigFSM_inst._073_ ;
 wire \ConfigFSM_inst._074_ ;
 wire \ConfigFSM_inst._075_ ;
 wire \ConfigFSM_inst._076_ ;
 wire \ConfigFSM_inst._077_ ;
 wire \ConfigFSM_inst._078_ ;
 wire \ConfigFSM_inst._079_ ;
 wire \ConfigFSM_inst._080_ ;
 wire \ConfigFSM_inst._081_ ;
 wire \ConfigFSM_inst._082_ ;
 wire \ConfigFSM_inst._083_ ;
 wire \ConfigFSM_inst._084_ ;
 wire \ConfigFSM_inst._085_ ;
 wire \ConfigFSM_inst._086_ ;
 wire \ConfigFSM_inst._087_ ;
 wire \ConfigFSM_inst._088_ ;
 wire \ConfigFSM_inst._089_ ;
 wire \ConfigFSM_inst._090_ ;
 wire \ConfigFSM_inst._091_ ;
 wire \ConfigFSM_inst._092_ ;
 wire \ConfigFSM_inst._093_ ;
 wire \ConfigFSM_inst._094_ ;
 wire \ConfigFSM_inst._095_ ;
 wire \ConfigFSM_inst._096_ ;
 wire \ConfigFSM_inst._097_ ;
 wire \ConfigFSM_inst._098_ ;
 wire \ConfigFSM_inst._099_ ;
 wire \ConfigFSM_inst._100_ ;
 wire \ConfigFSM_inst._101_ ;
 wire \ConfigFSM_inst._102_ ;
 wire \ConfigFSM_inst._103_ ;
 wire \ConfigFSM_inst._104_ ;
 wire \ConfigFSM_inst._105_ ;
 wire \ConfigFSM_inst._106_ ;
 wire \ConfigFSM_inst._107_ ;
 wire \ConfigFSM_inst._108_ ;
 wire \ConfigFSM_inst._109_ ;
 wire \ConfigFSM_inst._110_ ;
 wire \ConfigFSM_inst._111_ ;
 wire \ConfigFSM_inst._112_ ;
 wire \ConfigFSM_inst._113_ ;
 wire \ConfigFSM_inst._114_ ;
 wire \ConfigFSM_inst._115_ ;
 wire \ConfigFSM_inst._116_ ;
 wire \ConfigFSM_inst._117_ ;
 wire \ConfigFSM_inst._118_ ;
 wire \ConfigFSM_inst._119_ ;
 wire \ConfigFSM_inst.oldFrameStrobe ;
 wire \ConfigFSM_inst.old_reset ;
 wire \ConfigFSM_inst.state[0] ;
 wire \ConfigFSM_inst.state[1] ;
 wire \ConfigFSM_inst.state[2] ;
 wire \INST_config_UART.ByteWriteStrobe ;
 wire \INST_config_UART.CRCReg[0] ;
 wire \INST_config_UART.CRCReg[10] ;
 wire \INST_config_UART.CRCReg[11] ;
 wire \INST_config_UART.CRCReg[12] ;
 wire \INST_config_UART.CRCReg[13] ;
 wire \INST_config_UART.CRCReg[14] ;
 wire \INST_config_UART.CRCReg[15] ;
 wire \INST_config_UART.CRCReg[16] ;
 wire \INST_config_UART.CRCReg[17] ;
 wire \INST_config_UART.CRCReg[18] ;
 wire \INST_config_UART.CRCReg[19] ;
 wire \INST_config_UART.CRCReg[1] ;
 wire \INST_config_UART.CRCReg[2] ;
 wire \INST_config_UART.CRCReg[3] ;
 wire \INST_config_UART.CRCReg[4] ;
 wire \INST_config_UART.CRCReg[5] ;
 wire \INST_config_UART.CRCReg[6] ;
 wire \INST_config_UART.CRCReg[7] ;
 wire \INST_config_UART.CRCReg[8] ;
 wire \INST_config_UART.CRCReg[9] ;
 wire \INST_config_UART.ComCount[0] ;
 wire \INST_config_UART.ComCount[10] ;
 wire \INST_config_UART.ComCount[11] ;
 wire \INST_config_UART.ComCount[1] ;
 wire \INST_config_UART.ComCount[2] ;
 wire \INST_config_UART.ComCount[3] ;
 wire \INST_config_UART.ComCount[4] ;
 wire \INST_config_UART.ComCount[5] ;
 wire \INST_config_UART.ComCount[6] ;
 wire \INST_config_UART.ComCount[7] ;
 wire \INST_config_UART.ComCount[8] ;
 wire \INST_config_UART.ComCount[9] ;
 wire \INST_config_UART.ComState[0] ;
 wire \INST_config_UART.ComState[10] ;
 wire \INST_config_UART.ComState[1] ;
 wire \INST_config_UART.ComState[2] ;
 wire \INST_config_UART.ComState[3] ;
 wire \INST_config_UART.ComState[4] ;
 wire \INST_config_UART.ComState[5] ;
 wire \INST_config_UART.ComState[6] ;
 wire \INST_config_UART.ComState[7] ;
 wire \INST_config_UART.ComState[8] ;
 wire \INST_config_UART.ComState[9] ;
 wire \INST_config_UART.ComTick ;
 wire \INST_config_UART.Command[0] ;
 wire \INST_config_UART.Command[1] ;
 wire \INST_config_UART.Command[2] ;
 wire \INST_config_UART.Command[3] ;
 wire \INST_config_UART.Command[4] ;
 wire \INST_config_UART.Command[5] ;
 wire \INST_config_UART.Command[6] ;
 wire \INST_config_UART.Command[7] ;
 wire \INST_config_UART.Data_Reg[0] ;
 wire \INST_config_UART.Data_Reg[1] ;
 wire \INST_config_UART.Data_Reg[2] ;
 wire \INST_config_UART.Data_Reg[3] ;
 wire \INST_config_UART.Data_Reg[4] ;
 wire \INST_config_UART.Data_Reg[5] ;
 wire \INST_config_UART.Data_Reg[6] ;
 wire \INST_config_UART.Data_Reg[7] ;
 wire \INST_config_UART.GetWordState[0] ;
 wire \INST_config_UART.GetWordState[1] ;
 wire \INST_config_UART.GetWordState[2] ;
 wire \INST_config_UART.GetWordState[3] ;
 wire \INST_config_UART.HexData[0] ;
 wire \INST_config_UART.HexData[1] ;
 wire \INST_config_UART.HexData[2] ;
 wire \INST_config_UART.HexData[3] ;
 wire \INST_config_UART.HexData[4] ;
 wire \INST_config_UART.HexData[5] ;
 wire \INST_config_UART.HexData[6] ;
 wire \INST_config_UART.HexData[7] ;
 wire \INST_config_UART.HexWriteStrobe ;
 wire \INST_config_UART.HighReg[0] ;
 wire \INST_config_UART.HighReg[1] ;
 wire \INST_config_UART.HighReg[2] ;
 wire \INST_config_UART.HighReg[3] ;
 wire \INST_config_UART.ID_Reg[0] ;
 wire \INST_config_UART.ID_Reg[10] ;
 wire \INST_config_UART.ID_Reg[11] ;
 wire \INST_config_UART.ID_Reg[12] ;
 wire \INST_config_UART.ID_Reg[13] ;
 wire \INST_config_UART.ID_Reg[14] ;
 wire \INST_config_UART.ID_Reg[15] ;
 wire \INST_config_UART.ID_Reg[16] ;
 wire \INST_config_UART.ID_Reg[17] ;
 wire \INST_config_UART.ID_Reg[18] ;
 wire \INST_config_UART.ID_Reg[19] ;
 wire \INST_config_UART.ID_Reg[1] ;
 wire \INST_config_UART.ID_Reg[20] ;
 wire \INST_config_UART.ID_Reg[21] ;
 wire \INST_config_UART.ID_Reg[22] ;
 wire \INST_config_UART.ID_Reg[23] ;
 wire \INST_config_UART.ID_Reg[2] ;
 wire \INST_config_UART.ID_Reg[3] ;
 wire \INST_config_UART.ID_Reg[4] ;
 wire \INST_config_UART.ID_Reg[5] ;
 wire \INST_config_UART.ID_Reg[6] ;
 wire \INST_config_UART.ID_Reg[7] ;
 wire \INST_config_UART.ID_Reg[8] ;
 wire \INST_config_UART.ID_Reg[9] ;
 wire \INST_config_UART.LocalWriteStrobe ;
 wire \INST_config_UART.PresentState[0] ;
 wire \INST_config_UART.PresentState[1] ;
 wire \INST_config_UART.PresentState[2] ;
 wire \INST_config_UART.PresentState[4] ;
 wire \INST_config_UART.PresentState[5] ;
 wire \INST_config_UART.PresentState[6] ;
 wire \INST_config_UART.ReceiveLED ;
 wire \INST_config_UART.ReceiveState ;
 wire \INST_config_UART.ReceivedWord[0] ;
 wire \INST_config_UART.ReceivedWord[1] ;
 wire \INST_config_UART.ReceivedWord[2] ;
 wire \INST_config_UART.ReceivedWord[3] ;
 wire \INST_config_UART.ReceivedWord[4] ;
 wire \INST_config_UART.ReceivedWord[5] ;
 wire \INST_config_UART.ReceivedWord[6] ;
 wire \INST_config_UART.ReceivedWord[7] ;
 wire \INST_config_UART.RxLocal ;
 wire \INST_config_UART.TimeToSend ;
 wire \INST_config_UART.TimeToSendCounter[0] ;
 wire \INST_config_UART.TimeToSendCounter[10] ;
 wire \INST_config_UART.TimeToSendCounter[11] ;
 wire \INST_config_UART.TimeToSendCounter[12] ;
 wire \INST_config_UART.TimeToSendCounter[13] ;
 wire \INST_config_UART.TimeToSendCounter[14] ;
 wire \INST_config_UART.TimeToSendCounter[1] ;
 wire \INST_config_UART.TimeToSendCounter[2] ;
 wire \INST_config_UART.TimeToSendCounter[3] ;
 wire \INST_config_UART.TimeToSendCounter[4] ;
 wire \INST_config_UART.TimeToSendCounter[5] ;
 wire \INST_config_UART.TimeToSendCounter[6] ;
 wire \INST_config_UART.TimeToSendCounter[7] ;
 wire \INST_config_UART.TimeToSendCounter[8] ;
 wire \INST_config_UART.TimeToSendCounter[9] ;
 wire \INST_config_UART.WriteData[0] ;
 wire \INST_config_UART.WriteData[10] ;
 wire \INST_config_UART.WriteData[11] ;
 wire \INST_config_UART.WriteData[12] ;
 wire \INST_config_UART.WriteData[13] ;
 wire \INST_config_UART.WriteData[14] ;
 wire \INST_config_UART.WriteData[15] ;
 wire \INST_config_UART.WriteData[16] ;
 wire \INST_config_UART.WriteData[17] ;
 wire \INST_config_UART.WriteData[18] ;
 wire \INST_config_UART.WriteData[19] ;
 wire \INST_config_UART.WriteData[1] ;
 wire \INST_config_UART.WriteData[20] ;
 wire \INST_config_UART.WriteData[21] ;
 wire \INST_config_UART.WriteData[22] ;
 wire \INST_config_UART.WriteData[23] ;
 wire \INST_config_UART.WriteData[24] ;
 wire \INST_config_UART.WriteData[25] ;
 wire \INST_config_UART.WriteData[26] ;
 wire \INST_config_UART.WriteData[27] ;
 wire \INST_config_UART.WriteData[28] ;
 wire \INST_config_UART.WriteData[29] ;
 wire \INST_config_UART.WriteData[2] ;
 wire \INST_config_UART.WriteData[30] ;
 wire \INST_config_UART.WriteData[31] ;
 wire \INST_config_UART.WriteData[3] ;
 wire \INST_config_UART.WriteData[4] ;
 wire \INST_config_UART.WriteData[5] ;
 wire \INST_config_UART.WriteData[6] ;
 wire \INST_config_UART.WriteData[7] ;
 wire \INST_config_UART.WriteData[8] ;
 wire \INST_config_UART.WriteData[9] ;
 wire \INST_config_UART.WriteStrobe ;
 wire \INST_config_UART._0000_ ;
 wire \INST_config_UART._0001_ ;
 wire \INST_config_UART._0002_ ;
 wire \INST_config_UART._0003_ ;
 wire \INST_config_UART._0004_ ;
 wire \INST_config_UART._0005_ ;
 wire \INST_config_UART._0006_ ;
 wire \INST_config_UART._0007_ ;
 wire \INST_config_UART._0008_ ;
 wire \INST_config_UART._0009_ ;
 wire \INST_config_UART._0010_ ;
 wire \INST_config_UART._0011_ ;
 wire \INST_config_UART._0012_ ;
 wire \INST_config_UART._0013_ ;
 wire \INST_config_UART._0014_ ;
 wire \INST_config_UART._0015_ ;
 wire \INST_config_UART._0016_ ;
 wire \INST_config_UART._0017_ ;
 wire \INST_config_UART._0018_ ;
 wire \INST_config_UART._0019_ ;
 wire \INST_config_UART._0020_ ;
 wire \INST_config_UART._0021_ ;
 wire \INST_config_UART._0022_ ;
 wire \INST_config_UART._0023_ ;
 wire \INST_config_UART._0024_ ;
 wire \INST_config_UART._0025_ ;
 wire \INST_config_UART._0026_ ;
 wire \INST_config_UART._0027_ ;
 wire \INST_config_UART._0028_ ;
 wire \INST_config_UART._0029_ ;
 wire \INST_config_UART._0030_ ;
 wire \INST_config_UART._0031_ ;
 wire \INST_config_UART._0032_ ;
 wire \INST_config_UART._0033_ ;
 wire \INST_config_UART._0034_ ;
 wire \INST_config_UART._0035_ ;
 wire \INST_config_UART._0036_ ;
 wire \INST_config_UART._0037_ ;
 wire \INST_config_UART._0038_ ;
 wire \INST_config_UART._0039_ ;
 wire \INST_config_UART._0040_ ;
 wire \INST_config_UART._0041_ ;
 wire \INST_config_UART._0042_ ;
 wire \INST_config_UART._0043_ ;
 wire \INST_config_UART._0044_ ;
 wire \INST_config_UART._0045_ ;
 wire \INST_config_UART._0046_ ;
 wire \INST_config_UART._0047_ ;
 wire \INST_config_UART._0048_ ;
 wire \INST_config_UART._0049_ ;
 wire \INST_config_UART._0050_ ;
 wire \INST_config_UART._0051_ ;
 wire \INST_config_UART._0052_ ;
 wire \INST_config_UART._0053_ ;
 wire \INST_config_UART._0054_ ;
 wire \INST_config_UART._0055_ ;
 wire \INST_config_UART._0056_ ;
 wire \INST_config_UART._0057_ ;
 wire \INST_config_UART._0058_ ;
 wire \INST_config_UART._0059_ ;
 wire \INST_config_UART._0060_ ;
 wire \INST_config_UART._0061_ ;
 wire \INST_config_UART._0062_ ;
 wire \INST_config_UART._0063_ ;
 wire \INST_config_UART._0064_ ;
 wire \INST_config_UART._0065_ ;
 wire \INST_config_UART._0066_ ;
 wire \INST_config_UART._0067_ ;
 wire \INST_config_UART._0068_ ;
 wire \INST_config_UART._0069_ ;
 wire \INST_config_UART._0070_ ;
 wire \INST_config_UART._0071_ ;
 wire \INST_config_UART._0072_ ;
 wire \INST_config_UART._0073_ ;
 wire \INST_config_UART._0074_ ;
 wire \INST_config_UART._0075_ ;
 wire \INST_config_UART._0076_ ;
 wire \INST_config_UART._0077_ ;
 wire \INST_config_UART._0078_ ;
 wire \INST_config_UART._0079_ ;
 wire \INST_config_UART._0080_ ;
 wire \INST_config_UART._0081_ ;
 wire \INST_config_UART._0082_ ;
 wire \INST_config_UART._0083_ ;
 wire \INST_config_UART._0084_ ;
 wire \INST_config_UART._0085_ ;
 wire \INST_config_UART._0086_ ;
 wire \INST_config_UART._0087_ ;
 wire \INST_config_UART._0088_ ;
 wire \INST_config_UART._0089_ ;
 wire \INST_config_UART._0090_ ;
 wire \INST_config_UART._0091_ ;
 wire \INST_config_UART._0092_ ;
 wire \INST_config_UART._0093_ ;
 wire \INST_config_UART._0094_ ;
 wire \INST_config_UART._0095_ ;
 wire \INST_config_UART._0096_ ;
 wire \INST_config_UART._0097_ ;
 wire \INST_config_UART._0098_ ;
 wire \INST_config_UART._0099_ ;
 wire \INST_config_UART._0100_ ;
 wire \INST_config_UART._0101_ ;
 wire \INST_config_UART._0102_ ;
 wire \INST_config_UART._0103_ ;
 wire \INST_config_UART._0104_ ;
 wire \INST_config_UART._0105_ ;
 wire \INST_config_UART._0106_ ;
 wire \INST_config_UART._0107_ ;
 wire \INST_config_UART._0108_ ;
 wire \INST_config_UART._0109_ ;
 wire \INST_config_UART._0110_ ;
 wire \INST_config_UART._0111_ ;
 wire \INST_config_UART._0112_ ;
 wire \INST_config_UART._0113_ ;
 wire \INST_config_UART._0114_ ;
 wire \INST_config_UART._0115_ ;
 wire \INST_config_UART._0116_ ;
 wire \INST_config_UART._0117_ ;
 wire \INST_config_UART._0118_ ;
 wire \INST_config_UART._0119_ ;
 wire \INST_config_UART._0120_ ;
 wire \INST_config_UART._0121_ ;
 wire \INST_config_UART._0122_ ;
 wire \INST_config_UART._0123_ ;
 wire \INST_config_UART._0124_ ;
 wire \INST_config_UART._0125_ ;
 wire \INST_config_UART._0126_ ;
 wire \INST_config_UART._0127_ ;
 wire \INST_config_UART._0128_ ;
 wire \INST_config_UART._0129_ ;
 wire \INST_config_UART._0130_ ;
 wire \INST_config_UART._0131_ ;
 wire \INST_config_UART._0132_ ;
 wire \INST_config_UART._0133_ ;
 wire \INST_config_UART._0134_ ;
 wire \INST_config_UART._0135_ ;
 wire \INST_config_UART._0136_ ;
 wire \INST_config_UART._0137_ ;
 wire \INST_config_UART._0138_ ;
 wire \INST_config_UART._0139_ ;
 wire \INST_config_UART._0140_ ;
 wire \INST_config_UART._0141_ ;
 wire \INST_config_UART._0142_ ;
 wire \INST_config_UART._0143_ ;
 wire \INST_config_UART._0144_ ;
 wire \INST_config_UART._0145_ ;
 wire \INST_config_UART._0146_ ;
 wire \INST_config_UART._0147_ ;
 wire \INST_config_UART._0148_ ;
 wire \INST_config_UART._0149_ ;
 wire \INST_config_UART._0150_ ;
 wire \INST_config_UART._0151_ ;
 wire \INST_config_UART._0152_ ;
 wire \INST_config_UART._0153_ ;
 wire \INST_config_UART._0154_ ;
 wire \INST_config_UART._0155_ ;
 wire \INST_config_UART._0156_ ;
 wire \INST_config_UART._0157_ ;
 wire \INST_config_UART._0158_ ;
 wire \INST_config_UART._0159_ ;
 wire \INST_config_UART._0160_ ;
 wire \INST_config_UART._0161_ ;
 wire \INST_config_UART._0162_ ;
 wire \INST_config_UART._0163_ ;
 wire \INST_config_UART._0164_ ;
 wire \INST_config_UART._0165_ ;
 wire \INST_config_UART._0166_ ;
 wire \INST_config_UART._0167_ ;
 wire \INST_config_UART._0168_ ;
 wire \INST_config_UART._0169_ ;
 wire \INST_config_UART._0170_ ;
 wire \INST_config_UART._0171_ ;
 wire \INST_config_UART._0172_ ;
 wire \INST_config_UART._0173_ ;
 wire \INST_config_UART._0174_ ;
 wire \INST_config_UART._0175_ ;
 wire \INST_config_UART._0176_ ;
 wire \INST_config_UART._0177_ ;
 wire \INST_config_UART._0178_ ;
 wire \INST_config_UART._0179_ ;
 wire \INST_config_UART._0180_ ;
 wire \INST_config_UART._0181_ ;
 wire \INST_config_UART._0182_ ;
 wire \INST_config_UART._0183_ ;
 wire \INST_config_UART._0184_ ;
 wire \INST_config_UART._0185_ ;
 wire \INST_config_UART._0186_ ;
 wire \INST_config_UART._0187_ ;
 wire \INST_config_UART._0188_ ;
 wire \INST_config_UART._0189_ ;
 wire \INST_config_UART._0190_ ;
 wire \INST_config_UART._0191_ ;
 wire \INST_config_UART._0192_ ;
 wire \INST_config_UART._0193_ ;
 wire \INST_config_UART._0194_ ;
 wire \INST_config_UART._0195_ ;
 wire \INST_config_UART._0196_ ;
 wire \INST_config_UART._0197_ ;
 wire \INST_config_UART._0198_ ;
 wire \INST_config_UART._0199_ ;
 wire \INST_config_UART._0200_ ;
 wire \INST_config_UART._0201_ ;
 wire \INST_config_UART._0202_ ;
 wire \INST_config_UART._0203_ ;
 wire \INST_config_UART._0204_ ;
 wire \INST_config_UART._0205_ ;
 wire \INST_config_UART._0206_ ;
 wire \INST_config_UART._0207_ ;
 wire \INST_config_UART._0208_ ;
 wire \INST_config_UART._0209_ ;
 wire \INST_config_UART._0210_ ;
 wire \INST_config_UART._0211_ ;
 wire \INST_config_UART._0212_ ;
 wire \INST_config_UART._0213_ ;
 wire \INST_config_UART._0214_ ;
 wire \INST_config_UART._0215_ ;
 wire \INST_config_UART._0216_ ;
 wire \INST_config_UART._0217_ ;
 wire \INST_config_UART._0218_ ;
 wire \INST_config_UART._0219_ ;
 wire \INST_config_UART._0220_ ;
 wire \INST_config_UART._0221_ ;
 wire \INST_config_UART._0222_ ;
 wire \INST_config_UART._0223_ ;
 wire \INST_config_UART._0224_ ;
 wire \INST_config_UART._0225_ ;
 wire \INST_config_UART._0226_ ;
 wire \INST_config_UART._0227_ ;
 wire \INST_config_UART._0228_ ;
 wire \INST_config_UART._0229_ ;
 wire \INST_config_UART._0230_ ;
 wire \INST_config_UART._0231_ ;
 wire \INST_config_UART._0232_ ;
 wire \INST_config_UART._0233_ ;
 wire \INST_config_UART._0234_ ;
 wire \INST_config_UART._0235_ ;
 wire \INST_config_UART._0236_ ;
 wire \INST_config_UART._0237_ ;
 wire \INST_config_UART._0238_ ;
 wire \INST_config_UART._0239_ ;
 wire \INST_config_UART._0240_ ;
 wire \INST_config_UART._0241_ ;
 wire \INST_config_UART._0242_ ;
 wire \INST_config_UART._0243_ ;
 wire \INST_config_UART._0244_ ;
 wire \INST_config_UART._0245_ ;
 wire \INST_config_UART._0246_ ;
 wire \INST_config_UART._0247_ ;
 wire \INST_config_UART._0248_ ;
 wire \INST_config_UART._0249_ ;
 wire \INST_config_UART._0250_ ;
 wire \INST_config_UART._0251_ ;
 wire \INST_config_UART._0252_ ;
 wire \INST_config_UART._0253_ ;
 wire \INST_config_UART._0254_ ;
 wire \INST_config_UART._0255_ ;
 wire \INST_config_UART._0256_ ;
 wire \INST_config_UART._0257_ ;
 wire \INST_config_UART._0258_ ;
 wire \INST_config_UART._0259_ ;
 wire \INST_config_UART._0260_ ;
 wire \INST_config_UART._0261_ ;
 wire \INST_config_UART._0262_ ;
 wire \INST_config_UART._0263_ ;
 wire \INST_config_UART._0264_ ;
 wire \INST_config_UART._0265_ ;
 wire \INST_config_UART._0266_ ;
 wire \INST_config_UART._0267_ ;
 wire \INST_config_UART._0268_ ;
 wire \INST_config_UART._0269_ ;
 wire \INST_config_UART._0270_ ;
 wire \INST_config_UART._0271_ ;
 wire \INST_config_UART._0272_ ;
 wire \INST_config_UART._0273_ ;
 wire \INST_config_UART._0274_ ;
 wire \INST_config_UART._0275_ ;
 wire \INST_config_UART._0276_ ;
 wire \INST_config_UART._0277_ ;
 wire \INST_config_UART._0278_ ;
 wire \INST_config_UART._0279_ ;
 wire \INST_config_UART._0280_ ;
 wire \INST_config_UART._0281_ ;
 wire \INST_config_UART._0282_ ;
 wire \INST_config_UART._0283_ ;
 wire \INST_config_UART._0284_ ;
 wire \INST_config_UART._0285_ ;
 wire \INST_config_UART._0286_ ;
 wire \INST_config_UART._0287_ ;
 wire \INST_config_UART._0288_ ;
 wire \INST_config_UART._0289_ ;
 wire \INST_config_UART._0290_ ;
 wire \INST_config_UART._0291_ ;
 wire \INST_config_UART._0292_ ;
 wire \INST_config_UART._0293_ ;
 wire \INST_config_UART._0294_ ;
 wire \INST_config_UART._0295_ ;
 wire \INST_config_UART._0296_ ;
 wire \INST_config_UART._0297_ ;
 wire \INST_config_UART._0298_ ;
 wire \INST_config_UART._0299_ ;
 wire \INST_config_UART._0300_ ;
 wire \INST_config_UART._0301_ ;
 wire \INST_config_UART._0302_ ;
 wire \INST_config_UART._0303_ ;
 wire \INST_config_UART._0304_ ;
 wire \INST_config_UART._0305_ ;
 wire \INST_config_UART._0306_ ;
 wire \INST_config_UART._0307_ ;
 wire \INST_config_UART._0308_ ;
 wire \INST_config_UART._0309_ ;
 wire \INST_config_UART._0310_ ;
 wire \INST_config_UART._0311_ ;
 wire \INST_config_UART._0312_ ;
 wire \INST_config_UART._0313_ ;
 wire \INST_config_UART._0314_ ;
 wire \INST_config_UART._0315_ ;
 wire \INST_config_UART._0316_ ;
 wire \INST_config_UART._0317_ ;
 wire \INST_config_UART._0318_ ;
 wire \INST_config_UART._0319_ ;
 wire \INST_config_UART._0320_ ;
 wire \INST_config_UART._0321_ ;
 wire \INST_config_UART._0322_ ;
 wire \INST_config_UART._0323_ ;
 wire \INST_config_UART._0324_ ;
 wire \INST_config_UART._0325_ ;
 wire \INST_config_UART._0326_ ;
 wire \INST_config_UART._0327_ ;
 wire \INST_config_UART._0328_ ;
 wire \INST_config_UART._0329_ ;
 wire \INST_config_UART._0330_ ;
 wire \INST_config_UART._0331_ ;
 wire \INST_config_UART._0332_ ;
 wire \INST_config_UART._0333_ ;
 wire \INST_config_UART._0334_ ;
 wire \INST_config_UART._0335_ ;
 wire \INST_config_UART._0336_ ;
 wire \INST_config_UART._0337_ ;
 wire \INST_config_UART._0338_ ;
 wire \INST_config_UART._0339_ ;
 wire \INST_config_UART._0340_ ;
 wire \INST_config_UART._0341_ ;
 wire \INST_config_UART._0342_ ;
 wire \INST_config_UART._0343_ ;
 wire \INST_config_UART._0344_ ;
 wire \INST_config_UART._0345_ ;
 wire \INST_config_UART._0346_ ;
 wire \INST_config_UART._0347_ ;
 wire \INST_config_UART._0348_ ;
 wire \INST_config_UART._0349_ ;
 wire \INST_config_UART._0350_ ;
 wire \INST_config_UART._0351_ ;
 wire \INST_config_UART._0352_ ;
 wire \INST_config_UART._0353_ ;
 wire \INST_config_UART._0354_ ;
 wire \INST_config_UART._0355_ ;
 wire \INST_config_UART._0356_ ;
 wire \INST_config_UART._0357_ ;
 wire \INST_config_UART._0358_ ;
 wire \INST_config_UART._0359_ ;
 wire \INST_config_UART._0360_ ;
 wire \INST_config_UART._0361_ ;
 wire \INST_config_UART._0362_ ;
 wire \INST_config_UART._0363_ ;
 wire \INST_config_UART._0364_ ;
 wire \INST_config_UART._0365_ ;
 wire \INST_config_UART._0366_ ;
 wire \INST_config_UART._0367_ ;
 wire \INST_config_UART._0368_ ;
 wire \INST_config_UART._0369_ ;
 wire \INST_config_UART._0370_ ;
 wire \INST_config_UART._0371_ ;
 wire \INST_config_UART._0372_ ;
 wire \INST_config_UART._0373_ ;
 wire \INST_config_UART._0374_ ;
 wire \INST_config_UART._0375_ ;
 wire \INST_config_UART._0376_ ;
 wire \INST_config_UART._0377_ ;
 wire \INST_config_UART._0378_ ;
 wire \INST_config_UART._0379_ ;
 wire \INST_config_UART._0380_ ;
 wire \INST_config_UART._0381_ ;
 wire \INST_config_UART._0382_ ;
 wire \INST_config_UART._0383_ ;
 wire \INST_config_UART._0384_ ;
 wire \INST_config_UART._0385_ ;
 wire \INST_config_UART._0386_ ;
 wire \INST_config_UART._0387_ ;
 wire \INST_config_UART._0388_ ;
 wire \INST_config_UART._0389_ ;
 wire \INST_config_UART._0390_ ;
 wire \INST_config_UART._0391_ ;
 wire \INST_config_UART._0392_ ;
 wire \INST_config_UART._0393_ ;
 wire \INST_config_UART._0394_ ;
 wire \INST_config_UART._0395_ ;
 wire \INST_config_UART._0396_ ;
 wire \INST_config_UART._0397_ ;
 wire \INST_config_UART._0398_ ;
 wire \INST_config_UART._0399_ ;
 wire \INST_config_UART._0400_ ;
 wire \INST_config_UART._0401_ ;
 wire \INST_config_UART._0402_ ;
 wire \INST_config_UART._0403_ ;
 wire \INST_config_UART._0404_ ;
 wire \INST_config_UART._0405_ ;
 wire \INST_config_UART._0406_ ;
 wire \INST_config_UART._0407_ ;
 wire \INST_config_UART._0408_ ;
 wire \INST_config_UART._0409_ ;
 wire \INST_config_UART._0410_ ;
 wire \INST_config_UART._0411_ ;
 wire \INST_config_UART._0412_ ;
 wire \INST_config_UART._0413_ ;
 wire \INST_config_UART._0414_ ;
 wire \INST_config_UART._0415_ ;
 wire \INST_config_UART._0416_ ;
 wire \INST_config_UART._0417_ ;
 wire \INST_config_UART._0418_ ;
 wire \INST_config_UART._0419_ ;
 wire \INST_config_UART._0420_ ;
 wire \INST_config_UART._0421_ ;
 wire \INST_config_UART._0422_ ;
 wire \INST_config_UART._0423_ ;
 wire \INST_config_UART._0424_ ;
 wire \INST_config_UART._0425_ ;
 wire \INST_config_UART._0426_ ;
 wire \INST_config_UART._0427_ ;
 wire \INST_config_UART._0428_ ;
 wire \INST_config_UART._0429_ ;
 wire \INST_config_UART._0430_ ;
 wire \INST_config_UART._0431_ ;
 wire \INST_config_UART._0432_ ;
 wire \INST_config_UART._0433_ ;
 wire \INST_config_UART._0434_ ;
 wire \INST_config_UART._0435_ ;
 wire \INST_config_UART._0436_ ;
 wire \INST_config_UART._0437_ ;
 wire \INST_config_UART._0438_ ;
 wire \INST_config_UART._0439_ ;
 wire \INST_config_UART._0440_ ;
 wire \INST_config_UART._0441_ ;
 wire \INST_config_UART._0442_ ;
 wire \INST_config_UART._0443_ ;
 wire \INST_config_UART._0444_ ;
 wire \INST_config_UART._0445_ ;
 wire \INST_config_UART._0446_ ;
 wire \INST_config_UART._0447_ ;
 wire \INST_config_UART._0448_ ;
 wire \INST_config_UART._0449_ ;
 wire \INST_config_UART._0450_ ;
 wire \INST_config_UART._0451_ ;
 wire \INST_config_UART._0452_ ;
 wire \INST_config_UART._0453_ ;
 wire \INST_config_UART._0454_ ;
 wire \INST_config_UART._0455_ ;
 wire \INST_config_UART._0456_ ;
 wire \INST_config_UART._0457_ ;
 wire \INST_config_UART._0458_ ;
 wire \INST_config_UART._0459_ ;
 wire \INST_config_UART._0460_ ;
 wire \INST_config_UART._0461_ ;
 wire \INST_config_UART._0462_ ;
 wire \INST_config_UART._0463_ ;
 wire \INST_config_UART._0464_ ;
 wire \INST_config_UART._0465_ ;
 wire \INST_config_UART._0466_ ;
 wire \INST_config_UART._0467_ ;
 wire \INST_config_UART._0468_ ;
 wire \INST_config_UART._0469_ ;
 wire \INST_config_UART._0470_ ;
 wire \INST_config_UART._0471_ ;
 wire \INST_config_UART._0472_ ;
 wire \INST_config_UART._0473_ ;
 wire \INST_config_UART._0474_ ;
 wire \INST_config_UART._0475_ ;
 wire \INST_config_UART._0476_ ;
 wire \INST_config_UART._0477_ ;
 wire \INST_config_UART._0478_ ;
 wire \INST_config_UART._0479_ ;
 wire \INST_config_UART._0480_ ;
 wire \INST_config_UART._0481_ ;
 wire \INST_config_UART._0482_ ;
 wire \INST_config_UART._0483_ ;
 wire \INST_config_UART._0484_ ;
 wire \INST_config_UART._0485_ ;
 wire \INST_config_UART._0486_ ;
 wire \INST_config_UART._0487_ ;
 wire \INST_config_UART._0488_ ;
 wire \INST_config_UART._0489_ ;
 wire \INST_config_UART._0490_ ;
 wire \INST_config_UART._0491_ ;
 wire \INST_config_UART._0492_ ;
 wire \INST_config_UART._0493_ ;
 wire \INST_config_UART._0494_ ;
 wire \INST_config_UART._0495_ ;
 wire \INST_config_UART._0496_ ;
 wire \INST_config_UART._0497_ ;
 wire \INST_config_UART._0498_ ;
 wire \INST_config_UART._0499_ ;
 wire \INST_config_UART._0500_ ;
 wire \INST_config_UART._0501_ ;
 wire \INST_config_UART._0502_ ;
 wire \INST_config_UART._0503_ ;
 wire \INST_config_UART._0504_ ;
 wire \INST_config_UART._0505_ ;
 wire \INST_config_UART._0506_ ;
 wire \INST_config_UART._0507_ ;
 wire \INST_config_UART._0508_ ;
 wire \INST_config_UART._0509_ ;
 wire \INST_config_UART._0510_ ;
 wire \INST_config_UART._0511_ ;
 wire \INST_config_UART._0512_ ;
 wire \INST_config_UART._0513_ ;
 wire \INST_config_UART._0514_ ;
 wire \INST_config_UART._0515_ ;
 wire \INST_config_UART._0516_ ;
 wire \INST_config_UART._0517_ ;
 wire \INST_config_UART._0518_ ;
 wire \INST_config_UART._0519_ ;
 wire \INST_config_UART._0520_ ;
 wire \INST_config_UART._0521_ ;
 wire \INST_config_UART._0522_ ;
 wire \INST_config_UART._0523_ ;
 wire \INST_config_UART._0524_ ;
 wire \INST_config_UART._0525_ ;
 wire \INST_config_UART._0526_ ;
 wire \INST_config_UART._0527_ ;
 wire \INST_config_UART._0528_ ;
 wire \INST_config_UART._0529_ ;
 wire \INST_config_UART._0530_ ;
 wire \INST_config_UART._0531_ ;
 wire \INST_config_UART._0532_ ;
 wire \INST_config_UART._0533_ ;
 wire \INST_config_UART._0534_ ;
 wire \INST_config_UART._0535_ ;
 wire \INST_config_UART._0536_ ;
 wire \INST_config_UART._0537_ ;
 wire \INST_config_UART._0538_ ;
 wire \INST_config_UART._0539_ ;
 wire \INST_config_UART._0540_ ;
 wire \INST_config_UART._0541_ ;
 wire \INST_config_UART._0542_ ;
 wire \INST_config_UART._0543_ ;
 wire \INST_config_UART._0544_ ;
 wire \INST_config_UART._0545_ ;
 wire \INST_config_UART._0546_ ;
 wire \INST_config_UART._0547_ ;
 wire \INST_config_UART._0548_ ;
 wire \INST_config_UART._0549_ ;
 wire \INST_config_UART._0550_ ;
 wire \INST_config_UART._0551_ ;
 wire \INST_config_UART._0552_ ;
 wire \INST_config_UART._0553_ ;
 wire \INST_config_UART._0554_ ;
 wire \INST_config_UART._0555_ ;
 wire \INST_config_UART._0556_ ;
 wire \INST_config_UART._0557_ ;
 wire \INST_config_UART._0558_ ;
 wire \INST_config_UART._0559_ ;
 wire \INST_config_UART._0560_ ;
 wire \INST_config_UART._0561_ ;
 wire \INST_config_UART._0562_ ;
 wire \INST_config_UART._0563_ ;
 wire \INST_config_UART._0564_ ;
 wire \INST_config_UART._0565_ ;
 wire \INST_config_UART._0566_ ;
 wire \INST_config_UART._0567_ ;
 wire \INST_config_UART._0568_ ;
 wire \INST_config_UART._0569_ ;
 wire \INST_config_UART._0570_ ;
 wire \INST_config_UART._0571_ ;
 wire \INST_config_UART._0572_ ;
 wire \INST_config_UART._0573_ ;
 wire \INST_config_UART._0574_ ;
 wire \INST_config_UART._0575_ ;
 wire \INST_config_UART._0576_ ;
 wire \INST_config_UART._0577_ ;
 wire \INST_config_UART._0578_ ;
 wire \INST_config_UART._0579_ ;
 wire \INST_config_UART._0580_ ;
 wire \INST_config_UART._0581_ ;
 wire \INST_config_UART._0582_ ;
 wire \INST_config_UART._0583_ ;
 wire \INST_config_UART._0584_ ;
 wire \INST_config_UART._0585_ ;
 wire \INST_config_UART._0586_ ;
 wire \INST_config_UART._0587_ ;
 wire \INST_config_UART._0588_ ;
 wire \INST_config_UART.blink[0] ;
 wire \INST_config_UART.blink[10] ;
 wire \INST_config_UART.blink[11] ;
 wire \INST_config_UART.blink[12] ;
 wire \INST_config_UART.blink[13] ;
 wire \INST_config_UART.blink[14] ;
 wire \INST_config_UART.blink[15] ;
 wire \INST_config_UART.blink[16] ;
 wire \INST_config_UART.blink[17] ;
 wire \INST_config_UART.blink[18] ;
 wire \INST_config_UART.blink[19] ;
 wire \INST_config_UART.blink[1] ;
 wire \INST_config_UART.blink[20] ;
 wire \INST_config_UART.blink[21] ;
 wire \INST_config_UART.blink[22] ;
 wire \INST_config_UART.blink[2] ;
 wire \INST_config_UART.blink[3] ;
 wire \INST_config_UART.blink[4] ;
 wire \INST_config_UART.blink[5] ;
 wire \INST_config_UART.blink[6] ;
 wire \INST_config_UART.blink[7] ;
 wire \INST_config_UART.blink[8] ;
 wire \INST_config_UART.blink[9] ;
 wire \Inst_bitbang._000_ ;
 wire \Inst_bitbang._001_ ;
 wire \Inst_bitbang._002_ ;
 wire \Inst_bitbang._003_ ;
 wire \Inst_bitbang._004_ ;
 wire \Inst_bitbang._005_ ;
 wire \Inst_bitbang._006_ ;
 wire \Inst_bitbang._007_ ;
 wire \Inst_bitbang._008_ ;
 wire \Inst_bitbang._009_ ;
 wire \Inst_bitbang._010_ ;
 wire \Inst_bitbang._011_ ;
 wire \Inst_bitbang._012_ ;
 wire \Inst_bitbang._013_ ;
 wire \Inst_bitbang._014_ ;
 wire \Inst_bitbang._015_ ;
 wire \Inst_bitbang._016_ ;
 wire \Inst_bitbang._017_ ;
 wire \Inst_bitbang._018_ ;
 wire \Inst_bitbang._019_ ;
 wire \Inst_bitbang._020_ ;
 wire \Inst_bitbang._021_ ;
 wire \Inst_bitbang._022_ ;
 wire \Inst_bitbang._023_ ;
 wire \Inst_bitbang._024_ ;
 wire \Inst_bitbang._025_ ;
 wire \Inst_bitbang._026_ ;
 wire \Inst_bitbang._027_ ;
 wire \Inst_bitbang._028_ ;
 wire \Inst_bitbang._029_ ;
 wire \Inst_bitbang._030_ ;
 wire \Inst_bitbang._031_ ;
 wire \Inst_bitbang._032_ ;
 wire \Inst_bitbang._033_ ;
 wire \Inst_bitbang._034_ ;
 wire \Inst_bitbang._035_ ;
 wire \Inst_bitbang._036_ ;
 wire \Inst_bitbang._037_ ;
 wire \Inst_bitbang._038_ ;
 wire \Inst_bitbang._039_ ;
 wire \Inst_bitbang._040_ ;
 wire \Inst_bitbang._041_ ;
 wire \Inst_bitbang._042_ ;
 wire \Inst_bitbang._043_ ;
 wire \Inst_bitbang._044_ ;
 wire \Inst_bitbang._045_ ;
 wire \Inst_bitbang._046_ ;
 wire \Inst_bitbang._047_ ;
 wire \Inst_bitbang._048_ ;
 wire \Inst_bitbang._049_ ;
 wire \Inst_bitbang._050_ ;
 wire \Inst_bitbang._051_ ;
 wire \Inst_bitbang._052_ ;
 wire \Inst_bitbang._053_ ;
 wire \Inst_bitbang._054_ ;
 wire \Inst_bitbang._055_ ;
 wire \Inst_bitbang._056_ ;
 wire \Inst_bitbang._057_ ;
 wire \Inst_bitbang._058_ ;
 wire \Inst_bitbang._059_ ;
 wire \Inst_bitbang._060_ ;
 wire \Inst_bitbang._061_ ;
 wire \Inst_bitbang._062_ ;
 wire \Inst_bitbang._063_ ;
 wire \Inst_bitbang._064_ ;
 wire \Inst_bitbang._065_ ;
 wire \Inst_bitbang._066_ ;
 wire \Inst_bitbang._067_ ;
 wire \Inst_bitbang._068_ ;
 wire \Inst_bitbang._069_ ;
 wire \Inst_bitbang._070_ ;
 wire \Inst_bitbang._071_ ;
 wire \Inst_bitbang._072_ ;
 wire \Inst_bitbang._073_ ;
 wire \Inst_bitbang._074_ ;
 wire \Inst_bitbang._075_ ;
 wire \Inst_bitbang._076_ ;
 wire \Inst_bitbang._077_ ;
 wire \Inst_bitbang._078_ ;
 wire \Inst_bitbang._079_ ;
 wire \Inst_bitbang._080_ ;
 wire \Inst_bitbang._081_ ;
 wire \Inst_bitbang._082_ ;
 wire \Inst_bitbang._083_ ;
 wire \Inst_bitbang._084_ ;
 wire \Inst_bitbang._085_ ;
 wire \Inst_bitbang._086_ ;
 wire \Inst_bitbang._087_ ;
 wire \Inst_bitbang._088_ ;
 wire \Inst_bitbang._089_ ;
 wire \Inst_bitbang._090_ ;
 wire \Inst_bitbang._091_ ;
 wire \Inst_bitbang._092_ ;
 wire \Inst_bitbang._093_ ;
 wire \Inst_bitbang._094_ ;
 wire \Inst_bitbang._095_ ;
 wire \Inst_bitbang._096_ ;
 wire \Inst_bitbang._097_ ;
 wire \Inst_bitbang._098_ ;
 wire \Inst_bitbang._099_ ;
 wire \Inst_bitbang._100_ ;
 wire \Inst_bitbang._101_ ;
 wire \Inst_bitbang._102_ ;
 wire \Inst_bitbang._103_ ;
 wire \Inst_bitbang._104_ ;
 wire \Inst_bitbang._105_ ;
 wire \Inst_bitbang._106_ ;
 wire \Inst_bitbang._107_ ;
 wire \Inst_bitbang._108_ ;
 wire \Inst_bitbang._109_ ;
 wire \Inst_bitbang._110_ ;
 wire \Inst_bitbang._111_ ;
 wire \Inst_bitbang._112_ ;
 wire \Inst_bitbang._113_ ;
 wire \Inst_bitbang._114_ ;
 wire \Inst_bitbang._115_ ;
 wire \Inst_bitbang._116_ ;
 wire \Inst_bitbang._117_ ;
 wire \Inst_bitbang._118_ ;
 wire \Inst_bitbang._119_ ;
 wire \Inst_bitbang._120_ ;
 wire \Inst_bitbang._121_ ;
 wire \Inst_bitbang._122_ ;
 wire \Inst_bitbang._123_ ;
 wire \Inst_bitbang._124_ ;
 wire \Inst_bitbang._125_ ;
 wire \Inst_bitbang._126_ ;
 wire \Inst_bitbang._127_ ;
 wire \Inst_bitbang._128_ ;
 wire \Inst_bitbang._129_ ;
 wire \Inst_bitbang._130_ ;
 wire \Inst_bitbang._131_ ;
 wire \Inst_bitbang._132_ ;
 wire \Inst_bitbang._133_ ;
 wire \Inst_bitbang._134_ ;
 wire \Inst_bitbang._135_ ;
 wire \Inst_bitbang._136_ ;
 wire \Inst_bitbang._137_ ;
 wire \Inst_bitbang._138_ ;
 wire \Inst_bitbang._139_ ;
 wire \Inst_bitbang._140_ ;
 wire \Inst_bitbang._141_ ;
 wire \Inst_bitbang._142_ ;
 wire \Inst_bitbang._143_ ;
 wire \Inst_bitbang._144_ ;
 wire \Inst_bitbang._145_ ;
 wire \Inst_bitbang._146_ ;
 wire \Inst_bitbang._147_ ;
 wire \Inst_bitbang._148_ ;
 wire \Inst_bitbang._149_ ;
 wire \Inst_bitbang._150_ ;
 wire \Inst_bitbang._151_ ;
 wire \Inst_bitbang._152_ ;
 wire \Inst_bitbang._153_ ;
 wire \Inst_bitbang._154_ ;
 wire \Inst_bitbang._155_ ;
 wire \Inst_bitbang._156_ ;
 wire \Inst_bitbang._157_ ;
 wire \Inst_bitbang._158_ ;
 wire \Inst_bitbang._159_ ;
 wire \Inst_bitbang._160_ ;
 wire \Inst_bitbang._161_ ;
 wire \Inst_bitbang._162_ ;
 wire \Inst_bitbang._163_ ;
 wire \Inst_bitbang._164_ ;
 wire \Inst_bitbang._165_ ;
 wire \Inst_bitbang._166_ ;
 wire \Inst_bitbang._167_ ;
 wire \Inst_bitbang._168_ ;
 wire \Inst_bitbang._169_ ;
 wire \Inst_bitbang._170_ ;
 wire \Inst_bitbang._171_ ;
 wire \Inst_bitbang._172_ ;
 wire \Inst_bitbang._173_ ;
 wire \Inst_bitbang._174_ ;
 wire \Inst_bitbang._175_ ;
 wire \Inst_bitbang._176_ ;
 wire \Inst_bitbang._177_ ;
 wire \Inst_bitbang._178_ ;
 wire \Inst_bitbang._179_ ;
 wire \Inst_bitbang._180_ ;
 wire \Inst_bitbang.active ;
 wire \Inst_bitbang.data[0] ;
 wire \Inst_bitbang.data[10] ;
 wire \Inst_bitbang.data[11] ;
 wire \Inst_bitbang.data[12] ;
 wire \Inst_bitbang.data[13] ;
 wire \Inst_bitbang.data[14] ;
 wire \Inst_bitbang.data[15] ;
 wire \Inst_bitbang.data[16] ;
 wire \Inst_bitbang.data[17] ;
 wire \Inst_bitbang.data[18] ;
 wire \Inst_bitbang.data[19] ;
 wire \Inst_bitbang.data[1] ;
 wire \Inst_bitbang.data[20] ;
 wire \Inst_bitbang.data[21] ;
 wire \Inst_bitbang.data[22] ;
 wire \Inst_bitbang.data[23] ;
 wire \Inst_bitbang.data[24] ;
 wire \Inst_bitbang.data[25] ;
 wire \Inst_bitbang.data[26] ;
 wire \Inst_bitbang.data[27] ;
 wire \Inst_bitbang.data[28] ;
 wire \Inst_bitbang.data[29] ;
 wire \Inst_bitbang.data[2] ;
 wire \Inst_bitbang.data[30] ;
 wire \Inst_bitbang.data[31] ;
 wire \Inst_bitbang.data[3] ;
 wire \Inst_bitbang.data[4] ;
 wire \Inst_bitbang.data[5] ;
 wire \Inst_bitbang.data[6] ;
 wire \Inst_bitbang.data[7] ;
 wire \Inst_bitbang.data[8] ;
 wire \Inst_bitbang.data[9] ;
 wire \Inst_bitbang.local_strobe ;
 wire \Inst_bitbang.old_local_strobe ;
 wire \Inst_bitbang.s_clk_sample[0] ;
 wire \Inst_bitbang.s_clk_sample[1] ;
 wire \Inst_bitbang.s_clk_sample[2] ;
 wire \Inst_bitbang.s_clk_sample[3] ;
 wire \Inst_bitbang.s_data_sample[0] ;
 wire \Inst_bitbang.s_data_sample[1] ;
 wire \Inst_bitbang.s_data_sample[2] ;
 wire \Inst_bitbang.s_data_sample[3] ;
 wire \Inst_bitbang.serial_control[0] ;
 wire \Inst_bitbang.serial_control[10] ;
 wire \Inst_bitbang.serial_control[11] ;
 wire \Inst_bitbang.serial_control[12] ;
 wire \Inst_bitbang.serial_control[13] ;
 wire \Inst_bitbang.serial_control[14] ;
 wire \Inst_bitbang.serial_control[15] ;
 wire \Inst_bitbang.serial_control[1] ;
 wire \Inst_bitbang.serial_control[2] ;
 wire \Inst_bitbang.serial_control[3] ;
 wire \Inst_bitbang.serial_control[4] ;
 wire \Inst_bitbang.serial_control[5] ;
 wire \Inst_bitbang.serial_control[6] ;
 wire \Inst_bitbang.serial_control[7] ;
 wire \Inst_bitbang.serial_control[8] ;
 wire \Inst_bitbang.serial_control[9] ;
 wire \Inst_bitbang.serial_data[0] ;
 wire \Inst_bitbang.serial_data[10] ;
 wire \Inst_bitbang.serial_data[11] ;
 wire \Inst_bitbang.serial_data[12] ;
 wire \Inst_bitbang.serial_data[13] ;
 wire \Inst_bitbang.serial_data[14] ;
 wire \Inst_bitbang.serial_data[15] ;
 wire \Inst_bitbang.serial_data[16] ;
 wire \Inst_bitbang.serial_data[17] ;
 wire \Inst_bitbang.serial_data[18] ;
 wire \Inst_bitbang.serial_data[19] ;
 wire \Inst_bitbang.serial_data[1] ;
 wire \Inst_bitbang.serial_data[20] ;
 wire \Inst_bitbang.serial_data[21] ;
 wire \Inst_bitbang.serial_data[22] ;
 wire \Inst_bitbang.serial_data[23] ;
 wire \Inst_bitbang.serial_data[24] ;
 wire \Inst_bitbang.serial_data[25] ;
 wire \Inst_bitbang.serial_data[26] ;
 wire \Inst_bitbang.serial_data[27] ;
 wire \Inst_bitbang.serial_data[28] ;
 wire \Inst_bitbang.serial_data[29] ;
 wire \Inst_bitbang.serial_data[2] ;
 wire \Inst_bitbang.serial_data[30] ;
 wire \Inst_bitbang.serial_data[31] ;
 wire \Inst_bitbang.serial_data[3] ;
 wire \Inst_bitbang.serial_data[4] ;
 wire \Inst_bitbang.serial_data[5] ;
 wire \Inst_bitbang.serial_data[6] ;
 wire \Inst_bitbang.serial_data[7] ;
 wire \Inst_bitbang.serial_data[8] ;
 wire \Inst_bitbang.serial_data[9] ;
 wire \Inst_bitbang.strobe ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\ConfigFSM_inst.WriteData[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\ConfigFSM_inst.WriteData[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._121__A  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._121__C  (.DIODE(\ConfigFSM_inst.WriteData[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._122__A  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._124__A  (.DIODE(\ConfigFSM_inst.WriteData[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._124__B  (.DIODE(\ConfigFSM_inst.WriteData[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._124__C_N  (.DIODE(\ConfigFSM_inst.WriteData[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._124__D_N  (.DIODE(\ConfigFSM_inst.WriteData[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._125__A  (.DIODE(\ConfigFSM_inst.WriteData[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._125__B  (.DIODE(\ConfigFSM_inst.WriteData[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._125__C  (.DIODE(\ConfigFSM_inst.WriteData[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._125__D_N  (.DIODE(\ConfigFSM_inst.WriteData[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._126__A  (.DIODE(\ConfigFSM_inst.WriteData[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._126__B  (.DIODE(\ConfigFSM_inst.WriteData[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._126__D_N  (.DIODE(\ConfigFSM_inst.WriteData[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._127__B  (.DIODE(\ConfigFSM_inst.WriteData[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._127__C  (.DIODE(\ConfigFSM_inst.WriteData[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._127__D  (.DIODE(\ConfigFSM_inst.WriteData[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._129__A  (.DIODE(\ConfigFSM_inst.WriteData[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._129__B  (.DIODE(\ConfigFSM_inst.WriteData[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._129__C_N  (.DIODE(\ConfigFSM_inst.WriteData[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._129__D_N  (.DIODE(\ConfigFSM_inst.WriteData[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._130__A  (.DIODE(\ConfigFSM_inst.WriteData[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._130__B  (.DIODE(\ConfigFSM_inst.WriteData[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._130__C_N  (.DIODE(\ConfigFSM_inst.WriteData[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._130__D_N  (.DIODE(\ConfigFSM_inst.WriteData[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._131__A  (.DIODE(\ConfigFSM_inst.WriteData[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._131__B  (.DIODE(\ConfigFSM_inst.WriteData[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._131__C_N  (.DIODE(\ConfigFSM_inst.WriteData[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._131__D_N  (.DIODE(\ConfigFSM_inst.WriteData[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._132__A  (.DIODE(\ConfigFSM_inst.WriteData[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._132__B  (.DIODE(\ConfigFSM_inst.WriteData[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._132__C  (.DIODE(\ConfigFSM_inst.WriteData[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._132__D  (.DIODE(\ConfigFSM_inst.WriteData[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._141__A  (.DIODE(\ConfigFSM_inst.WriteData[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._143__B1  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._181__A0  (.DIODE(\ConfigFSM_inst.WriteData[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._181__S  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._183__A0  (.DIODE(\ConfigFSM_inst.WriteData[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._183__S  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._185__A0  (.DIODE(\ConfigFSM_inst.WriteData[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._185__S  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._187__A0  (.DIODE(\ConfigFSM_inst.WriteData[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._187__S  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._189__A0  (.DIODE(\ConfigFSM_inst.WriteData[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._189__S  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._191__A0  (.DIODE(\ConfigFSM_inst.WriteData[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._191__S  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._193__A0  (.DIODE(\ConfigFSM_inst.WriteData[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._193__S  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._195__A0  (.DIODE(\ConfigFSM_inst.WriteData[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._195__S  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._197__A0  (.DIODE(\ConfigFSM_inst.WriteData[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._197__S  (.DIODE(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._200__A0  (.DIODE(\ConfigFSM_inst.WriteData[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._202__A0  (.DIODE(\ConfigFSM_inst.WriteData[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._204__A0  (.DIODE(\ConfigFSM_inst.WriteData[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._206__A0  (.DIODE(\ConfigFSM_inst.WriteData[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._208__A0  (.DIODE(\ConfigFSM_inst.WriteData[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._210__A0  (.DIODE(\ConfigFSM_inst.WriteData[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._212__A0  (.DIODE(\ConfigFSM_inst.WriteData[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._214__A0  (.DIODE(\ConfigFSM_inst.WriteData[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._216__A0  (.DIODE(\ConfigFSM_inst.WriteData[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._218__A0  (.DIODE(\ConfigFSM_inst.WriteData[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._221__A0  (.DIODE(\ConfigFSM_inst.WriteData[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._223__A0  (.DIODE(\ConfigFSM_inst.WriteData[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._225__A0  (.DIODE(\ConfigFSM_inst.WriteData[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._227__A0  (.DIODE(\ConfigFSM_inst.WriteData[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._229__A0  (.DIODE(\ConfigFSM_inst.WriteData[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._231__A0  (.DIODE(\ConfigFSM_inst.WriteData[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._233__A0  (.DIODE(\ConfigFSM_inst.WriteData[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._237__A0  (.DIODE(\ConfigFSM_inst.WriteData[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._241__A0  (.DIODE(\ConfigFSM_inst.WriteData[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._243__A0  (.DIODE(\ConfigFSM_inst.WriteData[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._245__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._245__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._246__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._246__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._247__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._247__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._248__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._248__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._249__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._249__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._250__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._250__SET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._251__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._251__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._252__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._252__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._253__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._253__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._254__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._254__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._255__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._255__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._256__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._256__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._257__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._257__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._258__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._258__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._259__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._259__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._260__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._260__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._261__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._261__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._262__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._262__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._263__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._263__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._264__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._264__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._265__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._265__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._266__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._266__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._267__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._267__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._268__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._268__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._269__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._269__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._270__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._270__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._271__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._271__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._272__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._272__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._273__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._273__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._274__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._274__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._275__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._275__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._276__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._276__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._277__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._277__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._278__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._278__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._279__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._279__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._280__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._280__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._281__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._281__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._282__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._282__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._283__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._283__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._284__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._284__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._285__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._285__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._286__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._286__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._287__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_ConfigFSM_inst._287__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0597__A_N  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0612__A  (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0623__B  (.DIODE(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0623__C_N  (.DIODE(\INST_config_UART.ReceivedWord[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0623__D_N  (.DIODE(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0624__A  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0629__A  (.DIODE(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0629__C_N  (.DIODE(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0632__B  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0633__B_N  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0636__A1  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0636__A2  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0655__B1  (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0656__A  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0662__A  (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0759__A1  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0763__A0  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0763__A1  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0829__A1  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0829__B2  (.DIODE(\INST_config_UART.ReceivedWord[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0833__A1  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0840__A1  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0842__A1  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0844__A1  (.DIODE(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0846__A1  (.DIODE(\INST_config_UART.ReceivedWord[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0848__A1  (.DIODE(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0855__A1  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0855__B2  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0859__A1  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0859__B2  (.DIODE(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0863__A1  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0870__A1  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0872__A1  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0874__A1  (.DIODE(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0876__A1  (.DIODE(\INST_config_UART.ReceivedWord[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0878__A1  (.DIODE(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0892__B1  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0911__S  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0976__A  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0978__A1  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0978__B2  (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._0999__B1  (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1013__A0  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1018__A0  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1027__A0  (.DIODE(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1034__A0  (.DIODE(\INST_config_UART.ReceivedWord[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1040__A0  (.DIODE(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1107__A1  (.DIODE(\INST_config_UART.RxLocal ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1107__B2  (.DIODE(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1114__A1  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1116__A1  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1118__A1  (.DIODE(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1120__A1  (.DIODE(\INST_config_UART.ReceivedWord[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1122__A1  (.DIODE(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1132__A1  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1134__A1  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1136__A1  (.DIODE(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1138__A1  (.DIODE(\INST_config_UART.ReceivedWord[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1140__A1  (.DIODE(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1144__A  (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1144__B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1150__A1  (.DIODE(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1152__A1  (.DIODE(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1154__A1  (.DIODE(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1156__A1  (.DIODE(\INST_config_UART.ReceivedWord[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1158__A1  (.DIODE(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1178__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1178__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1179__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1179__SET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1180__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1180__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1181__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1181__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1182__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1182__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1183__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1183__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1184__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1184__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1185__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1185__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1186__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1186__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1187__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1187__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1188__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1188__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1189__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1189__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1190__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1190__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1191__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1191__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1192__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1192__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1193__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1193__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1194__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1194__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1195__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1195__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1196__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1196__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1197__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1197__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1198__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1198__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1199__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1199__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1200__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1200__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1201__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1201__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1202__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1202__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1203__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1203__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1204__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1204__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1205__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1205__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1206__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1206__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1207__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1207__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1208__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1208__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1209__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1209__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1210__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1210__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1211__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1211__SET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1212__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1212__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1213__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1213__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1214__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1214__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1215__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1215__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1216__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1216__SET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1217__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1217__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1218__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1218__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1219__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1219__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1220__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1220__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1221__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1221__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1222__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1222__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1223__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1223__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1224__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1224__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1225__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1225__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1226__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1226__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1227__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1227__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1228__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1228__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1229__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1229__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1230__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1230__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1231__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1231__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1232__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1232__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1233__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1233__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1234__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1234__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1235__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1235__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1236__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1236__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1237__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1237__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1238__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1238__SET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1239__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1239__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1240__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1240__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1241__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1241__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1242__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1242__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1243__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1243__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1244__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1245__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1245__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1246__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1246__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1247__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1247__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1248__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1248__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1249__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1249__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1250__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1250__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1251__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1251__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1252__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1252__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1253__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1253__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1254__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1254__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1255__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1255__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1256__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1256__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1257__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1257__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1258__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1258__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1259__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1259__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1260__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1260__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1261__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1261__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1262__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1262__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1263__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1263__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1264__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1264__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1265__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1265__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1266__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1266__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1267__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1267__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1268__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1268__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1269__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1269__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1270__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1270__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1271__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1272__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1272__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1273__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1273__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1274__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1274__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1275__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1275__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1276__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1276__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1277__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1277__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1278__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1278__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1279__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1279__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1280__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1280__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1281__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1281__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1282__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1282__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1283__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1283__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1284__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1284__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1285__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1285__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1286__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1286__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1287__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1287__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1288__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1288__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1289__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1289__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1290__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1290__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1291__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1291__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1292__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1292__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1293__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1293__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1294__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1294__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1295__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1295__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1296__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1296__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1297__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1297__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1298__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1298__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1299__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1299__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1300__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1300__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1301__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1301__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1302__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1302__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1303__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1303__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1304__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1304__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1305__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1305__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1306__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1306__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1307__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1307__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1308__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1308__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1309__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1309__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1310__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1310__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1311__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1311__SET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1312__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1312__SET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1313__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1313__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1314__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1314__SET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1315__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1315__SET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1316__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1316__SET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1317__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1317__SET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1318__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1318__SET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1319__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1319__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1320__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1320__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1321__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1321__SET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1322__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1322__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1323__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1323__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1324__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1324__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1325__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1325__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1326__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1326__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1327__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1327__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1328__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1328__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1329__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1329__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1330__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1330__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1331__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1331__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1332__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1332__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1333__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1333__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1334__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1334__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1335__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1335__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1336__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1336__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1337__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1337__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1338__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1338__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1339__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1339__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1340__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1340__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1341__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1341__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1342__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1342__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1343__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1343__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1344__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1344__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1345__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1345__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1346__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1346__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1347__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1347__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1348__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1348__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1349__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1349__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1350__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1350__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1351__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1351__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1352__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1352__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1353__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1353__SET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1354__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1355__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1356__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1357__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1358__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1359__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1360__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1361__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1362__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1362__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1363__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1363__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1364__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1364__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1365__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1365__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1366__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1366__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1367__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1367__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1368__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1368__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1369__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1369__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1370__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_INST_config_UART._1370__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._186__A  (.DIODE(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._187__A  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._191__A  (.DIODE(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._193__A  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._194__S  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._196__S  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._198__S  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._200__S  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._202__S  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._204__S  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._206__S  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._208__S  (.DIODE(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._210__A  (.DIODE(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._231__A  (.DIODE(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._252__S  (.DIODE(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._254__S  (.DIODE(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._256__S  (.DIODE(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._258__S  (.DIODE(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._261__A  (.DIODE(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._282__A  (.DIODE(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._303__A  (.DIODE(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._324__S  (.DIODE(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._326__S  (.DIODE(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._362__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._362__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._363__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._363__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._364__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._364__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._365__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._365__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._366__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._366__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._367__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._367__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._368__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._368__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._369__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._369__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._370__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._370__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._371__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._371__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._372__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._372__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._373__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._373__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._374__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._374__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._375__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._375__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._376__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._376__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._377__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._377__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._378__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._378__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._379__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._379__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._380__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._380__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._381__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._381__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._382__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._382__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._383__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._383__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._384__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._384__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._385__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._385__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._386__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._386__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._387__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._387__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._388__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._388__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._389__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._389__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._390__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._390__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._391__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._391__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._392__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._392__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._393__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._393__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._394__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._394__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._395__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._395__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._396__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._396__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._397__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._397__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._398__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._398__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._399__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._399__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._400__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._400__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._401__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._401__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._402__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._402__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._403__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._403__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._404__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._404__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._405__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._405__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._406__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._406__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._407__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._407__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._408__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._408__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._409__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._409__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._410__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._410__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._411__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._411__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._412__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._412__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._413__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._413__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._414__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._414__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._415__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._415__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._416__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._416__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._417__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._417__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._418__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._418__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._419__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._419__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._420__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._420__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._421__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._421__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._422__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._422__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._423__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._423__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._424__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._424__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._425__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._425__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._426__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._426__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._427__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._427__RESET_B  (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._428__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._428__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._429__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._429__RESET_B  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._430__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._430__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._431__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._431__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._432__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._432__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._433__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._433__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._434__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._434__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._435__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._435__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._436__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._436__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._437__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._437__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._438__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._438__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._439__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._439__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._440__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._440__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._441__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._441__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._442__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._442__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._443__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._443__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._444__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._444__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._445__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._445__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._446__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._446__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._447__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._447__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._448__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._448__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._449__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._449__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._450__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._450__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._451__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._451__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._452__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._452__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._453__CLK  (.DIODE(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_bitbang._453__RESET_B  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__A (.DIODE(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__A (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__104__A (.DIODE(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__105__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__106__A (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__109__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__112__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__115__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__118__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__S (.DIODE(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__A (.DIODE(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__A (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__168__S (.DIODE(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__169__S (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__171__S (.DIODE(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__172__S (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__S (.DIODE(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__175__S (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__177__S (.DIODE(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__178__S (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(\ConfigFSM_inst.WriteData[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__182__A (.DIODE(\ConfigFSM_inst.WriteData[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__183__A (.DIODE(\ConfigFSM_inst.WriteData[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__A (.DIODE(\ConfigFSM_inst.WriteData[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__185__A (.DIODE(\ConfigFSM_inst.WriteData[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__186__A (.DIODE(\ConfigFSM_inst.WriteData[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__187__A (.DIODE(\ConfigFSM_inst.WriteData[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__A (.DIODE(\ConfigFSM_inst.WriteData[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__A (.DIODE(\ConfigFSM_inst.WriteData[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__190__A (.DIODE(\ConfigFSM_inst.WriteData[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__A (.DIODE(\ConfigFSM_inst.WriteData[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A (.DIODE(\ConfigFSM_inst.WriteData[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A (.DIODE(\ConfigFSM_inst.WriteData[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__194__A (.DIODE(\ConfigFSM_inst.WriteData[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__A (.DIODE(\ConfigFSM_inst.WriteData[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__196__A (.DIODE(\ConfigFSM_inst.WriteData[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A (.DIODE(\ConfigFSM_inst.WriteData[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__198__A (.DIODE(\ConfigFSM_inst.WriteData[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__199__A (.DIODE(\ConfigFSM_inst.WriteData[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__200__A (.DIODE(\ConfigFSM_inst.WriteData[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__201__A (.DIODE(\ConfigFSM_inst.WriteData[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__202__A (.DIODE(\ConfigFSM_inst.WriteData[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__203__A (.DIODE(\ConfigFSM_inst.WriteData[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__204__A (.DIODE(\ConfigFSM_inst.WriteData[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__205__A (.DIODE(\ConfigFSM_inst.WriteData[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__206__A (.DIODE(\ConfigFSM_inst.WriteData[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__207__A (.DIODE(\ConfigFSM_inst.WriteData[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__209__A (.DIODE(\ConfigFSM_inst.WriteData[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__A (.DIODE(\ConfigFSM_inst.WriteData[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA__212__A (.DIODE(\ConfigFSM_inst.WriteData[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew111_A (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_load_slew112_A (.DIODE(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2b_1 \ConfigFSM_inst._120_  (.A_N(\ConfigFSM_inst.old_reset ),
    .B(\ConfigFSM_inst.FSM_Reset ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._041_ ));
 sky130_fd_sc_hd__and3_1 \ConfigFSM_inst._121_  (.A(net72),
    .B(\ConfigFSM_inst.state[2] ),
    .C(\ConfigFSM_inst.WriteData[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._042_ ));
 sky130_fd_sc_hd__clkbuf_2 \ConfigFSM_inst._122_  (.A(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._043_ ));
 sky130_fd_sc_hd__nor2_1 \ConfigFSM_inst._123_  (.A(\ConfigFSM_inst._043_ ),
    .B(\ConfigFSM_inst._041_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._044_ ));
 sky130_fd_sc_hd__or4bb_1 \ConfigFSM_inst._124_  (.A(\ConfigFSM_inst.WriteData[18] ),
    .B(\ConfigFSM_inst.WriteData[22] ),
    .C_N(\ConfigFSM_inst.WriteData[23] ),
    .D_N(\ConfigFSM_inst.WriteData[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._045_ ));
 sky130_fd_sc_hd__or4b_1 \ConfigFSM_inst._125_  (.A(\ConfigFSM_inst.WriteData[17] ),
    .B(\ConfigFSM_inst.WriteData[16] ),
    .C(\ConfigFSM_inst.WriteData[19] ),
    .D_N(\ConfigFSM_inst.WriteData[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._046_ ));
 sky130_fd_sc_hd__or4bb_1 \ConfigFSM_inst._126_  (.A(\ConfigFSM_inst.WriteData[24] ),
    .B(\ConfigFSM_inst.WriteData[26] ),
    .C_N(\ConfigFSM_inst.WriteData[27] ),
    .D_N(\ConfigFSM_inst.WriteData[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._047_ ));
 sky130_fd_sc_hd__and4_1 \ConfigFSM_inst._127_  (.A(\ConfigFSM_inst.WriteData[29] ),
    .B(\ConfigFSM_inst.WriteData[28] ),
    .C(\ConfigFSM_inst.WriteData[31] ),
    .D(\ConfigFSM_inst.WriteData[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._048_ ));
 sky130_fd_sc_hd__or4b_1 \ConfigFSM_inst._128_  (.A(\ConfigFSM_inst._045_ ),
    .B(\ConfigFSM_inst._046_ ),
    .C(\ConfigFSM_inst._047_ ),
    .D_N(\ConfigFSM_inst._048_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._049_ ));
 sky130_fd_sc_hd__or4bb_1 \ConfigFSM_inst._129_  (.A(\ConfigFSM_inst.WriteData[2] ),
    .B(\ConfigFSM_inst.WriteData[6] ),
    .C_N(\ConfigFSM_inst.WriteData[5] ),
    .D_N(\ConfigFSM_inst.WriteData[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._050_ ));
 sky130_fd_sc_hd__or4bb_1 \ConfigFSM_inst._130_  (.A(\ConfigFSM_inst.WriteData[1] ),
    .B(\ConfigFSM_inst.WriteData[3] ),
    .C_N(\ConfigFSM_inst.WriteData[20] ),
    .D_N(\ConfigFSM_inst.WriteData[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._051_ ));
 sky130_fd_sc_hd__or4bb_1 \ConfigFSM_inst._131_  (.A(\ConfigFSM_inst.WriteData[8] ),
    .B(\ConfigFSM_inst.WriteData[10] ),
    .C_N(\ConfigFSM_inst.WriteData[9] ),
    .D_N(\ConfigFSM_inst.WriteData[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._052_ ));
 sky130_fd_sc_hd__and4_1 \ConfigFSM_inst._132_  (.A(\ConfigFSM_inst.WriteData[11] ),
    .B(\ConfigFSM_inst.WriteData[13] ),
    .C(\ConfigFSM_inst.WriteData[12] ),
    .D(\ConfigFSM_inst.WriteData[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._053_ ));
 sky130_fd_sc_hd__or4b_1 \ConfigFSM_inst._133_  (.A(\ConfigFSM_inst._050_ ),
    .B(\ConfigFSM_inst._051_ ),
    .C(\ConfigFSM_inst._052_ ),
    .D_N(\ConfigFSM_inst._053_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._054_ ));
 sky130_fd_sc_hd__o31a_1 \ConfigFSM_inst._134_  (.A1(\ConfigFSM_inst._044_ ),
    .A2(\ConfigFSM_inst._049_ ),
    .A3(\ConfigFSM_inst._054_ ),
    .B1(\ConfigFSM_inst.state[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._055_ ));
 sky130_fd_sc_hd__or3_1 \ConfigFSM_inst._135_  (.A(\ConfigFSM_inst._041_ ),
    .B(\ConfigFSM_inst._042_ ),
    .C(\ConfigFSM_inst._055_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._056_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._136_  (.A(\ConfigFSM_inst._056_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._002_ ));
 sky130_fd_sc_hd__nand2b_2 \ConfigFSM_inst._137_  (.A_N(\ConfigFSM_inst.old_reset ),
    .B(\ConfigFSM_inst.FSM_Reset ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._057_ ));
 sky130_fd_sc_hd__nand2_1 \ConfigFSM_inst._138_  (.A(\ConfigFSM_inst.state[1] ),
    .B(\ConfigFSM_inst._057_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._058_ ));
 sky130_fd_sc_hd__or3_1 \ConfigFSM_inst._139_  (.A(\ConfigFSM_inst.FrameShiftState[3] ),
    .B(\ConfigFSM_inst.FrameShiftState[2] ),
    .C(\ConfigFSM_inst.FrameShiftState[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._059_ ));
 sky130_fd_sc_hd__and4bb_1 \ConfigFSM_inst._140_  (.A_N(\ConfigFSM_inst.FrameShiftState[1] ),
    .B_N(\ConfigFSM_inst._059_ ),
    .C(\ConfigFSM_inst._043_ ),
    .D(\ConfigFSM_inst.FrameShiftState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._060_ ));
 sky130_fd_sc_hd__or4bb_4 \ConfigFSM_inst._141_  (.A(\ConfigFSM_inst.WriteData[20] ),
    .B(\ConfigFSM_inst._041_ ),
    .C_N(\ConfigFSM_inst._043_ ),
    .D_N(\ConfigFSM_inst.state[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._061_ ));
 sky130_fd_sc_hd__buf_4 \ConfigFSM_inst._142_  (.A(\ConfigFSM_inst._061_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._062_ ));
 sky130_fd_sc_hd__o21ai_1 \ConfigFSM_inst._143_  (.A1(\ConfigFSM_inst._058_ ),
    .A2(\ConfigFSM_inst._060_ ),
    .B1(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._003_ ));
 sky130_fd_sc_hd__nor2_1 \ConfigFSM_inst._144_  (.A(\ConfigFSM_inst._049_ ),
    .B(\ConfigFSM_inst._054_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._063_ ));
 sky130_fd_sc_hd__and3_1 \ConfigFSM_inst._145_  (.A(\ConfigFSM_inst._043_ ),
    .B(\ConfigFSM_inst.state[0] ),
    .C(\ConfigFSM_inst._057_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._064_ ));
 sky130_fd_sc_hd__a32o_1 \ConfigFSM_inst._146_  (.A1(\ConfigFSM_inst.state[1] ),
    .A2(\ConfigFSM_inst._057_ ),
    .A3(\ConfigFSM_inst._060_ ),
    .B1(\ConfigFSM_inst._044_ ),
    .B2(\ConfigFSM_inst.state[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._065_ ));
 sky130_fd_sc_hd__a21o_1 \ConfigFSM_inst._147_  (.A1(\ConfigFSM_inst._063_ ),
    .A2(\ConfigFSM_inst._064_ ),
    .B1(\ConfigFSM_inst._065_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._004_ ));
 sky130_fd_sc_hd__or2_1 \ConfigFSM_inst._148_  (.A(\ConfigFSM_inst.oldFrameStrobe ),
    .B(\ConfigFSM_inst.FrameStrobe ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._066_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._149_  (.A(\ConfigFSM_inst._066_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._001_ ));
 sky130_fd_sc_hd__or2b_1 \ConfigFSM_inst._150_  (.A(\ConfigFSM_inst.FrameShiftState[0] ),
    .B_N(\ConfigFSM_inst._043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._067_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._151_  (.A(\ConfigFSM_inst._067_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.RowSelect[0] ));
 sky130_fd_sc_hd__or2b_1 \ConfigFSM_inst._152_  (.A(\ConfigFSM_inst.FrameShiftState[1] ),
    .B_N(\ConfigFSM_inst._043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._068_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._153_  (.A(\ConfigFSM_inst._068_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.RowSelect[1] ));
 sky130_fd_sc_hd__or2b_1 \ConfigFSM_inst._154_  (.A(\ConfigFSM_inst.FrameShiftState[2] ),
    .B_N(\ConfigFSM_inst._043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._069_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._155_  (.A(\ConfigFSM_inst._069_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.RowSelect[2] ));
 sky130_fd_sc_hd__inv_2 \ConfigFSM_inst._156_  (.A(\ConfigFSM_inst.FrameShiftState[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._070_ ));
 sky130_fd_sc_hd__nand2_1 \ConfigFSM_inst._157_  (.A(\ConfigFSM_inst._043_ ),
    .B(\ConfigFSM_inst._070_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst.RowSelect[3] ));
 sky130_fd_sc_hd__or2b_1 \ConfigFSM_inst._158_  (.A(\ConfigFSM_inst.FrameShiftState[4] ),
    .B_N(\ConfigFSM_inst._043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._071_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._159_  (.A(\ConfigFSM_inst._071_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.RowSelect[4] ));
 sky130_fd_sc_hd__and3_1 \ConfigFSM_inst._160_  (.A(\ConfigFSM_inst.state[1] ),
    .B(\ConfigFSM_inst._057_ ),
    .C(\ConfigFSM_inst._060_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._072_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._161_  (.A(\ConfigFSM_inst._072_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._000_ ));
 sky130_fd_sc_hd__o21ai_1 \ConfigFSM_inst._162_  (.A1(\ConfigFSM_inst.state[2] ),
    .A2(\ConfigFSM_inst.state[1] ),
    .B1(\ConfigFSM_inst._043_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._073_ ));
 sky130_fd_sc_hd__or2_1 \ConfigFSM_inst._163_  (.A(\ConfigFSM_inst._042_ ),
    .B(\ConfigFSM_inst._073_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._074_ ));
 sky130_fd_sc_hd__nor2_1 \ConfigFSM_inst._164_  (.A(\ConfigFSM_inst._058_ ),
    .B(\ConfigFSM_inst._074_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._075_ ));
 sky130_fd_sc_hd__o21a_1 \ConfigFSM_inst._165_  (.A1(\ConfigFSM_inst._042_ ),
    .A2(\ConfigFSM_inst._073_ ),
    .B1(\ConfigFSM_inst._057_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._076_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._166_  (.A0(\ConfigFSM_inst._075_ ),
    .A1(\ConfigFSM_inst._076_ ),
    .S(\ConfigFSM_inst.FrameShiftState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._077_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._167_  (.A(\ConfigFSM_inst._077_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._005_ ));
 sky130_fd_sc_hd__xnor2_1 \ConfigFSM_inst._168_  (.A(\ConfigFSM_inst.FrameShiftState[0] ),
    .B(\ConfigFSM_inst.FrameShiftState[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._078_ ));
 sky130_fd_sc_hd__a22o_1 \ConfigFSM_inst._169_  (.A1(\ConfigFSM_inst.FrameShiftState[1] ),
    .A2(\ConfigFSM_inst._076_ ),
    .B1(\ConfigFSM_inst._075_ ),
    .B2(\ConfigFSM_inst._078_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._006_ ));
 sky130_fd_sc_hd__or3_2 \ConfigFSM_inst._170_  (.A(\ConfigFSM_inst.FrameShiftState[0] ),
    .B(\ConfigFSM_inst.FrameShiftState[1] ),
    .C(\ConfigFSM_inst.FrameShiftState[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._079_ ));
 sky130_fd_sc_hd__o21ai_1 \ConfigFSM_inst._171_  (.A1(\ConfigFSM_inst.FrameShiftState[0] ),
    .A2(\ConfigFSM_inst.FrameShiftState[1] ),
    .B1(\ConfigFSM_inst.FrameShiftState[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._080_ ));
 sky130_fd_sc_hd__nand2_1 \ConfigFSM_inst._172_  (.A(\ConfigFSM_inst._079_ ),
    .B(\ConfigFSM_inst._080_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._081_ ));
 sky130_fd_sc_hd__a22o_1 \ConfigFSM_inst._173_  (.A1(\ConfigFSM_inst.FrameShiftState[2] ),
    .A2(\ConfigFSM_inst._076_ ),
    .B1(\ConfigFSM_inst._075_ ),
    .B2(\ConfigFSM_inst._081_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._007_ ));
 sky130_fd_sc_hd__nor2_1 \ConfigFSM_inst._174_  (.A(\ConfigFSM_inst._076_ ),
    .B(\ConfigFSM_inst._079_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._082_ ));
 sky130_fd_sc_hd__o211a_1 \ConfigFSM_inst._175_  (.A1(\ConfigFSM_inst._070_ ),
    .A2(\ConfigFSM_inst._079_ ),
    .B1(\ConfigFSM_inst._057_ ),
    .C1(\ConfigFSM_inst.state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._083_ ));
 sky130_fd_sc_hd__o22a_1 \ConfigFSM_inst._176_  (.A1(\ConfigFSM_inst.FrameShiftState[3] ),
    .A2(\ConfigFSM_inst._082_ ),
    .B1(\ConfigFSM_inst._083_ ),
    .B2(\ConfigFSM_inst._076_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._008_ ));
 sky130_fd_sc_hd__o31a_1 \ConfigFSM_inst._177_  (.A1(\ConfigFSM_inst.FrameShiftState[3] ),
    .A2(\ConfigFSM_inst.FrameShiftState[4] ),
    .A3(\ConfigFSM_inst._079_ ),
    .B1(\ConfigFSM_inst.state[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._084_ ));
 sky130_fd_sc_hd__nor2_1 \ConfigFSM_inst._178_  (.A(\ConfigFSM_inst._074_ ),
    .B(\ConfigFSM_inst._084_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\ConfigFSM_inst._085_ ));
 sky130_fd_sc_hd__o31a_1 \ConfigFSM_inst._179_  (.A1(\ConfigFSM_inst.FrameShiftState[3] ),
    .A2(\ConfigFSM_inst._074_ ),
    .A3(\ConfigFSM_inst._079_ ),
    .B1(\ConfigFSM_inst.FrameShiftState[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._086_ ));
 sky130_fd_sc_hd__o21a_1 \ConfigFSM_inst._180_  (.A1(\ConfigFSM_inst._085_ ),
    .A2(\ConfigFSM_inst._086_ ),
    .B1(\ConfigFSM_inst._057_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._009_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._181_  (.A0(\ConfigFSM_inst.WriteData[0] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[0] ),
    .S(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._087_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._182_  (.A(\ConfigFSM_inst._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._010_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._183_  (.A0(\ConfigFSM_inst.WriteData[1] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[1] ),
    .S(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._088_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._184_  (.A(\ConfigFSM_inst._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._011_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._185_  (.A0(\ConfigFSM_inst.WriteData[2] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[2] ),
    .S(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._089_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._186_  (.A(\ConfigFSM_inst._089_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._012_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._187_  (.A0(\ConfigFSM_inst.WriteData[3] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[3] ),
    .S(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._090_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._188_  (.A(\ConfigFSM_inst._090_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._013_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._189_  (.A0(\ConfigFSM_inst.WriteData[4] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[4] ),
    .S(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._091_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._190_  (.A(\ConfigFSM_inst._091_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._014_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._191_  (.A0(\ConfigFSM_inst.WriteData[5] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[5] ),
    .S(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._092_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._192_  (.A(\ConfigFSM_inst._092_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._015_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._193_  (.A0(\ConfigFSM_inst.WriteData[6] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[6] ),
    .S(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._093_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._194_  (.A(\ConfigFSM_inst._093_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._016_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._195_  (.A0(\ConfigFSM_inst.WriteData[7] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[7] ),
    .S(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._094_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._196_  (.A(\ConfigFSM_inst._094_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._017_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._197_  (.A0(\ConfigFSM_inst.WriteData[8] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[8] ),
    .S(\ConfigFSM_inst._062_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._095_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._198_  (.A(\ConfigFSM_inst._095_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._018_ ));
 sky130_fd_sc_hd__clkbuf_4 \ConfigFSM_inst._199_  (.A(\ConfigFSM_inst._061_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._096_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._200_  (.A0(\ConfigFSM_inst.WriteData[9] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[9] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._097_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._201_  (.A(\ConfigFSM_inst._097_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._019_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._202_  (.A0(\ConfigFSM_inst.WriteData[10] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[10] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._098_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._203_  (.A(\ConfigFSM_inst._098_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._020_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._204_  (.A0(\ConfigFSM_inst.WriteData[11] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[11] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._099_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._205_  (.A(\ConfigFSM_inst._099_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._021_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._206_  (.A0(\ConfigFSM_inst.WriteData[12] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[12] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._100_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._207_  (.A(\ConfigFSM_inst._100_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._022_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._208_  (.A0(\ConfigFSM_inst.WriteData[13] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[13] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._101_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._209_  (.A(\ConfigFSM_inst._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._023_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._210_  (.A0(\ConfigFSM_inst.WriteData[14] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[14] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._102_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._211_  (.A(\ConfigFSM_inst._102_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._024_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._212_  (.A0(\ConfigFSM_inst.WriteData[15] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[15] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._103_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._213_  (.A(\ConfigFSM_inst._103_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._025_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._214_  (.A0(\ConfigFSM_inst.WriteData[16] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[16] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._104_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._215_  (.A(\ConfigFSM_inst._104_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._026_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._216_  (.A0(\ConfigFSM_inst.WriteData[17] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[17] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._105_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._217_  (.A(\ConfigFSM_inst._105_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._027_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._218_  (.A0(\ConfigFSM_inst.WriteData[18] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[18] ),
    .S(\ConfigFSM_inst._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._106_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._219_  (.A(\ConfigFSM_inst._106_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._028_ ));
 sky130_fd_sc_hd__clkbuf_4 \ConfigFSM_inst._220_  (.A(\ConfigFSM_inst._061_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._107_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._221_  (.A0(\ConfigFSM_inst.WriteData[19] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[19] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._108_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._222_  (.A(\ConfigFSM_inst._108_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._029_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._223_  (.A0(\ConfigFSM_inst.WriteData[21] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[21] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._109_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._224_  (.A(\ConfigFSM_inst._109_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._030_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._225_  (.A0(\ConfigFSM_inst.WriteData[22] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[22] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._110_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._226_  (.A(\ConfigFSM_inst._110_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._031_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._227_  (.A0(\ConfigFSM_inst.WriteData[23] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[23] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._111_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._228_  (.A(\ConfigFSM_inst._111_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._032_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._229_  (.A0(\ConfigFSM_inst.WriteData[24] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[24] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._112_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._230_  (.A(\ConfigFSM_inst._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._033_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._231_  (.A0(\ConfigFSM_inst.WriteData[25] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[25] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._113_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._232_  (.A(\ConfigFSM_inst._113_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._034_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._233_  (.A0(\ConfigFSM_inst.WriteData[26] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[26] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._114_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._234_  (.A(\ConfigFSM_inst._114_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._035_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._235_  (.A0(\ConfigFSM_inst.WriteData[27] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[27] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._115_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._236_  (.A(\ConfigFSM_inst._115_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._036_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._237_  (.A0(\ConfigFSM_inst.WriteData[28] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[28] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._116_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._238_  (.A(\ConfigFSM_inst._116_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._037_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._239_  (.A0(\ConfigFSM_inst.WriteData[29] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[29] ),
    .S(\ConfigFSM_inst._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._117_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._240_  (.A(\ConfigFSM_inst._117_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._038_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._241_  (.A0(\ConfigFSM_inst.WriteData[30] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[30] ),
    .S(\ConfigFSM_inst._061_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._118_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._242_  (.A(\ConfigFSM_inst._118_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._039_ ));
 sky130_fd_sc_hd__mux2_1 \ConfigFSM_inst._243_  (.A0(\ConfigFSM_inst.WriteData[31] ),
    .A1(\ConfigFSM_inst.FrameAddressRegister[31] ),
    .S(\ConfigFSM_inst._061_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._119_ ));
 sky130_fd_sc_hd__clkbuf_1 \ConfigFSM_inst._244_  (.A(\ConfigFSM_inst._119_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst._040_ ));
 sky130_fd_sc_hd__dfrtp_2 \ConfigFSM_inst._245_  (.CLK(net1),
    .D(\ConfigFSM_inst._005_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameShiftState[0] ));
 sky130_fd_sc_hd__dfrtp_2 \ConfigFSM_inst._246_  (.CLK(net1),
    .D(\ConfigFSM_inst._006_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameShiftState[1] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._247_  (.CLK(net1),
    .D(\ConfigFSM_inst._007_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameShiftState[2] ));
 sky130_fd_sc_hd__dfrtp_2 \ConfigFSM_inst._248_  (.CLK(net1),
    .D(\ConfigFSM_inst._008_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameShiftState[3] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._249_  (.CLK(net1),
    .D(\ConfigFSM_inst._009_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameShiftState[4] ));
 sky130_fd_sc_hd__dfstp_1 \ConfigFSM_inst._250_  (.CLK(net1),
    .D(\ConfigFSM_inst._002_ ),
    .SET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 \ConfigFSM_inst._251_  (.CLK(net1),
    .D(\ConfigFSM_inst._003_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._252_  (.CLK(net1),
    .D(\ConfigFSM_inst._004_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._253_  (.CLK(net1),
    .D(\ConfigFSM_inst._001_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._254_  (.CLK(net1),
    .D(\ConfigFSM_inst.FrameStrobe ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.oldFrameStrobe ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._255_  (.CLK(net1),
    .D(\ConfigFSM_inst._010_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[0] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._256_  (.CLK(net1),
    .D(\ConfigFSM_inst._011_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[1] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._257_  (.CLK(net1),
    .D(\ConfigFSM_inst._012_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[2] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._258_  (.CLK(net1),
    .D(\ConfigFSM_inst._013_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[3] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._259_  (.CLK(net1),
    .D(\ConfigFSM_inst._014_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[4] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._260_  (.CLK(net1),
    .D(\ConfigFSM_inst._015_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[5] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._261_  (.CLK(net1),
    .D(\ConfigFSM_inst._016_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[6] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._262_  (.CLK(net1),
    .D(\ConfigFSM_inst._017_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[7] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._263_  (.CLK(net1),
    .D(\ConfigFSM_inst._018_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[8] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._264_  (.CLK(net1),
    .D(\ConfigFSM_inst._019_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[9] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._265_  (.CLK(net1),
    .D(\ConfigFSM_inst._020_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[10] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._266_  (.CLK(net1),
    .D(\ConfigFSM_inst._021_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[11] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._267_  (.CLK(net1),
    .D(\ConfigFSM_inst._022_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[12] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._268_  (.CLK(net1),
    .D(\ConfigFSM_inst._023_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[13] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._269_  (.CLK(net1),
    .D(\ConfigFSM_inst._024_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[14] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._270_  (.CLK(net1),
    .D(\ConfigFSM_inst._025_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[15] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._271_  (.CLK(net1),
    .D(\ConfigFSM_inst._026_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[16] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._272_  (.CLK(net1),
    .D(\ConfigFSM_inst._027_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[17] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._273_  (.CLK(net1),
    .D(\ConfigFSM_inst._028_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[18] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._274_  (.CLK(net1),
    .D(\ConfigFSM_inst._029_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[19] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._275_  (.CLK(net1),
    .D(\ConfigFSM_inst._030_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[21] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._276_  (.CLK(net1),
    .D(\ConfigFSM_inst._031_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[22] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._277_  (.CLK(net1),
    .D(\ConfigFSM_inst._032_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[23] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._278_  (.CLK(net1),
    .D(\ConfigFSM_inst._033_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[24] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._279_  (.CLK(net1),
    .D(\ConfigFSM_inst._034_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[25] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._280_  (.CLK(net1),
    .D(\ConfigFSM_inst._035_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[26] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._281_  (.CLK(net1),
    .D(\ConfigFSM_inst._036_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[27] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._282_  (.CLK(net1),
    .D(\ConfigFSM_inst._037_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[28] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._283_  (.CLK(net1),
    .D(\ConfigFSM_inst._038_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[29] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._284_  (.CLK(net1),
    .D(\ConfigFSM_inst._039_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[30] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._285_  (.CLK(net1),
    .D(\ConfigFSM_inst._040_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameAddressRegister[31] ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._286_  (.CLK(net1),
    .D(\ConfigFSM_inst._000_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.FrameStrobe ));
 sky130_fd_sc_hd__dfrtp_1 \ConfigFSM_inst._287_  (.CLK(net1),
    .D(\ConfigFSM_inst.FSM_Reset ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigFSM_inst.old_reset ));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_371 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_480 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_336 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_370 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_404 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_478 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_482 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_486 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_375 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_319 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_433 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_355 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_463 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_463 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_471 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_310 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_400 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_452 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_476 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_480 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_484 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_368 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_463 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_471 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_383 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_339 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_343 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_450 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_454 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_433 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_437 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_320 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_347 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_351 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_381 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_478 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_482 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_486 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_339 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_343 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_347 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_351 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_355 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_394 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_404 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_427 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_403 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_355 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_400 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_404 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_478 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_482 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_486 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_448 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_452 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_392 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_344 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_371 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_368 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_420 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_471 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_479 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_483 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_336 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_371 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_375 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_348 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_423 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_338 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_463 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_471 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_450 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_454 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_424 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_480 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_336 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_375 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_394 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_316 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_340 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_403 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_407 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_463 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_471 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_366 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_400 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_404 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_372 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_407 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_481 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_485 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_471 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_479 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_483 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0589_  (.A(\INST_config_UART.blink[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0031_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._0590_  (.A(\INST_config_UART.PresentState[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0192_ ));
 sky130_fd_sc_hd__and2_1 \INST_config_UART._0591_  (.A(\INST_config_UART.ComTick ),
    .B(\INST_config_UART.ComState[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0193_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0592_  (.A(\INST_config_UART.TimeToSend ),
    .B(\INST_config_UART._0193_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0194_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0593_  (.A(\INST_config_UART.ComTick ),
    .B(\INST_config_UART.ComState[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0195_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0594_  (.A(\INST_config_UART.TimeToSend ),
    .B(\INST_config_UART._0195_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0196_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0595_  (.A1(\INST_config_UART._0192_ ),
    .A2(\INST_config_UART._0194_ ),
    .B1(\INST_config_UART._0196_ ),
    .B2(\INST_config_UART.PresentState[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0026_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0596_  (.A(\INST_config_UART.ComTick ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0197_ ));
 sky130_fd_sc_hd__and2b_1 \INST_config_UART._0597_  (.A_N(\INST_config_UART.RxLocal ),
    .B(\INST_config_UART.ComState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0198_ ));
 sky130_fd_sc_hd__a21o_1 \INST_config_UART._0598_  (.A1(\INST_config_UART._0197_ ),
    .A2(\INST_config_UART.ComState[6] ),
    .B1(\INST_config_UART._0198_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0020_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0599_  (.A(\INST_config_UART._0198_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0199_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0600_  (.A(\INST_config_UART.Command[1] ),
    .B(\INST_config_UART.Command[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0200_ ));
 sky130_fd_sc_hd__or4_1 \INST_config_UART._0601_  (.A(\INST_config_UART.ID_Reg[23] ),
    .B(\INST_config_UART.ID_Reg[22] ),
    .C(\INST_config_UART.Command[3] ),
    .D(\INST_config_UART.Command[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0201_ ));
 sky130_fd_sc_hd__or4_1 \INST_config_UART._0602_  (.A(\INST_config_UART.Command[5] ),
    .B(\INST_config_UART.Command[4] ),
    .C(\INST_config_UART.Command[6] ),
    .D(\INST_config_UART._0201_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0202_ ));
 sky130_fd_sc_hd__and4b_1 \INST_config_UART._0603_  (.A_N(\INST_config_UART.ID_Reg[8] ),
    .B(\INST_config_UART.ID_Reg[9] ),
    .C(\INST_config_UART.ID_Reg[7] ),
    .D(\INST_config_UART.ID_Reg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0203_ ));
 sky130_fd_sc_hd__and4bb_1 \INST_config_UART._0604_  (.A_N(\INST_config_UART.ID_Reg[10] ),
    .B_N(\INST_config_UART.ID_Reg[12] ),
    .C(\INST_config_UART.ID_Reg[13] ),
    .D(\INST_config_UART.ID_Reg[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0204_ ));
 sky130_fd_sc_hd__and4_1 \INST_config_UART._0605_  (.A(\INST_config_UART.ID_Reg[3] ),
    .B(\INST_config_UART.ID_Reg[2] ),
    .C(\INST_config_UART.ID_Reg[5] ),
    .D(\INST_config_UART.ID_Reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0205_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0606_  (.A(\INST_config_UART.ID_Reg[1] ),
    .B(\INST_config_UART.ID_Reg[0] ),
    .C(\INST_config_UART._0205_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0206_ ));
 sky130_fd_sc_hd__or4_1 \INST_config_UART._0607_  (.A(\INST_config_UART.ID_Reg[19] ),
    .B(\INST_config_UART.ID_Reg[18] ),
    .C(\INST_config_UART.ID_Reg[21] ),
    .D(\INST_config_UART.ID_Reg[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0207_ ));
 sky130_fd_sc_hd__or4b_1 \INST_config_UART._0608_  (.A(\INST_config_UART.ID_Reg[14] ),
    .B(\INST_config_UART.ID_Reg[17] ),
    .C(\INST_config_UART.ID_Reg[16] ),
    .D_N(\INST_config_UART.ID_Reg[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0208_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0609_  (.A(\INST_config_UART._0207_ ),
    .B(\INST_config_UART._0208_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0209_ ));
 sky130_fd_sc_hd__and4_1 \INST_config_UART._0610_  (.A(\INST_config_UART._0203_ ),
    .B(\INST_config_UART._0204_ ),
    .C(\INST_config_UART._0206_ ),
    .D(\INST_config_UART._0209_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0210_ ));
 sky130_fd_sc_hd__or3b_2 \INST_config_UART._0611_  (.A(\INST_config_UART._0200_ ),
    .B(\INST_config_UART._0202_ ),
    .C_N(\INST_config_UART._0210_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0211_ ));
 sky130_fd_sc_hd__or4_1 \INST_config_UART._0612_  (.A(net39),
    .B(\INST_config_UART._0192_ ),
    .C(\INST_config_UART.PresentState[2] ),
    .D(\INST_config_UART.PresentState[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0212_ ));
 sky130_fd_sc_hd__o21a_1 \INST_config_UART._0613_  (.A1(\INST_config_UART.PresentState[6] ),
    .A2(\INST_config_UART._0212_ ),
    .B1(\INST_config_UART.TimeToSend ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0213_ ));
 sky130_fd_sc_hd__a221o_1 \INST_config_UART._0614_  (.A1(\INST_config_UART.PresentState[0] ),
    .A2(\INST_config_UART._0199_ ),
    .B1(\INST_config_UART._0211_ ),
    .B2(\INST_config_UART.PresentState[5] ),
    .C1(\INST_config_UART._0213_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0025_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._0615_  (.A(\INST_config_UART.ByteWriteStrobe ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0214_ ));
 sky130_fd_sc_hd__nand2_4 \INST_config_UART._0616_  (.A(\INST_config_UART._0214_ ),
    .B(\INST_config_UART.GetWordState[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0215_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._0617_  (.A(\INST_config_UART.ByteWriteStrobe ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0216_ ));
 sky130_fd_sc_hd__or2b_1 \INST_config_UART._0618_  (.A(\INST_config_UART._0216_ ),
    .B_N(\INST_config_UART.GetWordState[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0217_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0619_  (.A1(\INST_config_UART._0215_ ),
    .A2(\INST_config_UART._0217_ ),
    .B1(\INST_config_UART.PresentState[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0024_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0620_  (.A1(\INST_config_UART.PresentState[2] ),
    .A2(\INST_config_UART._0194_ ),
    .B1(\INST_config_UART._0196_ ),
    .B2(\INST_config_UART.PresentState[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0027_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0621_  (.A1(\INST_config_UART.PresentState[6] ),
    .A2(\INST_config_UART._0194_ ),
    .B1(\INST_config_UART._0196_ ),
    .B2(\INST_config_UART.PresentState[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0030_ ));
 sky130_fd_sc_hd__buf_4 \INST_config_UART._0622_  (.A(\INST_config_UART.ReceivedWord[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0218_ ));
 sky130_fd_sc_hd__or4bb_2 \INST_config_UART._0623_  (.A(\INST_config_UART.ReceivedWord[7] ),
    .B(\INST_config_UART.ReceivedWord[6] ),
    .C_N(\INST_config_UART.ReceivedWord[5] ),
    .D_N(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0219_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0624_  (.A(\INST_config_UART._0218_ ),
    .B(\INST_config_UART._0219_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0220_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._0625_  (.A(\INST_config_UART.ReceivedWord[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0221_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._0626_  (.A(\INST_config_UART.ReceivedWord[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0222_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._0627_  (.A(\INST_config_UART.ReceivedWord[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0223_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0628_  (.A(\INST_config_UART._0222_ ),
    .B(\INST_config_UART._0223_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0224_ ));
 sky130_fd_sc_hd__or3b_1 \INST_config_UART._0629_  (.A(\INST_config_UART.ReceivedWord[4] ),
    .B(\INST_config_UART.ReceivedWord[7] ),
    .C_N(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0225_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0630_  (.A(\INST_config_UART._0222_ ),
    .B(\INST_config_UART._0223_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0226_ ));
 sky130_fd_sc_hd__or3b_2 \INST_config_UART._0631_  (.A(\INST_config_UART._0224_ ),
    .B(\INST_config_UART._0225_ ),
    .C_N(\INST_config_UART._0226_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0227_ ));
 sky130_fd_sc_hd__or4b_2 \INST_config_UART._0632_  (.A(\INST_config_UART._0222_ ),
    .B(\INST_config_UART._0221_ ),
    .C(\INST_config_UART._0219_ ),
    .D_N(\INST_config_UART.ReceivedWord[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0228_ ));
 sky130_fd_sc_hd__or2b_1 \INST_config_UART._0633_  (.A(\INST_config_UART.ReceivedWord[3] ),
    .B_N(\INST_config_UART._0221_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0229_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0634_  (.A1(\INST_config_UART.ReceivedWord[3] ),
    .A2(\INST_config_UART.ReceivedWord[2] ),
    .B1(\INST_config_UART.ReceivedWord[1] ),
    .C1(\INST_config_UART.ReceivedWord[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0230_ ));
 sky130_fd_sc_hd__a211o_1 \INST_config_UART._0635_  (.A1(\INST_config_UART._0226_ ),
    .A2(\INST_config_UART._0229_ ),
    .B1(\INST_config_UART._0230_ ),
    .C1(\INST_config_UART._0225_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0231_ ));
 sky130_fd_sc_hd__o311ai_4 \INST_config_UART._0636_  (.A1(\INST_config_UART._0218_ ),
    .A2(\INST_config_UART._0221_ ),
    .A3(\INST_config_UART._0227_ ),
    .B1(\INST_config_UART._0228_ ),
    .C1(\INST_config_UART._0231_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0232_ ));
 sky130_fd_sc_hd__o21ai_2 \INST_config_UART._0637_  (.A1(\INST_config_UART._0220_ ),
    .A2(\INST_config_UART._0232_ ),
    .B1(\INST_config_UART._0193_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0233_ ));
 sky130_fd_sc_hd__nor2_4 \INST_config_UART._0638_  (.A(\INST_config_UART.ReceiveState ),
    .B(\INST_config_UART._0233_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0014_ ));
 sky130_fd_sc_hd__nand2_4 \INST_config_UART._0639_  (.A(\INST_config_UART._0214_ ),
    .B(\INST_config_UART.GetWordState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0234_ ));
 sky130_fd_sc_hd__or2b_1 \INST_config_UART._0640_  (.A(\INST_config_UART._0216_ ),
    .B_N(\INST_config_UART.GetWordState[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0235_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0641_  (.A1(\INST_config_UART._0234_ ),
    .A2(\INST_config_UART._0235_ ),
    .B1(\INST_config_UART.PresentState[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0023_ ));
 sky130_fd_sc_hd__nand2_4 \INST_config_UART._0642_  (.A(\INST_config_UART._0214_ ),
    .B(\INST_config_UART.GetWordState[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0236_ ));
 sky130_fd_sc_hd__or2b_1 \INST_config_UART._0643_  (.A(\INST_config_UART.ByteWriteStrobe ),
    .B_N(\INST_config_UART.GetWordState[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0237_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0644_  (.A1(\INST_config_UART._0236_ ),
    .A2(\INST_config_UART._0237_ ),
    .B1(\INST_config_UART.PresentState[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0022_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0645_  (.A(\INST_config_UART.GetWordState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0238_ ));
 sky130_fd_sc_hd__and2_1 \INST_config_UART._0646_  (.A(\INST_config_UART.ByteWriteStrobe ),
    .B(\INST_config_UART.GetWordState[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0239_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._0647_  (.A(\INST_config_UART._0239_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0017_ ));
 sky130_fd_sc_hd__nor2_4 \INST_config_UART._0648_  (.A(\INST_config_UART.PresentState[5] ),
    .B(\INST_config_UART._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0240_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0649_  (.A1(\INST_config_UART._0214_ ),
    .A2(\INST_config_UART._0238_ ),
    .B1(\INST_config_UART._0240_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0021_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0650_  (.A1(\INST_config_UART.PresentState[4] ),
    .A2(\INST_config_UART._0194_ ),
    .B1(\INST_config_UART._0198_ ),
    .B2(\INST_config_UART.PresentState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0029_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0651_  (.A(\INST_config_UART.PresentState[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0241_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._0652_  (.A(\INST_config_UART._0241_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0242_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._0653_  (.A(\INST_config_UART._0242_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0243_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0654_  (.A(\INST_config_UART.TimeToSend ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0244_ ));
 sky130_fd_sc_hd__a2bb2o_1 \INST_config_UART._0655_  (.A1_N(\INST_config_UART._0243_ ),
    .A2_N(\INST_config_UART._0211_ ),
    .B1(net39),
    .B2(\INST_config_UART._0244_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0028_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0656_  (.A(\INST_config_UART.RxLocal ),
    .B(\INST_config_UART.ComState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0245_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0657_  (.A(\INST_config_UART._0195_ ),
    .B(\INST_config_UART._0245_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0019_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._0658_  (.A(\INST_config_UART.Command[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0246_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._0659_  (.A(\INST_config_UART._0246_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0247_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0660_  (.A0(\INST_config_UART.LocalWriteStrobe ),
    .A1(\INST_config_UART.HexWriteStrobe ),
    .S(\INST_config_UART._0247_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0248_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0661_  (.A(\INST_config_UART._0248_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0000_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0662_  (.A(net39),
    .B(\INST_config_UART._0242_ ),
    .C(\INST_config_UART._0193_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0249_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0663_  (.A(\INST_config_UART._0249_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0015_ ));
 sky130_fd_sc_hd__clkbuf_2 \INST_config_UART._0664_  (.A(\INST_config_UART.ComState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0250_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._0665_  (.A(\INST_config_UART._0250_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0251_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._0666_  (.A(\INST_config_UART.ComCount[1] ),
    .B(\INST_config_UART.ComCount[0] ),
    .C(\INST_config_UART.ComCount[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0252_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0667_  (.A(\INST_config_UART.ComCount[3] ),
    .B(\INST_config_UART._0252_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0253_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._0668_  (.A(\INST_config_UART.ComCount[5] ),
    .B(\INST_config_UART.ComCount[4] ),
    .C(\INST_config_UART._0253_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0254_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0669_  (.A(\INST_config_UART.ComCount[6] ),
    .B(\INST_config_UART._0254_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0255_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._0670_  (.A(\INST_config_UART.ComCount[7] ),
    .B(\INST_config_UART.ComCount[8] ),
    .C(\INST_config_UART._0255_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0256_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0671_  (.A(\INST_config_UART.ComCount[9] ),
    .B(\INST_config_UART._0256_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0257_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0672_  (.A(\INST_config_UART.ComCount[10] ),
    .B(\INST_config_UART._0257_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0258_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0673_  (.A(\INST_config_UART.ComCount[11] ),
    .B(\INST_config_UART._0258_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0259_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0674_  (.A(\INST_config_UART._0251_ ),
    .B(\INST_config_UART._0259_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0013_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0675_  (.A(\INST_config_UART._0251_ ),
    .B(\INST_config_UART.ComCount[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0001_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0676_  (.A(\INST_config_UART.ComCount[1] ),
    .B(\INST_config_UART.ComCount[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0260_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0677_  (.A(\INST_config_UART.ComCount[1] ),
    .B(\INST_config_UART.ComCount[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0261_ ));
 sky130_fd_sc_hd__nand2b_1 \INST_config_UART._0678_  (.A_N(\INST_config_UART._0250_ ),
    .B(\INST_config_UART._0259_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0262_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0679_  (.A1(\INST_config_UART._0260_ ),
    .A2(\INST_config_UART._0261_ ),
    .B1(\INST_config_UART._0262_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0004_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0680_  (.A(\INST_config_UART.ComCount[2] ),
    .B(\INST_config_UART._0260_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0263_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0681_  (.A(\INST_config_UART._0252_ ),
    .B(\INST_config_UART._0263_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0264_ ));
 sky130_fd_sc_hd__a21o_1 \INST_config_UART._0682_  (.A1(\INST_config_UART._0259_ ),
    .A2(\INST_config_UART._0264_ ),
    .B1(\INST_config_UART._0251_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0005_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0683_  (.A1(\INST_config_UART.ComCount[3] ),
    .A2(\INST_config_UART._0252_ ),
    .B1(\INST_config_UART._0251_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0265_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0684_  (.A(\INST_config_UART._0253_ ),
    .B(\INST_config_UART._0265_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0006_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0685_  (.A(\INST_config_UART.ComCount[4] ),
    .B(\INST_config_UART._0253_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0266_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0686_  (.A(\INST_config_UART.ComCount[4] ),
    .B(\INST_config_UART._0253_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0267_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0687_  (.A1(\INST_config_UART._0266_ ),
    .A2(\INST_config_UART._0267_ ),
    .B1(\INST_config_UART._0251_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0007_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0688_  (.A1(\INST_config_UART.ComCount[4] ),
    .A2(\INST_config_UART._0253_ ),
    .B1(\INST_config_UART.ComCount[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0268_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0689_  (.A(\INST_config_UART._0254_ ),
    .B(\INST_config_UART._0268_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0269_ ));
 sky130_fd_sc_hd__a21o_1 \INST_config_UART._0690_  (.A1(\INST_config_UART._0259_ ),
    .A2(\INST_config_UART._0269_ ),
    .B1(\INST_config_UART._0251_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0008_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0691_  (.A1(\INST_config_UART.ComCount[6] ),
    .A2(\INST_config_UART._0254_ ),
    .B1(\INST_config_UART._0251_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0270_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0692_  (.A(\INST_config_UART._0255_ ),
    .B(\INST_config_UART._0270_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0009_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0693_  (.A(\INST_config_UART.ComCount[7] ),
    .B(\INST_config_UART._0255_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0271_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0694_  (.A(\INST_config_UART.ComCount[7] ),
    .B(\INST_config_UART._0255_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0272_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0695_  (.A1(\INST_config_UART._0271_ ),
    .A2(\INST_config_UART._0272_ ),
    .B1(\INST_config_UART._0251_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0010_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0696_  (.A1(\INST_config_UART.ComCount[7] ),
    .A2(\INST_config_UART._0255_ ),
    .B1(\INST_config_UART.ComCount[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0273_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0697_  (.A1(\INST_config_UART._0256_ ),
    .A2(\INST_config_UART._0273_ ),
    .B1(\INST_config_UART._0262_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0011_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0698_  (.A(\INST_config_UART.ComCount[9] ),
    .B(\INST_config_UART._0256_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0274_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0699_  (.A1(\INST_config_UART._0257_ ),
    .A2(\INST_config_UART._0274_ ),
    .B1(\INST_config_UART._0262_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0012_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0700_  (.A(\INST_config_UART.ComCount[10] ),
    .B(\INST_config_UART._0257_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0275_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0701_  (.A1(\INST_config_UART._0258_ ),
    .A2(\INST_config_UART._0275_ ),
    .B1(\INST_config_UART._0262_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0002_ ));
 sky130_fd_sc_hd__and3b_1 \INST_config_UART._0702_  (.A_N(\INST_config_UART._0251_ ),
    .B(\INST_config_UART.ComCount[11] ),
    .C(\INST_config_UART._0258_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0276_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0703_  (.A(\INST_config_UART._0276_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0003_ ));
 sky130_fd_sc_hd__or4_1 \INST_config_UART._0704_  (.A(\INST_config_UART.PresentState[2] ),
    .B(\INST_config_UART.PresentState[4] ),
    .C(\INST_config_UART.PresentState[5] ),
    .D(\INST_config_UART.PresentState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0277_ ));
 sky130_fd_sc_hd__or4_1 \INST_config_UART._0705_  (.A(\INST_config_UART.PresentState[6] ),
    .B(\INST_config_UART._0192_ ),
    .C(\INST_config_UART._0233_ ),
    .D(\INST_config_UART._0277_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0278_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0706_  (.A(\INST_config_UART._0278_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0016_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0707_  (.A(\INST_config_UART._0244_ ),
    .B(\INST_config_UART._0192_ ),
    .C(\INST_config_UART._0193_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0279_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0708_  (.A(\INST_config_UART._0279_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0018_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0709_  (.A(\INST_config_UART.blink[0] ),
    .B(\INST_config_UART.blink[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0042_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._0710_  (.A(\INST_config_UART.blink[0] ),
    .B(\INST_config_UART.blink[1] ),
    .C(\INST_config_UART.blink[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0280_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0711_  (.A1(\INST_config_UART.blink[0] ),
    .A2(\INST_config_UART.blink[1] ),
    .B1(\INST_config_UART.blink[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0281_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0712_  (.A(\INST_config_UART._0280_ ),
    .B(\INST_config_UART._0281_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0046_ ));
 sky130_fd_sc_hd__or4_2 \INST_config_UART._0713_  (.A(\INST_config_UART.blink[0] ),
    .B(\INST_config_UART.blink[1] ),
    .C(\INST_config_UART.blink[2] ),
    .D(\INST_config_UART.blink[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0282_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0714_  (.A(\INST_config_UART.blink[3] ),
    .B(\INST_config_UART._0280_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0283_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0715_  (.A(\INST_config_UART._0282_ ),
    .B(\INST_config_UART._0283_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0047_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0716_  (.A(\INST_config_UART.blink[4] ),
    .B(\INST_config_UART._0282_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0284_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0717_  (.A(\INST_config_UART.blink[4] ),
    .B(\INST_config_UART._0282_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0285_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0718_  (.A(\INST_config_UART._0284_ ),
    .B(\INST_config_UART._0285_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0048_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0719_  (.A(\INST_config_UART.blink[5] ),
    .B(\INST_config_UART._0284_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0049_ ));
 sky130_fd_sc_hd__or4_2 \INST_config_UART._0720_  (.A(\INST_config_UART.blink[4] ),
    .B(\INST_config_UART.blink[5] ),
    .C(\INST_config_UART.blink[6] ),
    .D(\INST_config_UART._0282_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0286_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0721_  (.A1(\INST_config_UART.blink[5] ),
    .A2(\INST_config_UART._0284_ ),
    .B1(\INST_config_UART.blink[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0287_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0722_  (.A(\INST_config_UART._0286_ ),
    .B(\INST_config_UART._0287_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0050_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0723_  (.A(\INST_config_UART.blink[7] ),
    .B(\INST_config_UART._0286_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0051_ ));
 sky130_fd_sc_hd__or3_2 \INST_config_UART._0724_  (.A(\INST_config_UART.blink[7] ),
    .B(\INST_config_UART.blink[8] ),
    .C(\INST_config_UART._0286_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0288_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0725_  (.A1(\INST_config_UART.blink[7] ),
    .A2(\INST_config_UART._0286_ ),
    .B1(\INST_config_UART.blink[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0289_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0726_  (.A(\INST_config_UART._0288_ ),
    .B(\INST_config_UART._0289_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0052_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0727_  (.A(\INST_config_UART.blink[9] ),
    .B(\INST_config_UART._0288_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0053_ ));
 sky130_fd_sc_hd__or3_2 \INST_config_UART._0728_  (.A(\INST_config_UART.blink[9] ),
    .B(\INST_config_UART.blink[10] ),
    .C(\INST_config_UART._0288_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0290_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0729_  (.A1(\INST_config_UART.blink[9] ),
    .A2(\INST_config_UART._0288_ ),
    .B1(\INST_config_UART.blink[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0291_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0730_  (.A(\INST_config_UART._0290_ ),
    .B(\INST_config_UART._0291_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0032_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0731_  (.A(\INST_config_UART.blink[11] ),
    .B(\INST_config_UART._0290_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0292_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0732_  (.A(\INST_config_UART.blink[11] ),
    .B(\INST_config_UART._0290_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0293_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0733_  (.A(\INST_config_UART._0292_ ),
    .B(\INST_config_UART._0293_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0033_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0734_  (.A(\INST_config_UART.blink[12] ),
    .B(\INST_config_UART._0292_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0034_ ));
 sky130_fd_sc_hd__or4_2 \INST_config_UART._0735_  (.A(\INST_config_UART.blink[11] ),
    .B(\INST_config_UART.blink[12] ),
    .C(\INST_config_UART.blink[13] ),
    .D(\INST_config_UART._0290_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0294_ ));
 sky130_fd_sc_hd__o31ai_1 \INST_config_UART._0736_  (.A1(\INST_config_UART.blink[11] ),
    .A2(\INST_config_UART.blink[12] ),
    .A3(\INST_config_UART._0290_ ),
    .B1(\INST_config_UART.blink[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0295_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0737_  (.A(\INST_config_UART._0294_ ),
    .B(\INST_config_UART._0295_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0035_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0738_  (.A(\INST_config_UART.blink[14] ),
    .B(\INST_config_UART._0294_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0296_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0739_  (.A(\INST_config_UART.blink[14] ),
    .B(\INST_config_UART._0294_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0297_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0740_  (.A(\INST_config_UART._0296_ ),
    .B(\INST_config_UART._0297_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0036_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0741_  (.A(\INST_config_UART.blink[15] ),
    .B(\INST_config_UART._0296_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0037_ ));
 sky130_fd_sc_hd__or4_2 \INST_config_UART._0742_  (.A(\INST_config_UART.blink[14] ),
    .B(\INST_config_UART.blink[15] ),
    .C(\INST_config_UART.blink[16] ),
    .D(\INST_config_UART._0294_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0298_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0743_  (.A1(\INST_config_UART.blink[15] ),
    .A2(\INST_config_UART._0296_ ),
    .B1(\INST_config_UART.blink[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0299_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0744_  (.A(\INST_config_UART._0298_ ),
    .B(\INST_config_UART._0299_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0038_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0745_  (.A(\INST_config_UART.blink[17] ),
    .B(\INST_config_UART._0298_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0039_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._0746_  (.A(\INST_config_UART.blink[17] ),
    .B(\INST_config_UART.blink[18] ),
    .C(\INST_config_UART._0298_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0300_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0747_  (.A1(\INST_config_UART.blink[17] ),
    .A2(\INST_config_UART._0298_ ),
    .B1(\INST_config_UART.blink[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0301_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0748_  (.A(\INST_config_UART._0300_ ),
    .B(\INST_config_UART._0301_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0040_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0749_  (.A(\INST_config_UART.blink[19] ),
    .B(\INST_config_UART._0300_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0302_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0750_  (.A(\INST_config_UART.blink[19] ),
    .B(\INST_config_UART._0300_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0303_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0751_  (.A(\INST_config_UART._0302_ ),
    .B(\INST_config_UART._0303_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0041_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0752_  (.A(\INST_config_UART.blink[20] ),
    .B(\INST_config_UART._0302_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0043_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._0753_  (.A(\INST_config_UART.blink[20] ),
    .B(\INST_config_UART.blink[21] ),
    .C(\INST_config_UART._0302_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0304_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0754_  (.A1(\INST_config_UART.blink[20] ),
    .A2(\INST_config_UART._0302_ ),
    .B1(\INST_config_UART.blink[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0305_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0755_  (.A(\INST_config_UART._0304_ ),
    .B(\INST_config_UART._0305_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0044_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._0756_  (.A(\INST_config_UART.blink[22] ),
    .B(\INST_config_UART._0304_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0045_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0757_  (.A(\INST_config_UART._0197_ ),
    .B(\INST_config_UART.ComState[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0306_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0758_  (.A1(\INST_config_UART.ComState[0] ),
    .A2(\INST_config_UART.ComState[7] ),
    .B1(\INST_config_UART._0245_ ),
    .C1(\INST_config_UART._0306_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0307_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0759_  (.A0(\INST_config_UART.ReceivedWord[7] ),
    .A1(\INST_config_UART.RxLocal ),
    .S(\INST_config_UART._0307_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0308_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0760_  (.A(\INST_config_UART._0308_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0054_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0761_  (.A(\INST_config_UART._0197_ ),
    .B(\INST_config_UART.ComState[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0309_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0762_  (.A1(\INST_config_UART.ComState[0] ),
    .A2(\INST_config_UART.ComState[2] ),
    .B1(\INST_config_UART._0245_ ),
    .C1(\INST_config_UART._0309_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0310_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0763_  (.A0(\INST_config_UART._0221_ ),
    .A1(\INST_config_UART.RxLocal ),
    .S(\INST_config_UART._0310_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0311_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0764_  (.A(\INST_config_UART._0311_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0055_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0765_  (.A(\INST_config_UART._0246_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0312_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0766_  (.A(\INST_config_UART._0247_ ),
    .B(\INST_config_UART.Data_Reg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0313_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0767_  (.A1(\INST_config_UART._0312_ ),
    .A2(\INST_config_UART.HexData[0] ),
    .B1(\INST_config_UART._0313_ ),
    .C1(\INST_config_UART._0242_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0314_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0768_  (.A1(\INST_config_UART.WriteData[0] ),
    .A2(\INST_config_UART._0240_ ),
    .B1(\INST_config_UART._0314_ ),
    .B2(\INST_config_UART._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0056_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0769_  (.A(\INST_config_UART._0247_ ),
    .B(\INST_config_UART.Data_Reg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0315_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0770_  (.A1(\INST_config_UART._0312_ ),
    .A2(\INST_config_UART.HexData[1] ),
    .B1(\INST_config_UART._0315_ ),
    .C1(\INST_config_UART._0242_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0316_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0771_  (.A1(\INST_config_UART.WriteData[1] ),
    .A2(\INST_config_UART._0240_ ),
    .B1(\INST_config_UART._0316_ ),
    .B2(\INST_config_UART._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0057_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0772_  (.A(\INST_config_UART._0247_ ),
    .B(\INST_config_UART.Data_Reg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0317_ ));
 sky130_fd_sc_hd__o211a_2 \INST_config_UART._0773_  (.A1(\INST_config_UART._0312_ ),
    .A2(\INST_config_UART.HexData[2] ),
    .B1(\INST_config_UART._0317_ ),
    .C1(\INST_config_UART._0241_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0318_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0774_  (.A1(\INST_config_UART.WriteData[2] ),
    .A2(\INST_config_UART._0240_ ),
    .B1(\INST_config_UART._0318_ ),
    .B2(\INST_config_UART._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0058_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0775_  (.A(\INST_config_UART._0247_ ),
    .B(\INST_config_UART.Data_Reg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0319_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0776_  (.A1(\INST_config_UART._0312_ ),
    .A2(\INST_config_UART.HexData[3] ),
    .B1(\INST_config_UART._0319_ ),
    .C1(\INST_config_UART._0241_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0320_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0777_  (.A1(\INST_config_UART.WriteData[3] ),
    .A2(\INST_config_UART._0240_ ),
    .B1(\INST_config_UART._0320_ ),
    .B2(\INST_config_UART._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0059_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0778_  (.A(\INST_config_UART._0247_ ),
    .B(\INST_config_UART.Data_Reg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0321_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0779_  (.A1(\INST_config_UART._0312_ ),
    .A2(\INST_config_UART.HexData[4] ),
    .B1(\INST_config_UART._0321_ ),
    .C1(\INST_config_UART._0241_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0322_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0780_  (.A1(\INST_config_UART.WriteData[4] ),
    .A2(\INST_config_UART._0240_ ),
    .B1(\INST_config_UART._0322_ ),
    .B2(\INST_config_UART._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0060_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0781_  (.A(\INST_config_UART._0247_ ),
    .B(\INST_config_UART.Data_Reg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0323_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0782_  (.A1(\INST_config_UART._0312_ ),
    .A2(\INST_config_UART.HexData[5] ),
    .B1(\INST_config_UART._0323_ ),
    .C1(\INST_config_UART._0241_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0324_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0783_  (.A1(\INST_config_UART.WriteData[5] ),
    .A2(\INST_config_UART._0240_ ),
    .B1(\INST_config_UART._0324_ ),
    .B2(\INST_config_UART._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0061_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0784_  (.A(\INST_config_UART._0247_ ),
    .B(\INST_config_UART.Data_Reg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0325_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0785_  (.A1(\INST_config_UART._0312_ ),
    .A2(\INST_config_UART.HexData[6] ),
    .B1(\INST_config_UART._0325_ ),
    .C1(\INST_config_UART._0241_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0326_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0786_  (.A1(\INST_config_UART.WriteData[6] ),
    .A2(\INST_config_UART._0240_ ),
    .B1(\INST_config_UART._0326_ ),
    .B2(\INST_config_UART._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0062_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0787_  (.A(\INST_config_UART._0247_ ),
    .B(\INST_config_UART.Data_Reg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0327_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._0788_  (.A1(\INST_config_UART._0312_ ),
    .A2(\INST_config_UART.HexData[7] ),
    .B1(\INST_config_UART._0327_ ),
    .C1(\INST_config_UART._0241_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0328_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._0789_  (.A1(\INST_config_UART.WriteData[7] ),
    .A2(\INST_config_UART._0240_ ),
    .B1(\INST_config_UART._0328_ ),
    .B2(\INST_config_UART._0017_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0063_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0790_  (.A(\INST_config_UART._0214_ ),
    .B(\INST_config_UART.GetWordState[2] ),
    .C(\INST_config_UART._0314_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0329_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0791_  (.A1(\INST_config_UART._0243_ ),
    .A2(\INST_config_UART.WriteData[16] ),
    .A3(\INST_config_UART._0236_ ),
    .B1(\INST_config_UART._0329_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0064_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0792_  (.A(\INST_config_UART._0214_ ),
    .B(\INST_config_UART.GetWordState[2] ),
    .C(\INST_config_UART._0316_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0330_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0793_  (.A1(\INST_config_UART._0243_ ),
    .A2(\INST_config_UART.WriteData[17] ),
    .A3(\INST_config_UART._0236_ ),
    .B1(\INST_config_UART._0330_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0065_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0794_  (.A(\INST_config_UART._0214_ ),
    .B(\INST_config_UART.GetWordState[2] ),
    .C(\INST_config_UART._0318_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0331_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0795_  (.A1(\INST_config_UART._0243_ ),
    .A2(\INST_config_UART.WriteData[18] ),
    .A3(\INST_config_UART._0236_ ),
    .B1(\INST_config_UART._0331_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0066_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0796_  (.A(\INST_config_UART._0214_ ),
    .B(\INST_config_UART.GetWordState[2] ),
    .C(\INST_config_UART._0320_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0332_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0797_  (.A1(\INST_config_UART._0243_ ),
    .A2(\INST_config_UART.WriteData[19] ),
    .A3(\INST_config_UART._0236_ ),
    .B1(\INST_config_UART._0332_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0067_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0798_  (.A(\INST_config_UART._0214_ ),
    .B(\INST_config_UART.GetWordState[2] ),
    .C(\INST_config_UART._0322_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0333_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0799_  (.A1(\INST_config_UART._0243_ ),
    .A2(\INST_config_UART.WriteData[20] ),
    .A3(\INST_config_UART._0236_ ),
    .B1(\INST_config_UART._0333_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0068_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0800_  (.A(\INST_config_UART._0214_ ),
    .B(\INST_config_UART.GetWordState[2] ),
    .C(\INST_config_UART._0324_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0334_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0801_  (.A1(\INST_config_UART._0243_ ),
    .A2(\INST_config_UART.WriteData[21] ),
    .A3(\INST_config_UART._0236_ ),
    .B1(\INST_config_UART._0334_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0069_ ));
 sky130_fd_sc_hd__clkbuf_2 \INST_config_UART._0802_  (.A(\INST_config_UART.ByteWriteStrobe ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0335_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0803_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[2] ),
    .C(\INST_config_UART._0326_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0336_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0804_  (.A1(\INST_config_UART._0243_ ),
    .A2(\INST_config_UART.WriteData[22] ),
    .A3(\INST_config_UART._0236_ ),
    .B1(\INST_config_UART._0336_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0070_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0805_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[2] ),
    .C(\INST_config_UART._0328_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0337_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0806_  (.A1(\INST_config_UART._0243_ ),
    .A2(\INST_config_UART.WriteData[23] ),
    .A3(\INST_config_UART._0236_ ),
    .B1(\INST_config_UART._0337_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0071_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0807_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[1] ),
    .C(\INST_config_UART._0314_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0338_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0808_  (.A1(\INST_config_UART._0243_ ),
    .A2(\INST_config_UART.WriteData[8] ),
    .A3(\INST_config_UART._0215_ ),
    .B1(\INST_config_UART._0338_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0072_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._0809_  (.A(\INST_config_UART._0242_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0339_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0810_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[1] ),
    .C(\INST_config_UART._0316_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0340_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0811_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[9] ),
    .A3(\INST_config_UART._0215_ ),
    .B1(\INST_config_UART._0340_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0073_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0812_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[1] ),
    .C(\INST_config_UART._0318_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0341_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0813_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[10] ),
    .A3(\INST_config_UART._0215_ ),
    .B1(\INST_config_UART._0341_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0074_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0814_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[1] ),
    .C(\INST_config_UART._0320_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0342_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0815_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[11] ),
    .A3(\INST_config_UART._0215_ ),
    .B1(\INST_config_UART._0342_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0075_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0816_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[1] ),
    .C(\INST_config_UART._0322_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0343_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0817_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[12] ),
    .A3(\INST_config_UART._0215_ ),
    .B1(\INST_config_UART._0343_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0076_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0818_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[1] ),
    .C(\INST_config_UART._0324_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0344_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0819_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[13] ),
    .A3(\INST_config_UART._0215_ ),
    .B1(\INST_config_UART._0344_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0077_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0820_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[1] ),
    .C(\INST_config_UART._0326_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0345_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0821_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[14] ),
    .A3(\INST_config_UART._0215_ ),
    .B1(\INST_config_UART._0345_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0078_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0822_  (.A(\INST_config_UART._0335_ ),
    .B(\INST_config_UART.GetWordState[1] ),
    .C(\INST_config_UART._0328_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0346_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0823_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[15] ),
    .A3(\INST_config_UART._0215_ ),
    .B1(\INST_config_UART._0346_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0079_ ));
 sky130_fd_sc_hd__clkbuf_2 \INST_config_UART._0824_  (.A(\INST_config_UART.ComTick ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0347_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0825_  (.A0(\INST_config_UART._0250_ ),
    .A1(\INST_config_UART._0347_ ),
    .S(\INST_config_UART.ComState[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0348_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0826_  (.A(\INST_config_UART._0348_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0349_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._0827_  (.A(\INST_config_UART._0347_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0350_ ));
 sky130_fd_sc_hd__and3b_1 \INST_config_UART._0828_  (.A_N(\INST_config_UART._0251_ ),
    .B(\INST_config_UART._0350_ ),
    .C(\INST_config_UART.ComState[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0351_ ));
 sky130_fd_sc_hd__o22a_1 \INST_config_UART._0829_  (.A1(\INST_config_UART.RxLocal ),
    .A2(\INST_config_UART._0349_ ),
    .B1(\INST_config_UART._0351_ ),
    .B2(\INST_config_UART.ReceivedWord[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0080_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0830_  (.A0(\INST_config_UART._0250_ ),
    .A1(\INST_config_UART._0347_ ),
    .S(\INST_config_UART.ComState[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0352_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0831_  (.A(\INST_config_UART._0352_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0353_ ));
 sky130_fd_sc_hd__and3b_1 \INST_config_UART._0832_  (.A_N(\INST_config_UART._0250_ ),
    .B(\INST_config_UART._0347_ ),
    .C(\INST_config_UART.ComState[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0354_ ));
 sky130_fd_sc_hd__o22a_1 \INST_config_UART._0833_  (.A1(\INST_config_UART.RxLocal ),
    .A2(\INST_config_UART._0353_ ),
    .B1(\INST_config_UART._0354_ ),
    .B2(\INST_config_UART._0222_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0081_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0834_  (.A(\INST_config_UART.ComTick ),
    .B(\INST_config_UART.ComState[4] ),
    .C(\INST_config_UART.PresentState[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0355_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._0835_  (.A(\INST_config_UART._0355_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0356_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0836_  (.A0(\INST_config_UART.ID_Reg[16] ),
    .A1(\INST_config_UART._0223_ ),
    .S(\INST_config_UART._0356_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0357_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0837_  (.A(\INST_config_UART._0357_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0082_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0838_  (.A0(\INST_config_UART.ID_Reg[17] ),
    .A1(\INST_config_UART._0222_ ),
    .S(\INST_config_UART._0356_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0358_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0839_  (.A(\INST_config_UART._0358_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0083_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0840_  (.A0(\INST_config_UART.ID_Reg[18] ),
    .A1(\INST_config_UART._0221_ ),
    .S(\INST_config_UART._0356_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0359_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0841_  (.A(\INST_config_UART._0359_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0084_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0842_  (.A0(\INST_config_UART.ID_Reg[19] ),
    .A1(\INST_config_UART._0218_ ),
    .S(\INST_config_UART._0356_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0360_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0843_  (.A(\INST_config_UART._0360_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0085_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0844_  (.A0(\INST_config_UART.ID_Reg[20] ),
    .A1(\INST_config_UART.ReceivedWord[4] ),
    .S(\INST_config_UART._0356_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0361_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0845_  (.A(\INST_config_UART._0361_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0086_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0846_  (.A0(\INST_config_UART.ID_Reg[21] ),
    .A1(\INST_config_UART.ReceivedWord[5] ),
    .S(\INST_config_UART._0356_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0362_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0847_  (.A(\INST_config_UART._0362_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0087_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0848_  (.A0(\INST_config_UART.ID_Reg[22] ),
    .A1(\INST_config_UART.ReceivedWord[6] ),
    .S(\INST_config_UART._0356_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0363_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0849_  (.A(\INST_config_UART._0363_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0088_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0850_  (.A0(\INST_config_UART.ID_Reg[23] ),
    .A1(\INST_config_UART.ReceivedWord[7] ),
    .S(\INST_config_UART._0356_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0364_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0851_  (.A(\INST_config_UART._0364_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0089_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0852_  (.A0(\INST_config_UART._0250_ ),
    .A1(\INST_config_UART._0347_ ),
    .S(\INST_config_UART.ComState[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0365_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0853_  (.A(\INST_config_UART._0365_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0366_ ));
 sky130_fd_sc_hd__and3b_1 \INST_config_UART._0854_  (.A_N(\INST_config_UART._0250_ ),
    .B(\INST_config_UART._0347_ ),
    .C(\INST_config_UART.ComState[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0367_ ));
 sky130_fd_sc_hd__o22a_1 \INST_config_UART._0855_  (.A1(\INST_config_UART.RxLocal ),
    .A2(\INST_config_UART._0366_ ),
    .B1(\INST_config_UART._0367_ ),
    .B2(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0090_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0856_  (.A0(\INST_config_UART.ComState[0] ),
    .A1(\INST_config_UART._0347_ ),
    .S(\INST_config_UART.ComState[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0368_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0857_  (.A(\INST_config_UART._0368_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0369_ ));
 sky130_fd_sc_hd__and3b_1 \INST_config_UART._0858_  (.A_N(\INST_config_UART._0250_ ),
    .B(\INST_config_UART._0347_ ),
    .C(\INST_config_UART.ComState[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0370_ ));
 sky130_fd_sc_hd__o22a_1 \INST_config_UART._0859_  (.A1(\INST_config_UART.RxLocal ),
    .A2(\INST_config_UART._0369_ ),
    .B1(\INST_config_UART._0370_ ),
    .B2(\INST_config_UART.ReceivedWord[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0091_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0860_  (.A0(\INST_config_UART.ComState[0] ),
    .A1(\INST_config_UART.ComTick ),
    .S(\INST_config_UART.ComState[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0371_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0861_  (.A(\INST_config_UART._0371_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0372_ ));
 sky130_fd_sc_hd__and3b_1 \INST_config_UART._0862_  (.A_N(\INST_config_UART._0250_ ),
    .B(\INST_config_UART._0347_ ),
    .C(\INST_config_UART.ComState[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0373_ ));
 sky130_fd_sc_hd__o22a_1 \INST_config_UART._0863_  (.A1(\INST_config_UART.RxLocal ),
    .A2(\INST_config_UART._0372_ ),
    .B1(\INST_config_UART._0373_ ),
    .B2(\INST_config_UART._0223_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0092_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0864_  (.A(\INST_config_UART.ComTick ),
    .B(\INST_config_UART.ComState[4] ),
    .C(\INST_config_UART.PresentState[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0374_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._0865_  (.A(\INST_config_UART._0374_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0375_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0866_  (.A0(\INST_config_UART.ID_Reg[8] ),
    .A1(\INST_config_UART._0223_ ),
    .S(\INST_config_UART._0375_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0376_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0867_  (.A(\INST_config_UART._0376_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0093_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0868_  (.A0(\INST_config_UART.ID_Reg[9] ),
    .A1(\INST_config_UART._0222_ ),
    .S(\INST_config_UART._0375_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0377_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0869_  (.A(\INST_config_UART._0377_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0094_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0870_  (.A0(\INST_config_UART.ID_Reg[10] ),
    .A1(\INST_config_UART._0221_ ),
    .S(\INST_config_UART._0375_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0378_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0871_  (.A(\INST_config_UART._0378_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0095_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0872_  (.A0(\INST_config_UART.ID_Reg[11] ),
    .A1(\INST_config_UART._0218_ ),
    .S(\INST_config_UART._0375_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0379_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0873_  (.A(\INST_config_UART._0379_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0096_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0874_  (.A0(\INST_config_UART.ID_Reg[12] ),
    .A1(\INST_config_UART.ReceivedWord[4] ),
    .S(\INST_config_UART._0375_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0380_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0875_  (.A(\INST_config_UART._0380_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0097_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0876_  (.A0(\INST_config_UART.ID_Reg[13] ),
    .A1(\INST_config_UART.ReceivedWord[5] ),
    .S(\INST_config_UART._0375_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0381_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0877_  (.A(\INST_config_UART._0381_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0098_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0878_  (.A0(\INST_config_UART.ID_Reg[14] ),
    .A1(\INST_config_UART.ReceivedWord[6] ),
    .S(\INST_config_UART._0375_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0382_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0879_  (.A(\INST_config_UART._0382_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0099_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0880_  (.A0(\INST_config_UART.ID_Reg[15] ),
    .A1(\INST_config_UART.ReceivedWord[7] ),
    .S(\INST_config_UART._0375_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0383_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0881_  (.A(\INST_config_UART._0383_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0100_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0882_  (.A(\INST_config_UART.ReceivedWord[1] ),
    .B(\INST_config_UART.ReceivedWord[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0384_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0883_  (.A1(\INST_config_UART.ReceivedWord[3] ),
    .A2(\INST_config_UART._0384_ ),
    .B1(\INST_config_UART._0219_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0385_ ));
 sky130_fd_sc_hd__or4b_1 \INST_config_UART._0884_  (.A(\INST_config_UART.ReceivedWord[0] ),
    .B(\INST_config_UART.ReceivedWord[3] ),
    .C(\INST_config_UART._0225_ ),
    .D_N(\INST_config_UART._0384_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0386_ ));
 sky130_fd_sc_hd__a21bo_1 \INST_config_UART._0885_  (.A1(\INST_config_UART._0223_ ),
    .A2(\INST_config_UART._0385_ ),
    .B1_N(\INST_config_UART._0386_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0387_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0886_  (.A(\INST_config_UART.ReceiveState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0388_ ));
 sky130_fd_sc_hd__or2_2 \INST_config_UART._0887_  (.A(\INST_config_UART._0388_ ),
    .B(\INST_config_UART._0233_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0389_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0888_  (.A0(\INST_config_UART._0387_ ),
    .A1(\INST_config_UART.HighReg[0] ),
    .S(\INST_config_UART._0389_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0390_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0889_  (.A(\INST_config_UART._0390_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0101_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0890_  (.A(\INST_config_UART.ReceivedWord[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0391_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0891_  (.A(\INST_config_UART._0391_ ),
    .B(\INST_config_UART._0219_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0392_ ));
 sky130_fd_sc_hd__a21oi_2 \INST_config_UART._0892_  (.A1(\INST_config_UART._0227_ ),
    .A2(\INST_config_UART._0392_ ),
    .B1(\INST_config_UART._0218_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0393_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0893_  (.A0(\INST_config_UART._0393_ ),
    .A1(\INST_config_UART.HighReg[1] ),
    .S(\INST_config_UART._0389_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0394_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0894_  (.A(\INST_config_UART._0394_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0102_ ));
 sky130_fd_sc_hd__o21ai_2 \INST_config_UART._0895_  (.A1(\INST_config_UART._0219_ ),
    .A2(\INST_config_UART._0229_ ),
    .B1(\INST_config_UART._0231_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0395_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0896_  (.A0(\INST_config_UART._0395_ ),
    .A1(\INST_config_UART.HighReg[2] ),
    .S(\INST_config_UART._0389_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0396_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0897_  (.A(\INST_config_UART._0396_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0103_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0898_  (.A0(\INST_config_UART._0232_ ),
    .A1(\INST_config_UART.HighReg[3] ),
    .S(\INST_config_UART._0389_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0397_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0899_  (.A(\INST_config_UART._0397_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0104_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0900_  (.A(\INST_config_UART.ComState[4] ),
    .B(\INST_config_UART.PresentState[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0398_ ));
 sky130_fd_sc_hd__clkbuf_2 \INST_config_UART._0901_  (.A(\INST_config_UART._0398_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0399_ ));
 sky130_fd_sc_hd__or4_2 \INST_config_UART._0902_  (.A(\INST_config_UART.TimeToSendCounter[3] ),
    .B(\INST_config_UART.TimeToSendCounter[2] ),
    .C(\INST_config_UART.TimeToSendCounter[1] ),
    .D(\INST_config_UART.TimeToSendCounter[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0400_ ));
 sky130_fd_sc_hd__or4_2 \INST_config_UART._0903_  (.A(\INST_config_UART.TimeToSendCounter[6] ),
    .B(\INST_config_UART.TimeToSendCounter[5] ),
    .C(\INST_config_UART.TimeToSendCounter[4] ),
    .D(\INST_config_UART._0400_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0401_ ));
 sky130_fd_sc_hd__or3_2 \INST_config_UART._0904_  (.A(\INST_config_UART.TimeToSendCounter[8] ),
    .B(\INST_config_UART.TimeToSendCounter[7] ),
    .C(\INST_config_UART._0401_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0402_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0905_  (.A(\INST_config_UART.TimeToSendCounter[9] ),
    .B(\INST_config_UART._0402_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0403_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._0906_  (.A(\INST_config_UART.TimeToSendCounter[11] ),
    .B(\INST_config_UART.TimeToSendCounter[10] ),
    .C(\INST_config_UART._0403_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0404_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0907_  (.A(\INST_config_UART.TimeToSendCounter[12] ),
    .B(\INST_config_UART._0404_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0405_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._0908_  (.A(\INST_config_UART.TimeToSendCounter[13] ),
    .B(\INST_config_UART.TimeToSendCounter[14] ),
    .C(\INST_config_UART._0405_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0406_ ));
 sky130_fd_sc_hd__or2_2 \INST_config_UART._0909_  (.A(\INST_config_UART._0399_ ),
    .B(\INST_config_UART._0406_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0407_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0910_  (.A(\INST_config_UART._0407_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0408_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0911_  (.A0(\INST_config_UART.TimeToSend ),
    .A1(\INST_config_UART._0408_ ),
    .S(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0409_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0912_  (.A(\INST_config_UART._0409_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0105_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0913_  (.A0(\INST_config_UART.HexData[0] ),
    .A1(\INST_config_UART._0387_ ),
    .S(\INST_config_UART._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0410_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0914_  (.A(\INST_config_UART._0410_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0106_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0915_  (.A0(\INST_config_UART.HexData[1] ),
    .A1(\INST_config_UART._0393_ ),
    .S(\INST_config_UART._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0411_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0916_  (.A(\INST_config_UART._0411_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0107_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0917_  (.A0(\INST_config_UART.HexData[2] ),
    .A1(\INST_config_UART._0395_ ),
    .S(\INST_config_UART._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0412_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0918_  (.A(\INST_config_UART._0412_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0108_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0919_  (.A0(\INST_config_UART.HexData[3] ),
    .A1(\INST_config_UART._0232_ ),
    .S(\INST_config_UART._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0413_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0920_  (.A(\INST_config_UART._0413_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0109_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0921_  (.A0(\INST_config_UART.HexData[4] ),
    .A1(\INST_config_UART.HighReg[0] ),
    .S(\INST_config_UART._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0414_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0922_  (.A(\INST_config_UART._0414_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0110_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0923_  (.A0(\INST_config_UART.HexData[5] ),
    .A1(\INST_config_UART.HighReg[1] ),
    .S(\INST_config_UART._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0415_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0924_  (.A(\INST_config_UART._0415_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0111_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0925_  (.A0(\INST_config_UART.HexData[6] ),
    .A1(\INST_config_UART.HighReg[2] ),
    .S(\INST_config_UART._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0416_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0926_  (.A(\INST_config_UART._0416_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0112_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0927_  (.A0(\INST_config_UART.HexData[7] ),
    .A1(\INST_config_UART.HighReg[3] ),
    .S(\INST_config_UART._0014_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0417_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._0928_  (.A(\INST_config_UART._0417_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0113_ ));
 sky130_fd_sc_hd__or2b_1 \INST_config_UART._0929_  (.A(\INST_config_UART._0399_ ),
    .B_N(\INST_config_UART._0406_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0418_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._0930_  (.A(\INST_config_UART._0418_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0419_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0931_  (.A(\INST_config_UART.TimeToSendCounter[0] ),
    .B(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0114_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0932_  (.A(\INST_config_UART.TimeToSendCounter[1] ),
    .B(\INST_config_UART.TimeToSendCounter[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0420_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0933_  (.A(\INST_config_UART.TimeToSendCounter[1] ),
    .B(\INST_config_UART.TimeToSendCounter[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0421_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0934_  (.A1(\INST_config_UART._0420_ ),
    .A2(\INST_config_UART._0421_ ),
    .B1(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0115_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0935_  (.A(\INST_config_UART.TimeToSendCounter[2] ),
    .B(\INST_config_UART._0420_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0422_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0936_  (.A(\INST_config_UART.TimeToSendCounter[2] ),
    .B(\INST_config_UART._0420_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0423_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0937_  (.A1(\INST_config_UART._0422_ ),
    .A2(\INST_config_UART._0423_ ),
    .B1(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0116_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0938_  (.A(\INST_config_UART._0400_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0424_ ));
 sky130_fd_sc_hd__and2_1 \INST_config_UART._0939_  (.A(\INST_config_UART.TimeToSendCounter[3] ),
    .B(\INST_config_UART._0422_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0425_ ));
 sky130_fd_sc_hd__o31a_1 \INST_config_UART._0940_  (.A1(\INST_config_UART._0399_ ),
    .A2(\INST_config_UART._0424_ ),
    .A3(\INST_config_UART._0425_ ),
    .B1(\INST_config_UART._0407_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0117_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0941_  (.A(\INST_config_UART.TimeToSendCounter[4] ),
    .B(\INST_config_UART._0400_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0426_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0942_  (.A(\INST_config_UART.TimeToSendCounter[4] ),
    .B(\INST_config_UART._0400_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0427_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0943_  (.A1(\INST_config_UART._0426_ ),
    .A2(\INST_config_UART._0427_ ),
    .B1(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0118_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0944_  (.A(\INST_config_UART.TimeToSendCounter[5] ),
    .B(\INST_config_UART._0426_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0428_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0945_  (.A1(\INST_config_UART.TimeToSendCounter[4] ),
    .A2(\INST_config_UART._0400_ ),
    .B1(\INST_config_UART.TimeToSendCounter[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0429_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0946_  (.A1(\INST_config_UART._0428_ ),
    .A2(\INST_config_UART._0429_ ),
    .B1(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0119_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0947_  (.A(\INST_config_UART.TimeToSendCounter[6] ),
    .B(\INST_config_UART._0428_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0430_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0948_  (.A1(\INST_config_UART._0401_ ),
    .A2(\INST_config_UART._0430_ ),
    .B1(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0120_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0949_  (.A(\INST_config_UART.TimeToSendCounter[7] ),
    .B(\INST_config_UART._0401_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0431_ ));
 sky130_fd_sc_hd__and2_1 \INST_config_UART._0950_  (.A(\INST_config_UART.TimeToSendCounter[7] ),
    .B(\INST_config_UART._0401_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0432_ ));
 sky130_fd_sc_hd__o31a_1 \INST_config_UART._0951_  (.A1(\INST_config_UART._0399_ ),
    .A2(\INST_config_UART._0431_ ),
    .A3(\INST_config_UART._0432_ ),
    .B1(\INST_config_UART._0407_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0121_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0952_  (.A(\INST_config_UART._0402_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0433_ ));
 sky130_fd_sc_hd__o21a_1 \INST_config_UART._0953_  (.A1(\INST_config_UART.TimeToSendCounter[7] ),
    .A2(\INST_config_UART._0401_ ),
    .B1(\INST_config_UART.TimeToSendCounter[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0434_ ));
 sky130_fd_sc_hd__o31a_1 \INST_config_UART._0954_  (.A1(\INST_config_UART._0399_ ),
    .A2(\INST_config_UART._0433_ ),
    .A3(\INST_config_UART._0434_ ),
    .B1(\INST_config_UART._0407_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0122_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0955_  (.A(\INST_config_UART.TimeToSendCounter[9] ),
    .B(\INST_config_UART._0402_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0435_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0956_  (.A1(\INST_config_UART._0403_ ),
    .A2(\INST_config_UART._0435_ ),
    .B1(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0123_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0957_  (.A(\INST_config_UART.TimeToSendCounter[10] ),
    .B(\INST_config_UART._0403_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0436_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0958_  (.A(\INST_config_UART.TimeToSendCounter[10] ),
    .B(\INST_config_UART._0403_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0437_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0959_  (.A1(\INST_config_UART._0436_ ),
    .A2(\INST_config_UART._0437_ ),
    .B1(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0124_ ));
 sky130_fd_sc_hd__o21ai_1 \INST_config_UART._0960_  (.A1(\INST_config_UART.TimeToSendCounter[10] ),
    .A2(\INST_config_UART._0403_ ),
    .B1(\INST_config_UART.TimeToSendCounter[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0438_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0961_  (.A1(\INST_config_UART._0404_ ),
    .A2(\INST_config_UART._0438_ ),
    .B1(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0125_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0962_  (.A(\INST_config_UART.TimeToSendCounter[12] ),
    .B(\INST_config_UART._0404_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0439_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0963_  (.A1(\INST_config_UART._0405_ ),
    .A2(\INST_config_UART._0439_ ),
    .B1(\INST_config_UART._0419_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0126_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0964_  (.A(\INST_config_UART.TimeToSendCounter[13] ),
    .B(\INST_config_UART._0405_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0440_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0965_  (.A(\INST_config_UART.TimeToSendCounter[13] ),
    .B(\INST_config_UART._0405_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0441_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._0966_  (.A1(\INST_config_UART._0440_ ),
    .A2(\INST_config_UART._0441_ ),
    .B1(\INST_config_UART._0418_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0127_ ));
 sky130_fd_sc_hd__a21o_1 \INST_config_UART._0967_  (.A1(\INST_config_UART.TimeToSendCounter[14] ),
    .A2(\INST_config_UART._0440_ ),
    .B1(\INST_config_UART._0399_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0128_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0968_  (.A(\INST_config_UART.CRCReg[12] ),
    .B(\INST_config_UART.CRCReg[13] ),
    .C(\INST_config_UART.CRCReg[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0442_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0969_  (.A(\INST_config_UART.CRCReg[15] ),
    .B(\INST_config_UART._0442_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0443_ ));
 sky130_fd_sc_hd__or4_1 \INST_config_UART._0970_  (.A(\INST_config_UART.CRCReg[2] ),
    .B(\INST_config_UART.CRCReg[3] ),
    .C(\INST_config_UART.CRCReg[4] ),
    .D(\INST_config_UART.CRCReg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0444_ ));
 sky130_fd_sc_hd__and2_1 \INST_config_UART._0971_  (.A(\INST_config_UART.CRCReg[8] ),
    .B(\INST_config_UART.CRCReg[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0445_ ));
 sky130_fd_sc_hd__or4b_1 \INST_config_UART._0972_  (.A(\INST_config_UART.CRCReg[0] ),
    .B(\INST_config_UART.CRCReg[1] ),
    .C(\INST_config_UART._0444_ ),
    .D_N(\INST_config_UART._0445_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0446_ ));
 sky130_fd_sc_hd__or4b_1 \INST_config_UART._0973_  (.A(\INST_config_UART.CRCReg[6] ),
    .B(\INST_config_UART.CRCReg[7] ),
    .C(\INST_config_UART.CRCReg[10] ),
    .D_N(\INST_config_UART.CRCReg[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0447_ ));
 sky130_fd_sc_hd__or4b_1 \INST_config_UART._0974_  (.A(\INST_config_UART.CRCReg[16] ),
    .B(\INST_config_UART.CRCReg[17] ),
    .C(\INST_config_UART.CRCReg[19] ),
    .D_N(\INST_config_UART.CRCReg[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0448_ ));
 sky130_fd_sc_hd__or4_1 \INST_config_UART._0975_  (.A(\INST_config_UART._0443_ ),
    .B(\INST_config_UART._0446_ ),
    .C(\INST_config_UART._0447_ ),
    .D(\INST_config_UART._0448_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0449_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._0976_  (.A(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0450_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0977_  (.A1(\INST_config_UART.PresentState[0] ),
    .A2(\INST_config_UART.blink[22] ),
    .A3(\INST_config_UART._0449_ ),
    .B1(\INST_config_UART._0450_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0451_ ));
 sky130_fd_sc_hd__o22a_1 \INST_config_UART._0978_  (.A1(net111),
    .A2(\INST_config_UART.ReceiveLED ),
    .B1(\INST_config_UART._0451_ ),
    .B2(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0129_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0979_  (.A(\INST_config_UART._0216_ ),
    .B(\INST_config_UART.GetWordState[0] ),
    .C(\INST_config_UART._0314_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0452_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0980_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[24] ),
    .A3(\INST_config_UART._0234_ ),
    .B1(\INST_config_UART._0452_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0130_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0981_  (.A(\INST_config_UART._0216_ ),
    .B(\INST_config_UART.GetWordState[0] ),
    .C(\INST_config_UART._0316_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0453_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0982_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[25] ),
    .A3(\INST_config_UART._0234_ ),
    .B1(\INST_config_UART._0453_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0131_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0983_  (.A(\INST_config_UART._0216_ ),
    .B(\INST_config_UART.GetWordState[0] ),
    .C(\INST_config_UART._0318_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0454_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0984_  (.A1(\INST_config_UART._0339_ ),
    .A2(\INST_config_UART.WriteData[26] ),
    .A3(\INST_config_UART._0234_ ),
    .B1(\INST_config_UART._0454_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0132_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0985_  (.A(\INST_config_UART._0216_ ),
    .B(\INST_config_UART.GetWordState[0] ),
    .C(\INST_config_UART._0320_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0455_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0986_  (.A1(\INST_config_UART._0242_ ),
    .A2(\INST_config_UART.WriteData[27] ),
    .A3(\INST_config_UART._0234_ ),
    .B1(\INST_config_UART._0455_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0133_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0987_  (.A(\INST_config_UART._0216_ ),
    .B(\INST_config_UART.GetWordState[0] ),
    .C(\INST_config_UART._0322_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0456_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0988_  (.A1(\INST_config_UART._0242_ ),
    .A2(\INST_config_UART.WriteData[28] ),
    .A3(\INST_config_UART._0234_ ),
    .B1(\INST_config_UART._0456_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0134_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0989_  (.A(\INST_config_UART._0216_ ),
    .B(\INST_config_UART.GetWordState[0] ),
    .C(\INST_config_UART._0324_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0457_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0990_  (.A1(\INST_config_UART._0242_ ),
    .A2(\INST_config_UART.WriteData[29] ),
    .A3(\INST_config_UART._0234_ ),
    .B1(\INST_config_UART._0457_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0135_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0991_  (.A(\INST_config_UART._0216_ ),
    .B(\INST_config_UART.GetWordState[0] ),
    .C(\INST_config_UART._0326_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0458_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0992_  (.A1(\INST_config_UART._0242_ ),
    .A2(\INST_config_UART.WriteData[30] ),
    .A3(\INST_config_UART._0234_ ),
    .B1(\INST_config_UART._0458_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0136_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._0993_  (.A(\INST_config_UART._0216_ ),
    .B(\INST_config_UART.GetWordState[0] ),
    .C(\INST_config_UART._0328_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0459_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._0994_  (.A1(\INST_config_UART._0242_ ),
    .A2(\INST_config_UART.WriteData[31] ),
    .A3(\INST_config_UART._0234_ ),
    .B1(\INST_config_UART._0459_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0137_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._0995_  (.A0(\INST_config_UART._0223_ ),
    .A1(\INST_config_UART._0387_ ),
    .S(\INST_config_UART._0246_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0460_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._0996_  (.A(\INST_config_UART.CRCReg[0] ),
    .B(\INST_config_UART._0460_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0461_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._0997_  (.A(\INST_config_UART.CRCReg[0] ),
    .B(\INST_config_UART._0460_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0462_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._0998_  (.A(\INST_config_UART._0246_ ),
    .B(\INST_config_UART._0195_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0463_ ));
 sky130_fd_sc_hd__o21ai_2 \INST_config_UART._0999_  (.A1(\INST_config_UART._0014_ ),
    .A2(\INST_config_UART._0463_ ),
    .B1(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0464_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._1000_  (.A(\INST_config_UART._0192_ ),
    .B(\INST_config_UART._0464_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0465_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._1001_  (.A(\INST_config_UART._0465_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0466_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._1002_  (.A(\INST_config_UART._0464_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0467_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._1003_  (.A(\INST_config_UART._0192_ ),
    .B(\INST_config_UART._0467_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0468_ ));
 sky130_fd_sc_hd__buf_2 \INST_config_UART._1004_  (.A(\INST_config_UART._0468_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0469_ ));
 sky130_fd_sc_hd__a32o_1 \INST_config_UART._1005_  (.A1(\INST_config_UART._0461_ ),
    .A2(\INST_config_UART._0462_ ),
    .A3(\INST_config_UART._0466_ ),
    .B1(\INST_config_UART._0469_ ),
    .B2(\INST_config_UART.CRCReg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0138_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._1006_  (.A(\INST_config_UART._0222_ ),
    .B(\INST_config_UART._0246_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0470_ ));
 sky130_fd_sc_hd__o211ai_2 \INST_config_UART._1007_  (.A1(\INST_config_UART._0312_ ),
    .A2(\INST_config_UART._0393_ ),
    .B1(\INST_config_UART._0470_ ),
    .C1(\INST_config_UART.CRCReg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0471_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._1008_  (.A(\INST_config_UART._0391_ ),
    .B(\INST_config_UART._0246_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0472_ ));
 sky130_fd_sc_hd__a211o_1 \INST_config_UART._1009_  (.A1(\INST_config_UART._0246_ ),
    .A2(\INST_config_UART._0393_ ),
    .B1(\INST_config_UART._0472_ ),
    .C1(\INST_config_UART.CRCReg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0473_ ));
 sky130_fd_sc_hd__nand4_1 \INST_config_UART._1010_  (.A(\INST_config_UART.CRCReg[0] ),
    .B(\INST_config_UART._0460_ ),
    .C(\INST_config_UART._0471_ ),
    .D(\INST_config_UART._0473_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0474_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._1011_  (.A1(\INST_config_UART.CRCReg[0] ),
    .A2(\INST_config_UART._0460_ ),
    .B1(\INST_config_UART._0471_ ),
    .B2(\INST_config_UART._0473_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0475_ ));
 sky130_fd_sc_hd__a32o_1 \INST_config_UART._1012_  (.A1(\INST_config_UART._0466_ ),
    .A2(\INST_config_UART._0474_ ),
    .A3(\INST_config_UART._0475_ ),
    .B1(\INST_config_UART._0469_ ),
    .B2(\INST_config_UART.CRCReg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0139_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1013_  (.A0(\INST_config_UART._0221_ ),
    .A1(\INST_config_UART._0395_ ),
    .S(\INST_config_UART._0246_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0476_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._1014_  (.A(\INST_config_UART.CRCReg[2] ),
    .B(\INST_config_UART._0476_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0477_ ));
 sky130_fd_sc_hd__a21o_1 \INST_config_UART._1015_  (.A1(\INST_config_UART._0471_ ),
    .A2(\INST_config_UART._0474_ ),
    .B1(\INST_config_UART._0477_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0478_ ));
 sky130_fd_sc_hd__nand3_1 \INST_config_UART._1016_  (.A(\INST_config_UART._0471_ ),
    .B(\INST_config_UART._0474_ ),
    .C(\INST_config_UART._0477_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0479_ ));
 sky130_fd_sc_hd__a32o_1 \INST_config_UART._1017_  (.A1(\INST_config_UART._0466_ ),
    .A2(\INST_config_UART._0478_ ),
    .A3(\INST_config_UART._0479_ ),
    .B1(\INST_config_UART._0469_ ),
    .B2(\INST_config_UART.CRCReg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0140_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1018_  (.A0(\INST_config_UART._0218_ ),
    .A1(\INST_config_UART._0232_ ),
    .S(\INST_config_UART._0246_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0480_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._1019_  (.A(\INST_config_UART.CRCReg[3] ),
    .B(\INST_config_UART._0480_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0481_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1020_  (.A(\INST_config_UART.CRCReg[3] ),
    .B(\INST_config_UART._0480_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0482_ ));
 sky130_fd_sc_hd__or2b_1 \INST_config_UART._1021_  (.A(\INST_config_UART._0481_ ),
    .B_N(\INST_config_UART._0482_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0483_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1022_  (.A(\INST_config_UART.CRCReg[2] ),
    .B(\INST_config_UART._0476_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0484_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1023_  (.A(\INST_config_UART._0484_ ),
    .B(\INST_config_UART._0478_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0485_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._1024_  (.A(\INST_config_UART._0483_ ),
    .B(\INST_config_UART._0485_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0486_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._1025_  (.A1(\INST_config_UART.CRCReg[3] ),
    .A2(\INST_config_UART._0469_ ),
    .B1(\INST_config_UART._0466_ ),
    .B2(\INST_config_UART._0486_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0141_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._1026_  (.A1(\INST_config_UART._0484_ ),
    .A2(\INST_config_UART._0478_ ),
    .A3(\INST_config_UART._0482_ ),
    .B1(\INST_config_UART._0481_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0487_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1027_  (.A0(\INST_config_UART.ReceivedWord[4] ),
    .A1(\INST_config_UART.HighReg[0] ),
    .S(\INST_config_UART.Command[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0488_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._1028_  (.A(\INST_config_UART.CRCReg[4] ),
    .B(\INST_config_UART._0488_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0489_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1029_  (.A(\INST_config_UART.CRCReg[4] ),
    .B(\INST_config_UART._0488_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0490_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1030_  (.A(\INST_config_UART._0489_ ),
    .B(\INST_config_UART._0490_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0491_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1031_  (.A(\INST_config_UART._0487_ ),
    .B(\INST_config_UART._0491_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0492_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._1032_  (.A(\INST_config_UART._0487_ ),
    .B(\INST_config_UART._0491_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0493_ ));
 sky130_fd_sc_hd__a32o_1 \INST_config_UART._1033_  (.A1(\INST_config_UART._0466_ ),
    .A2(\INST_config_UART._0492_ ),
    .A3(\INST_config_UART._0493_ ),
    .B1(\INST_config_UART._0469_ ),
    .B2(\INST_config_UART.CRCReg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0142_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1034_  (.A0(\INST_config_UART.ReceivedWord[5] ),
    .A1(\INST_config_UART.HighReg[1] ),
    .S(\INST_config_UART.Command[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0494_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._1035_  (.A(\INST_config_UART.CRCReg[5] ),
    .B(\INST_config_UART._0494_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0495_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._1036_  (.A1(\INST_config_UART._0490_ ),
    .A2(\INST_config_UART._0493_ ),
    .B1(\INST_config_UART._0495_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0496_ ));
 sky130_fd_sc_hd__or2_2 \INST_config_UART._1037_  (.A(\INST_config_UART._0192_ ),
    .B(\INST_config_UART._0464_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0497_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._1038_  (.A1(\INST_config_UART._0490_ ),
    .A2(\INST_config_UART._0493_ ),
    .A3(\INST_config_UART._0495_ ),
    .B1(\INST_config_UART._0497_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0498_ ));
 sky130_fd_sc_hd__a2bb2o_1 \INST_config_UART._1039_  (.A1_N(\INST_config_UART._0496_ ),
    .A2_N(\INST_config_UART._0498_ ),
    .B1(\INST_config_UART.CRCReg[5] ),
    .B2(\INST_config_UART._0469_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0143_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1040_  (.A0(\INST_config_UART.ReceivedWord[6] ),
    .A1(\INST_config_UART.HighReg[2] ),
    .S(\INST_config_UART.Command[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0499_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._1041_  (.A(\INST_config_UART.CRCReg[6] ),
    .B(\INST_config_UART._0499_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0500_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1042_  (.A(\INST_config_UART.CRCReg[6] ),
    .B(\INST_config_UART._0499_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0501_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1043_  (.A(\INST_config_UART._0500_ ),
    .B(\INST_config_UART._0501_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0502_ ));
 sky130_fd_sc_hd__o211a_1 \INST_config_UART._1044_  (.A1(\INST_config_UART.CRCReg[5] ),
    .A2(\INST_config_UART._0494_ ),
    .B1(\INST_config_UART._0488_ ),
    .C1(\INST_config_UART.CRCReg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0503_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._1045_  (.A1(\INST_config_UART.CRCReg[5] ),
    .A2(\INST_config_UART._0494_ ),
    .B1(\INST_config_UART._0503_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0504_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._1046_  (.A(\INST_config_UART._0491_ ),
    .B(\INST_config_UART._0495_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0505_ ));
 sky130_fd_sc_hd__a311o_1 \INST_config_UART._1047_  (.A1(\INST_config_UART._0484_ ),
    .A2(\INST_config_UART._0478_ ),
    .A3(\INST_config_UART._0482_ ),
    .B1(\INST_config_UART._0505_ ),
    .C1(\INST_config_UART._0481_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0506_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1048_  (.A(\INST_config_UART._0504_ ),
    .B(\INST_config_UART._0506_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0507_ ));
 sky130_fd_sc_hd__xnor2_1 \INST_config_UART._1049_  (.A(\INST_config_UART._0502_ ),
    .B(\INST_config_UART._0507_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0508_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._1050_  (.A1(\INST_config_UART.CRCReg[6] ),
    .A2(\INST_config_UART._0469_ ),
    .B1(\INST_config_UART._0466_ ),
    .B2(\INST_config_UART._0508_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0144_ ));
 sky130_fd_sc_hd__a21o_1 \INST_config_UART._1051_  (.A1(\INST_config_UART._0504_ ),
    .A2(\INST_config_UART._0506_ ),
    .B1(\INST_config_UART._0502_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0509_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1052_  (.A0(\INST_config_UART.ReceivedWord[7] ),
    .A1(\INST_config_UART.HighReg[3] ),
    .S(\INST_config_UART._0246_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0510_ ));
 sky130_fd_sc_hd__nor2_1 \INST_config_UART._1053_  (.A(\INST_config_UART.CRCReg[7] ),
    .B(\INST_config_UART._0510_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0511_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1054_  (.A(\INST_config_UART.CRCReg[7] ),
    .B(\INST_config_UART._0510_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0512_ ));
 sky130_fd_sc_hd__or2b_1 \INST_config_UART._1055_  (.A(\INST_config_UART._0511_ ),
    .B_N(\INST_config_UART._0512_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0513_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._1056_  (.A1(\INST_config_UART._0501_ ),
    .A2(\INST_config_UART._0509_ ),
    .B1(\INST_config_UART._0513_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0514_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._1057_  (.A1(\INST_config_UART._0501_ ),
    .A2(\INST_config_UART._0509_ ),
    .A3(\INST_config_UART._0513_ ),
    .B1(\INST_config_UART._0497_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0515_ ));
 sky130_fd_sc_hd__a2bb2o_1 \INST_config_UART._1058_  (.A1_N(\INST_config_UART._0514_ ),
    .A2_N(\INST_config_UART._0515_ ),
    .B1(\INST_config_UART.CRCReg[7] ),
    .B2(\INST_config_UART._0469_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0145_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._1059_  (.A(\INST_config_UART._0502_ ),
    .B(\INST_config_UART._0505_ ),
    .C(\INST_config_UART._0513_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0516_ ));
 sky130_fd_sc_hd__a311o_2 \INST_config_UART._1060_  (.A1(\INST_config_UART._0484_ ),
    .A2(\INST_config_UART._0478_ ),
    .A3(\INST_config_UART._0482_ ),
    .B1(\INST_config_UART._0516_ ),
    .C1(\INST_config_UART._0481_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0517_ ));
 sky130_fd_sc_hd__or3_1 \INST_config_UART._1061_  (.A(\INST_config_UART._0502_ ),
    .B(\INST_config_UART._0504_ ),
    .C(\INST_config_UART._0513_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0518_ ));
 sky130_fd_sc_hd__o211a_2 \INST_config_UART._1062_  (.A1(\INST_config_UART._0501_ ),
    .A2(\INST_config_UART._0511_ ),
    .B1(\INST_config_UART._0512_ ),
    .C1(\INST_config_UART._0518_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0519_ ));
 sky130_fd_sc_hd__nand2_2 \INST_config_UART._1063_  (.A(\INST_config_UART._0517_ ),
    .B(\INST_config_UART._0519_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0520_ ));
 sky130_fd_sc_hd__or2_1 \INST_config_UART._1064_  (.A(\INST_config_UART.CRCReg[8] ),
    .B(\INST_config_UART._0520_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0521_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1065_  (.A(\INST_config_UART.CRCReg[8] ),
    .B(\INST_config_UART._0520_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0522_ ));
 sky130_fd_sc_hd__a32o_1 \INST_config_UART._1066_  (.A1(\INST_config_UART._0466_ ),
    .A2(\INST_config_UART._0521_ ),
    .A3(\INST_config_UART._0522_ ),
    .B1(\INST_config_UART._0469_ ),
    .B2(\INST_config_UART.CRCReg[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0146_ ));
 sky130_fd_sc_hd__a21o_1 \INST_config_UART._1067_  (.A1(\INST_config_UART.CRCReg[8] ),
    .A2(\INST_config_UART._0520_ ),
    .B1(\INST_config_UART.CRCReg[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0523_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1068_  (.A(\INST_config_UART._0445_ ),
    .B(\INST_config_UART._0520_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0524_ ));
 sky130_fd_sc_hd__a32o_1 \INST_config_UART._1069_  (.A1(\INST_config_UART._0466_ ),
    .A2(\INST_config_UART._0523_ ),
    .A3(\INST_config_UART._0524_ ),
    .B1(\INST_config_UART._0468_ ),
    .B2(\INST_config_UART.CRCReg[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0147_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._1070_  (.A1(\INST_config_UART._0445_ ),
    .A2(\INST_config_UART._0520_ ),
    .B1(\INST_config_UART.CRCReg[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0525_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._1071_  (.A(\INST_config_UART.CRCReg[10] ),
    .B(\INST_config_UART._0445_ ),
    .C(\INST_config_UART._0520_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0526_ ));
 sky130_fd_sc_hd__nand2_1 \INST_config_UART._1072_  (.A(\INST_config_UART.CRCReg[10] ),
    .B(\INST_config_UART._0468_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0527_ ));
 sky130_fd_sc_hd__o31ai_1 \INST_config_UART._1073_  (.A1(\INST_config_UART._0497_ ),
    .A2(\INST_config_UART._0525_ ),
    .A3(\INST_config_UART._0526_ ),
    .B1(\INST_config_UART._0527_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0148_ ));
 sky130_fd_sc_hd__nand3_2 \INST_config_UART._1074_  (.A(\INST_config_UART.CRCReg[10] ),
    .B(\INST_config_UART.CRCReg[11] ),
    .C(\INST_config_UART._0445_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0528_ ));
 sky130_fd_sc_hd__a21oi_4 \INST_config_UART._1075_  (.A1(\INST_config_UART._0517_ ),
    .A2(\INST_config_UART._0519_ ),
    .B1(\INST_config_UART._0528_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0529_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._1076_  (.A(\INST_config_UART._0529_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0530_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._1077_  (.A1(\INST_config_UART._0467_ ),
    .A2(\INST_config_UART._0529_ ),
    .B1(\INST_config_UART._0192_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0531_ ));
 sky130_fd_sc_hd__a32o_1 \INST_config_UART._1078_  (.A1(\INST_config_UART._0466_ ),
    .A2(\INST_config_UART._0526_ ),
    .A3(\INST_config_UART._0530_ ),
    .B1(\INST_config_UART._0531_ ),
    .B2(\INST_config_UART.CRCReg[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0149_ ));
 sky130_fd_sc_hd__a21oi_1 \INST_config_UART._1079_  (.A1(\INST_config_UART.CRCReg[12] ),
    .A2(\INST_config_UART._0529_ ),
    .B1(\INST_config_UART._0497_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0532_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._1080_  (.A1(\INST_config_UART.CRCReg[12] ),
    .A2(\INST_config_UART._0531_ ),
    .B1(\INST_config_UART._0532_ ),
    .B2(\INST_config_UART._0529_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0150_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._1081_  (.A(\INST_config_UART.CRCReg[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0533_ ));
 sky130_fd_sc_hd__a31o_1 \INST_config_UART._1082_  (.A1(\INST_config_UART.CRCReg[12] ),
    .A2(\INST_config_UART._0466_ ),
    .A3(\INST_config_UART._0529_ ),
    .B1(\INST_config_UART.CRCReg[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0534_ ));
 sky130_fd_sc_hd__o31a_1 \INST_config_UART._1083_  (.A1(\INST_config_UART._0533_ ),
    .A2(\INST_config_UART._0468_ ),
    .A3(\INST_config_UART._0532_ ),
    .B1(\INST_config_UART._0534_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0151_ ));
 sky130_fd_sc_hd__a31oi_1 \INST_config_UART._1084_  (.A1(\INST_config_UART._0442_ ),
    .A2(\INST_config_UART._0467_ ),
    .A3(\INST_config_UART._0529_ ),
    .B1(\INST_config_UART._0192_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0535_ ));
 sky130_fd_sc_hd__and4b_1 \INST_config_UART._1085_  (.A_N(\INST_config_UART._0442_ ),
    .B(\INST_config_UART._0465_ ),
    .C(\INST_config_UART._0529_ ),
    .D(\INST_config_UART.CRCReg[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0536_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._1086_  (.A1(\INST_config_UART.CRCReg[14] ),
    .A2(\INST_config_UART._0535_ ),
    .B1(\INST_config_UART._0536_ ),
    .B2(\INST_config_UART.CRCReg[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0152_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._1087_  (.A(\INST_config_UART._0442_ ),
    .B(\INST_config_UART._0465_ ),
    .C(\INST_config_UART._0529_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0537_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1088_  (.A0(\INST_config_UART._0537_ ),
    .A1(\INST_config_UART._0535_ ),
    .S(\INST_config_UART.CRCReg[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0538_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1089_  (.A(\INST_config_UART._0538_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0153_ ));
 sky130_fd_sc_hd__a211oi_4 \INST_config_UART._1090_  (.A1(\INST_config_UART._0517_ ),
    .A2(\INST_config_UART._0519_ ),
    .B1(\INST_config_UART._0528_ ),
    .C1(\INST_config_UART._0443_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0539_ ));
 sky130_fd_sc_hd__a31oi_2 \INST_config_UART._1091_  (.A1(\INST_config_UART.CRCReg[16] ),
    .A2(\INST_config_UART._0467_ ),
    .A3(\INST_config_UART._0539_ ),
    .B1(\INST_config_UART._0192_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0540_ ));
 sky130_fd_sc_hd__and3b_1 \INST_config_UART._1092_  (.A_N(\INST_config_UART.CRCReg[16] ),
    .B(\INST_config_UART._0465_ ),
    .C(\INST_config_UART._0539_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0541_ ));
 sky130_fd_sc_hd__a21o_1 \INST_config_UART._1093_  (.A1(\INST_config_UART.CRCReg[16] ),
    .A2(\INST_config_UART._0540_ ),
    .B1(\INST_config_UART._0541_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0154_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._1094_  (.A(\INST_config_UART.CRCReg[16] ),
    .B(\INST_config_UART._0465_ ),
    .C(\INST_config_UART._0539_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0542_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1095_  (.A0(\INST_config_UART._0542_ ),
    .A1(\INST_config_UART._0540_ ),
    .S(\INST_config_UART.CRCReg[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0543_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1096_  (.A(\INST_config_UART._0543_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0155_ ));
 sky130_fd_sc_hd__and2_1 \INST_config_UART._1097_  (.A(\INST_config_UART.CRCReg[16] ),
    .B(\INST_config_UART.CRCReg[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0544_ ));
 sky130_fd_sc_hd__a31oi_1 \INST_config_UART._1098_  (.A1(\INST_config_UART.CRCReg[18] ),
    .A2(\INST_config_UART._0539_ ),
    .A3(\INST_config_UART._0544_ ),
    .B1(\INST_config_UART._0497_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0545_ ));
 sky130_fd_sc_hd__a21o_1 \INST_config_UART._1099_  (.A1(\INST_config_UART._0539_ ),
    .A2(\INST_config_UART._0544_ ),
    .B1(\INST_config_UART.CRCReg[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0546_ ));
 sky130_fd_sc_hd__a22o_1 \INST_config_UART._1100_  (.A1(\INST_config_UART.CRCReg[18] ),
    .A2(\INST_config_UART._0469_ ),
    .B1(\INST_config_UART._0545_ ),
    .B2(\INST_config_UART._0546_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0156_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._1101_  (.A(\INST_config_UART.CRCReg[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0547_ ));
 sky130_fd_sc_hd__a41o_1 \INST_config_UART._1102_  (.A1(\INST_config_UART.CRCReg[18] ),
    .A2(\INST_config_UART._0465_ ),
    .A3(\INST_config_UART._0539_ ),
    .A4(\INST_config_UART._0544_ ),
    .B1(\INST_config_UART.CRCReg[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0548_ ));
 sky130_fd_sc_hd__o31a_1 \INST_config_UART._1103_  (.A1(\INST_config_UART._0547_ ),
    .A2(\INST_config_UART._0468_ ),
    .A3(\INST_config_UART._0545_ ),
    .B1(\INST_config_UART._0548_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0157_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1104_  (.A0(\INST_config_UART.ComState[0] ),
    .A1(\INST_config_UART.ComTick ),
    .S(\INST_config_UART.ComState[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0549_ ));
 sky130_fd_sc_hd__inv_2 \INST_config_UART._1105_  (.A(\INST_config_UART._0549_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\INST_config_UART._0550_ ));
 sky130_fd_sc_hd__and3b_1 \INST_config_UART._1106_  (.A_N(\INST_config_UART._0250_ ),
    .B(\INST_config_UART._0347_ ),
    .C(\INST_config_UART.ComState[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0551_ ));
 sky130_fd_sc_hd__o22a_1 \INST_config_UART._1107_  (.A1(\INST_config_UART.RxLocal ),
    .A2(\INST_config_UART._0550_ ),
    .B1(\INST_config_UART._0551_ ),
    .B2(\INST_config_UART.ReceivedWord[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0158_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._1108_  (.A(\INST_config_UART.ComTick ),
    .B(\INST_config_UART.ComState[4] ),
    .C(\INST_config_UART.PresentState[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0552_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._1109_  (.A(\INST_config_UART._0552_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0553_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1110_  (.A0(\INST_config_UART.ID_Reg[0] ),
    .A1(\INST_config_UART._0223_ ),
    .S(\INST_config_UART._0553_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0554_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1111_  (.A(\INST_config_UART._0554_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0159_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1112_  (.A0(\INST_config_UART.ID_Reg[1] ),
    .A1(\INST_config_UART._0222_ ),
    .S(\INST_config_UART._0553_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0555_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1113_  (.A(\INST_config_UART._0555_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0160_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1114_  (.A0(\INST_config_UART.ID_Reg[2] ),
    .A1(\INST_config_UART._0221_ ),
    .S(\INST_config_UART._0553_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0556_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1115_  (.A(\INST_config_UART._0556_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0161_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1116_  (.A0(\INST_config_UART.ID_Reg[3] ),
    .A1(\INST_config_UART._0218_ ),
    .S(\INST_config_UART._0553_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0557_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1117_  (.A(\INST_config_UART._0557_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0162_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1118_  (.A0(\INST_config_UART.ID_Reg[4] ),
    .A1(\INST_config_UART.ReceivedWord[4] ),
    .S(\INST_config_UART._0553_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0558_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1119_  (.A(\INST_config_UART._0558_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0163_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1120_  (.A0(\INST_config_UART.ID_Reg[5] ),
    .A1(\INST_config_UART.ReceivedWord[5] ),
    .S(\INST_config_UART._0553_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0559_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1121_  (.A(\INST_config_UART._0559_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0164_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1122_  (.A0(\INST_config_UART.ID_Reg[6] ),
    .A1(\INST_config_UART.ReceivedWord[6] ),
    .S(\INST_config_UART._0553_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0560_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1123_  (.A(\INST_config_UART._0560_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0165_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1124_  (.A0(\INST_config_UART.ID_Reg[7] ),
    .A1(\INST_config_UART.ReceivedWord[7] ),
    .S(\INST_config_UART._0553_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0561_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1125_  (.A(\INST_config_UART._0561_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0166_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._1126_  (.A(\INST_config_UART.ComTick ),
    .B(\INST_config_UART.ComState[4] ),
    .C(\INST_config_UART.PresentState[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0562_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._1127_  (.A(\INST_config_UART._0562_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0563_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1128_  (.A0(\INST_config_UART.Command[0] ),
    .A1(\INST_config_UART._0223_ ),
    .S(\INST_config_UART._0563_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0564_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1129_  (.A(\INST_config_UART._0564_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0167_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1130_  (.A0(\INST_config_UART.Command[1] ),
    .A1(\INST_config_UART._0222_ ),
    .S(\INST_config_UART._0563_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0565_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1131_  (.A(\INST_config_UART._0565_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0168_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1132_  (.A0(\INST_config_UART.Command[2] ),
    .A1(\INST_config_UART._0221_ ),
    .S(\INST_config_UART._0563_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0566_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1133_  (.A(\INST_config_UART._0566_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0169_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1134_  (.A0(\INST_config_UART.Command[3] ),
    .A1(\INST_config_UART._0218_ ),
    .S(\INST_config_UART._0563_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0567_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1135_  (.A(\INST_config_UART._0567_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0170_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1136_  (.A0(\INST_config_UART.Command[4] ),
    .A1(\INST_config_UART.ReceivedWord[4] ),
    .S(\INST_config_UART._0563_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0568_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1137_  (.A(\INST_config_UART._0568_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0171_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1138_  (.A0(\INST_config_UART.Command[5] ),
    .A1(\INST_config_UART.ReceivedWord[5] ),
    .S(\INST_config_UART._0563_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0569_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1139_  (.A(\INST_config_UART._0569_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0172_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1140_  (.A0(\INST_config_UART.Command[6] ),
    .A1(\INST_config_UART.ReceivedWord[6] ),
    .S(\INST_config_UART._0563_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0570_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1141_  (.A(\INST_config_UART._0570_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0173_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1142_  (.A0(\INST_config_UART._0247_ ),
    .A1(\INST_config_UART.ReceivedWord[7] ),
    .S(\INST_config_UART._0563_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0571_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1143_  (.A(\INST_config_UART._0571_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0174_ ));
 sky130_fd_sc_hd__and3_1 \INST_config_UART._1144_  (.A(net39),
    .B(net112),
    .C(\INST_config_UART._0193_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0572_ ));
 sky130_fd_sc_hd__clkbuf_4 \INST_config_UART._1145_  (.A(\INST_config_UART._0572_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0573_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1146_  (.A0(\INST_config_UART.Data_Reg[0] ),
    .A1(\INST_config_UART._0223_ ),
    .S(\INST_config_UART._0573_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0574_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1147_  (.A(\INST_config_UART._0574_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0175_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1148_  (.A0(\INST_config_UART.Data_Reg[1] ),
    .A1(\INST_config_UART._0222_ ),
    .S(\INST_config_UART._0573_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0575_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1149_  (.A(\INST_config_UART._0575_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0176_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1150_  (.A0(\INST_config_UART.Data_Reg[2] ),
    .A1(\INST_config_UART._0221_ ),
    .S(\INST_config_UART._0573_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0576_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1151_  (.A(\INST_config_UART._0576_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0177_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1152_  (.A0(\INST_config_UART.Data_Reg[3] ),
    .A1(\INST_config_UART._0218_ ),
    .S(\INST_config_UART._0573_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0577_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1153_  (.A(\INST_config_UART._0577_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0178_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1154_  (.A0(\INST_config_UART.Data_Reg[4] ),
    .A1(\INST_config_UART.ReceivedWord[4] ),
    .S(\INST_config_UART._0573_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0578_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1155_  (.A(\INST_config_UART._0578_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0179_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1156_  (.A0(\INST_config_UART.Data_Reg[5] ),
    .A1(\INST_config_UART.ReceivedWord[5] ),
    .S(\INST_config_UART._0573_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0579_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1157_  (.A(\INST_config_UART._0579_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0180_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1158_  (.A0(\INST_config_UART.Data_Reg[6] ),
    .A1(\INST_config_UART.ReceivedWord[6] ),
    .S(\INST_config_UART._0573_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0580_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1159_  (.A(\INST_config_UART._0580_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0181_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1160_  (.A0(\INST_config_UART.Data_Reg[7] ),
    .A1(\INST_config_UART.ReceivedWord[7] ),
    .S(\INST_config_UART._0573_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0581_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1161_  (.A(\INST_config_UART._0581_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0182_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1162_  (.A0(\INST_config_UART.ComState[10] ),
    .A1(\INST_config_UART.ComState[5] ),
    .S(\INST_config_UART._0350_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0582_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1163_  (.A(\INST_config_UART._0582_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0183_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1164_  (.A0(\INST_config_UART.ComState[9] ),
    .A1(\INST_config_UART.ComState[3] ),
    .S(\INST_config_UART._0350_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0583_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1165_  (.A(\INST_config_UART._0583_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0184_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1166_  (.A0(\INST_config_UART.ComState[8] ),
    .A1(\INST_config_UART.ComState[2] ),
    .S(\INST_config_UART._0350_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0584_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1167_  (.A(\INST_config_UART._0584_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0185_ ));
 sky130_fd_sc_hd__a21bo_1 \INST_config_UART._1168_  (.A1(\INST_config_UART._0350_ ),
    .A2(\INST_config_UART.ComState[1] ),
    .B1_N(\INST_config_UART._0306_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0186_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1169_  (.A0(\INST_config_UART.ComState[5] ),
    .A1(\INST_config_UART.ComState[8] ),
    .S(\INST_config_UART._0350_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0585_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1170_  (.A(\INST_config_UART._0585_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0187_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1171_  (.A0(\INST_config_UART.ComState[4] ),
    .A1(\INST_config_UART.ComState[7] ),
    .S(\INST_config_UART._0350_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0586_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1172_  (.A(\INST_config_UART._0586_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0188_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1173_  (.A0(\INST_config_UART.ComState[3] ),
    .A1(\INST_config_UART.ComState[6] ),
    .S(\INST_config_UART._0350_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0587_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1174_  (.A(\INST_config_UART._0587_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0189_ ));
 sky130_fd_sc_hd__a21bo_1 \INST_config_UART._1175_  (.A1(\INST_config_UART._0350_ ),
    .A2(\INST_config_UART.ComState[9] ),
    .B1_N(\INST_config_UART._0309_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0190_ ));
 sky130_fd_sc_hd__mux2_1 \INST_config_UART._1176_  (.A0(\INST_config_UART.ComState[1] ),
    .A1(\INST_config_UART.ComState[10] ),
    .S(\INST_config_UART._0350_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0588_ ));
 sky130_fd_sc_hd__clkbuf_1 \INST_config_UART._1177_  (.A(\INST_config_UART._0588_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\INST_config_UART._0191_ ));
 sky130_fd_sc_hd__dfrtp_4 \INST_config_UART._1178_  (.CLK(net1),
    .D(\INST_config_UART._0054_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceivedWord[7] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1179_  (.CLK(net1),
    .D(\INST_config_UART._0025_ ),
    .SET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.PresentState[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1180_  (.CLK(net1),
    .D(\INST_config_UART._0026_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.PresentState[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1181_  (.CLK(net1),
    .D(\INST_config_UART._0027_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.PresentState[2] ));
 sky130_fd_sc_hd__dfrtp_4 \INST_config_UART._1182_  (.CLK(net1),
    .D(\INST_config_UART._0028_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1183_  (.CLK(net1),
    .D(\INST_config_UART._0029_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.PresentState[4] ));
 sky130_fd_sc_hd__dfrtp_4 \INST_config_UART._1184_  (.CLK(net1),
    .D(\INST_config_UART._0018_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.PresentState[5] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1185_  (.CLK(net1),
    .D(\INST_config_UART._0030_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.PresentState[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1186_  (.CLK(net1),
    .D(\INST_config_UART._0055_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceivedWord[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1187_  (.CLK(net1),
    .D(\INST_config_UART._0056_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1188_  (.CLK(net1),
    .D(\INST_config_UART._0057_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1189_  (.CLK(net1),
    .D(\INST_config_UART._0058_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1190_  (.CLK(net1),
    .D(\INST_config_UART._0059_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1191_  (.CLK(net1),
    .D(\INST_config_UART._0060_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1192_  (.CLK(net1),
    .D(\INST_config_UART._0061_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[5] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1193_  (.CLK(net1),
    .D(\INST_config_UART._0062_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1194_  (.CLK(net1),
    .D(\INST_config_UART._0063_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[7] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1195_  (.CLK(net1),
    .D(\INST_config_UART._0064_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[16] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1196_  (.CLK(net1),
    .D(\INST_config_UART._0065_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[17] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1197_  (.CLK(net1),
    .D(\INST_config_UART._0066_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[18] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1198_  (.CLK(net1),
    .D(\INST_config_UART._0067_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[19] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1199_  (.CLK(net1),
    .D(\INST_config_UART._0068_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[20] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1200_  (.CLK(net1),
    .D(\INST_config_UART._0069_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[21] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1201_  (.CLK(net1),
    .D(\INST_config_UART._0070_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[22] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1202_  (.CLK(net1),
    .D(\INST_config_UART._0071_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[23] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1203_  (.CLK(net1),
    .D(\INST_config_UART._0072_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[8] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1204_  (.CLK(net1),
    .D(\INST_config_UART._0073_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[9] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1205_  (.CLK(net1),
    .D(\INST_config_UART._0074_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[10] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1206_  (.CLK(net1),
    .D(\INST_config_UART._0075_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[11] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1207_  (.CLK(net1),
    .D(\INST_config_UART._0076_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[12] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1208_  (.CLK(net1),
    .D(\INST_config_UART._0077_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[13] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1209_  (.CLK(net1),
    .D(\INST_config_UART._0078_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[14] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1210_  (.CLK(net1),
    .D(\INST_config_UART._0079_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[15] ));
 sky130_fd_sc_hd__dfstp_2 \INST_config_UART._1211_  (.CLK(net1),
    .D(\INST_config_UART._0021_ ),
    .SET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.GetWordState[0] ));
 sky130_fd_sc_hd__dfrtp_4 \INST_config_UART._1212_  (.CLK(net1),
    .D(\INST_config_UART._0022_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.GetWordState[1] ));
 sky130_fd_sc_hd__dfrtp_4 \INST_config_UART._1213_  (.CLK(net1),
    .D(\INST_config_UART._0023_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.GetWordState[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1214_  (.CLK(net1),
    .D(\INST_config_UART._0024_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.GetWordState[3] ));
 sky130_fd_sc_hd__dfrtp_4 \INST_config_UART._1215_  (.CLK(net1),
    .D(\INST_config_UART._0080_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceivedWord[5] ));
 sky130_fd_sc_hd__dfstp_2 \INST_config_UART._1216_  (.CLK(net1),
    .D(\INST_config_UART._0019_ ),
    .SET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1217_  (.CLK(net1),
    .D(\INST_config_UART._0020_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1218_  (.CLK(net1),
    .D(\INST_config_UART._0081_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceivedWord[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1219_  (.CLK(net1),
    .D(\INST_config_UART._0082_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1220_  (.CLK(net1),
    .D(\INST_config_UART._0083_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1221_  (.CLK(net1),
    .D(\INST_config_UART._0084_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1222_  (.CLK(net1),
    .D(\INST_config_UART._0085_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1223_  (.CLK(net1),
    .D(\INST_config_UART._0086_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1224_  (.CLK(net1),
    .D(\INST_config_UART._0087_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1225_  (.CLK(net1),
    .D(\INST_config_UART._0088_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1226_  (.CLK(net1),
    .D(\INST_config_UART._0089_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[23] ));
 sky130_fd_sc_hd__dfrtp_2 \INST_config_UART._1227_  (.CLK(net1),
    .D(\INST_config_UART._0090_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceivedWord[3] ));
 sky130_fd_sc_hd__dfrtp_4 \INST_config_UART._1228_  (.CLK(net1),
    .D(\INST_config_UART._0091_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceivedWord[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1229_  (.CLK(net1),
    .D(\INST_config_UART._0092_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceivedWord[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1230_  (.CLK(net1),
    .D(\INST_config_UART._0093_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1231_  (.CLK(net1),
    .D(\INST_config_UART._0094_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1232_  (.CLK(net1),
    .D(\INST_config_UART._0095_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1233_  (.CLK(net1),
    .D(\INST_config_UART._0096_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1234_  (.CLK(net1),
    .D(\INST_config_UART._0097_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1235_  (.CLK(net1),
    .D(\INST_config_UART._0098_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1236_  (.CLK(net1),
    .D(\INST_config_UART._0099_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1237_  (.CLK(net1),
    .D(\INST_config_UART._0100_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[15] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1238_  (.CLK(net1),
    .D(\INST_config_UART._0016_ ),
    .SET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceiveState ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1239_  (.CLK(net1),
    .D(\INST_config_UART._0101_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HighReg[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1240_  (.CLK(net1),
    .D(\INST_config_UART._0102_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HighReg[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1241_  (.CLK(net1),
    .D(\INST_config_UART._0103_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HighReg[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1242_  (.CLK(net1),
    .D(\INST_config_UART._0104_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HighReg[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1243_  (.CLK(net1),
    .D(\INST_config_UART._0014_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HexWriteStrobe ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1244_  (.CLK(net1),
    .D(\INST_config_UART._0105_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSend ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1245_  (.CLK(net1),
    .D(\INST_config_UART._0106_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HexData[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1246_  (.CLK(net1),
    .D(\INST_config_UART._0107_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HexData[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1247_  (.CLK(net1),
    .D(\INST_config_UART._0108_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HexData[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1248_  (.CLK(net1),
    .D(\INST_config_UART._0109_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HexData[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1249_  (.CLK(net1),
    .D(\INST_config_UART._0110_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HexData[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1250_  (.CLK(net1),
    .D(\INST_config_UART._0111_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HexData[5] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1251_  (.CLK(net1),
    .D(\INST_config_UART._0112_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HexData[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1252_  (.CLK(net1),
    .D(\INST_config_UART._0113_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.HexData[7] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1253_  (.CLK(net1),
    .D(\INST_config_UART._0114_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1254_  (.CLK(net1),
    .D(\INST_config_UART._0115_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1255_  (.CLK(net1),
    .D(\INST_config_UART._0116_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1256_  (.CLK(net1),
    .D(\INST_config_UART._0117_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1257_  (.CLK(net1),
    .D(\INST_config_UART._0118_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1258_  (.CLK(net1),
    .D(\INST_config_UART._0119_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[5] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1259_  (.CLK(net1),
    .D(\INST_config_UART._0120_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1260_  (.CLK(net1),
    .D(\INST_config_UART._0121_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[7] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1261_  (.CLK(net1),
    .D(\INST_config_UART._0122_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[8] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1262_  (.CLK(net1),
    .D(\INST_config_UART._0123_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[9] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1263_  (.CLK(net1),
    .D(\INST_config_UART._0124_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[10] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1264_  (.CLK(net1),
    .D(\INST_config_UART._0125_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[11] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1265_  (.CLK(net1),
    .D(\INST_config_UART._0126_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[12] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1266_  (.CLK(net1),
    .D(\INST_config_UART._0127_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[13] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1267_  (.CLK(net1),
    .D(\INST_config_UART._0128_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.TimeToSendCounter[14] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1268_  (.CLK(net1),
    .D(\INST_config_UART._0017_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteStrobe ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1269_  (.CLK(net1),
    .D(\INST_config_UART._0015_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.LocalWriteStrobe ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1270_  (.CLK(net1),
    .D(\INST_config_UART._0000_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ByteWriteStrobe ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1271_  (.CLK(net1),
    .D(\INST_config_UART._0129_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceiveLED ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1272_  (.CLK(net1),
    .D(\INST_config_UART._0130_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[24] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1273_  (.CLK(net1),
    .D(\INST_config_UART._0131_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[25] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1274_  (.CLK(net1),
    .D(\INST_config_UART._0132_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[26] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1275_  (.CLK(net1),
    .D(\INST_config_UART._0133_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[27] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1276_  (.CLK(net1),
    .D(\INST_config_UART._0134_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[28] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1277_  (.CLK(net1),
    .D(\INST_config_UART._0135_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[29] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1278_  (.CLK(net1),
    .D(\INST_config_UART._0136_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[30] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1279_  (.CLK(net1),
    .D(\INST_config_UART._0137_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.WriteData[31] ));
 sky130_fd_sc_hd__dfrtp_2 \INST_config_UART._1280_  (.CLK(net1),
    .D(\INST_config_UART._0031_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1281_  (.CLK(net1),
    .D(\INST_config_UART._0042_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1282_  (.CLK(net1),
    .D(\INST_config_UART._0046_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1283_  (.CLK(net1),
    .D(\INST_config_UART._0047_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1284_  (.CLK(net1),
    .D(\INST_config_UART._0048_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1285_  (.CLK(net1),
    .D(\INST_config_UART._0049_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[5] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1286_  (.CLK(net1),
    .D(\INST_config_UART._0050_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1287_  (.CLK(net1),
    .D(\INST_config_UART._0051_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[7] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1288_  (.CLK(net1),
    .D(\INST_config_UART._0052_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[8] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1289_  (.CLK(net1),
    .D(\INST_config_UART._0053_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[9] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1290_  (.CLK(net1),
    .D(\INST_config_UART._0032_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[10] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1291_  (.CLK(net1),
    .D(\INST_config_UART._0033_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[11] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1292_  (.CLK(net1),
    .D(\INST_config_UART._0034_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[12] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1293_  (.CLK(net1),
    .D(\INST_config_UART._0035_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[13] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1294_  (.CLK(net1),
    .D(\INST_config_UART._0036_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[14] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1295_  (.CLK(net1),
    .D(\INST_config_UART._0037_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[15] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1296_  (.CLK(net1),
    .D(\INST_config_UART._0038_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[16] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1297_  (.CLK(net1),
    .D(\INST_config_UART._0039_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[17] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1298_  (.CLK(net1),
    .D(\INST_config_UART._0040_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[18] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1299_  (.CLK(net1),
    .D(\INST_config_UART._0041_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[19] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1300_  (.CLK(net1),
    .D(\INST_config_UART._0043_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[20] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1301_  (.CLK(net1),
    .D(\INST_config_UART._0044_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[21] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1302_  (.CLK(net1),
    .D(\INST_config_UART._0045_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.blink[22] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1303_  (.CLK(net1),
    .D(\INST_config_UART._0138_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1304_  (.CLK(net1),
    .D(\INST_config_UART._0139_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1305_  (.CLK(net1),
    .D(\INST_config_UART._0140_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1306_  (.CLK(net1),
    .D(\INST_config_UART._0141_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1307_  (.CLK(net1),
    .D(\INST_config_UART._0142_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1308_  (.CLK(net1),
    .D(\INST_config_UART._0143_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[5] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1309_  (.CLK(net1),
    .D(\INST_config_UART._0144_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1310_  (.CLK(net1),
    .D(\INST_config_UART._0145_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[7] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1311_  (.CLK(net1),
    .D(\INST_config_UART._0146_ ),
    .SET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[8] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1312_  (.CLK(net1),
    .D(\INST_config_UART._0147_ ),
    .SET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[9] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1313_  (.CLK(net1),
    .D(\INST_config_UART._0148_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[10] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1314_  (.CLK(net1),
    .D(\INST_config_UART._0149_ ),
    .SET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[11] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1315_  (.CLK(net1),
    .D(\INST_config_UART._0150_ ),
    .SET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[12] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1316_  (.CLK(net1),
    .D(\INST_config_UART._0151_ ),
    .SET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[13] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1317_  (.CLK(net1),
    .D(\INST_config_UART._0152_ ),
    .SET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[14] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1318_  (.CLK(net1),
    .D(\INST_config_UART._0153_ ),
    .SET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[15] ));
 sky130_fd_sc_hd__dfrtp_2 \INST_config_UART._1319_  (.CLK(net1),
    .D(\INST_config_UART._0154_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[16] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1320_  (.CLK(net1),
    .D(\INST_config_UART._0155_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[17] ));
 sky130_fd_sc_hd__dfstp_1 \INST_config_UART._1321_  (.CLK(net1),
    .D(\INST_config_UART._0156_ ),
    .SET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[18] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1322_  (.CLK(net1),
    .D(\INST_config_UART._0157_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.CRCReg[19] ));
 sky130_fd_sc_hd__dfrtp_4 \INST_config_UART._1323_  (.CLK(net1),
    .D(\INST_config_UART._0158_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ReceivedWord[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1324_  (.CLK(net1),
    .D(\INST_config_UART._0159_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1325_  (.CLK(net1),
    .D(\INST_config_UART._0160_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1326_  (.CLK(net1),
    .D(\INST_config_UART._0161_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1327_  (.CLK(net1),
    .D(\INST_config_UART._0162_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1328_  (.CLK(net1),
    .D(\INST_config_UART._0163_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1329_  (.CLK(net1),
    .D(\INST_config_UART._0164_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1330_  (.CLK(net1),
    .D(\INST_config_UART._0165_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1331_  (.CLK(net1),
    .D(\INST_config_UART._0166_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ID_Reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1332_  (.CLK(net1),
    .D(\INST_config_UART._0167_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Command[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1333_  (.CLK(net1),
    .D(\INST_config_UART._0168_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Command[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1334_  (.CLK(net1),
    .D(\INST_config_UART._0169_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Command[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1335_  (.CLK(net1),
    .D(\INST_config_UART._0170_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Command[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1336_  (.CLK(net1),
    .D(\INST_config_UART._0171_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Command[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1337_  (.CLK(net1),
    .D(\INST_config_UART._0172_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Command[5] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1338_  (.CLK(net1),
    .D(\INST_config_UART._0173_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Command[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1339_  (.CLK(net1),
    .D(\INST_config_UART._0174_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Command[7] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1340_  (.CLK(net1),
    .D(\INST_config_UART._0001_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[0] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1341_  (.CLK(net1),
    .D(\INST_config_UART._0004_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[1] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1342_  (.CLK(net1),
    .D(\INST_config_UART._0005_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1343_  (.CLK(net1),
    .D(\INST_config_UART._0006_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1344_  (.CLK(net1),
    .D(\INST_config_UART._0007_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1345_  (.CLK(net1),
    .D(\INST_config_UART._0008_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[5] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1346_  (.CLK(net1),
    .D(\INST_config_UART._0009_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[6] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1347_  (.CLK(net1),
    .D(\INST_config_UART._0010_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[7] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1348_  (.CLK(net1),
    .D(\INST_config_UART._0011_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[8] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1349_  (.CLK(net1),
    .D(\INST_config_UART._0012_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[9] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1350_  (.CLK(net1),
    .D(\INST_config_UART._0002_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[10] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1351_  (.CLK(net1),
    .D(\INST_config_UART._0003_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComCount[11] ));
 sky130_fd_sc_hd__dfrtp_4 \INST_config_UART._1352_  (.CLK(net1),
    .D(\INST_config_UART._0013_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComTick ));
 sky130_fd_sc_hd__dfstp_4 \INST_config_UART._1353_  (.CLK(net1),
    .D(net2),
    .SET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.RxLocal ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1354_  (.CLK(net1),
    .D(\INST_config_UART._0175_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Data_Reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1355_  (.CLK(net1),
    .D(\INST_config_UART._0176_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Data_Reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1356_  (.CLK(net1),
    .D(\INST_config_UART._0177_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Data_Reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1357_  (.CLK(net1),
    .D(\INST_config_UART._0178_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Data_Reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1358_  (.CLK(net1),
    .D(\INST_config_UART._0179_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Data_Reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1359_  (.CLK(net1),
    .D(\INST_config_UART._0180_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Data_Reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1360_  (.CLK(net1),
    .D(\INST_config_UART._0181_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Data_Reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 \INST_config_UART._1361_  (.CLK(net1),
    .D(\INST_config_UART._0182_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.Data_Reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1362_  (.CLK(net1),
    .D(\INST_config_UART._0183_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[10] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1363_  (.CLK(net1),
    .D(\INST_config_UART._0184_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[9] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1364_  (.CLK(net1),
    .D(\INST_config_UART._0185_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[8] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1365_  (.CLK(net1),
    .D(\INST_config_UART._0186_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[7] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1366_  (.CLK(net1),
    .D(\INST_config_UART._0187_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[5] ));
 sky130_fd_sc_hd__dfrtp_2 \INST_config_UART._1367_  (.CLK(net1),
    .D(\INST_config_UART._0188_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[4] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1368_  (.CLK(net1),
    .D(\INST_config_UART._0189_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[3] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1369_  (.CLK(net1),
    .D(\INST_config_UART._0190_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[2] ));
 sky130_fd_sc_hd__dfrtp_1 \INST_config_UART._1370_  (.CLK(net1),
    .D(\INST_config_UART._0191_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\INST_config_UART.ComState[1] ));
 sky130_fd_sc_hd__and4_1 \Inst_bitbang._181_  (.A(\Inst_bitbang.serial_control[13] ),
    .B(\Inst_bitbang.serial_control[12] ),
    .C(\Inst_bitbang.serial_control[15] ),
    .D(\Inst_bitbang.serial_control[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._083_ ));
 sky130_fd_sc_hd__and4bb_1 \Inst_bitbang._182_  (.A_N(\Inst_bitbang.serial_control[8] ),
    .B_N(\Inst_bitbang.serial_control[10] ),
    .C(\Inst_bitbang.serial_control[11] ),
    .D(\Inst_bitbang.serial_control[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._084_ ));
 sky130_fd_sc_hd__and4b_1 \Inst_bitbang._183_  (.A_N(\Inst_bitbang.serial_control[6] ),
    .B(\Inst_bitbang.serial_control[7] ),
    .C(\Inst_bitbang.serial_control[5] ),
    .D(\Inst_bitbang.serial_control[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._085_ ));
 sky130_fd_sc_hd__nor4b_2 \Inst_bitbang._184_  (.A(\Inst_bitbang.serial_control[3] ),
    .B(\Inst_bitbang.serial_control[2] ),
    .C(\Inst_bitbang.serial_control[1] ),
    .D_N(\Inst_bitbang.serial_control[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_bitbang._086_ ));
 sky130_fd_sc_hd__nand4_4 \Inst_bitbang._185_  (.A(\Inst_bitbang._083_ ),
    .B(\Inst_bitbang._084_ ),
    .C(\Inst_bitbang._085_ ),
    .D(\Inst_bitbang._086_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_bitbang._087_ ));
 sky130_fd_sc_hd__buf_4 \Inst_bitbang._186_  (.A(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._088_ ));
 sky130_fd_sc_hd__inv_2 \Inst_bitbang._187_  (.A(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_bitbang._000_ ));
 sky130_fd_sc_hd__and2b_1 \Inst_bitbang._188_  (.A_N(\Inst_bitbang.old_local_strobe ),
    .B(\Inst_bitbang.local_strobe ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._089_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._189_  (.A(\Inst_bitbang._089_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._001_ ));
 sky130_fd_sc_hd__nor3_1 \Inst_bitbang._190_  (.A(\Inst_bitbang.serial_control[3] ),
    .B(\Inst_bitbang.serial_control[2] ),
    .C(\Inst_bitbang.serial_control[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_bitbang._090_ ));
 sky130_fd_sc_hd__inv_2 \Inst_bitbang._191_  (.A(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_bitbang._091_ ));
 sky130_fd_sc_hd__a41o_1 \Inst_bitbang._192_  (.A1(\Inst_bitbang._083_ ),
    .A2(\Inst_bitbang._084_ ),
    .A3(\Inst_bitbang._085_ ),
    .A4(\Inst_bitbang._090_ ),
    .B1(\Inst_bitbang._091_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._092_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_bitbang._193_  (.A(\Inst_bitbang._088_ ),
    .B(\Inst_bitbang._092_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_bitbang._002_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._194_  (.A0(\Inst_bitbang.serial_data[0] ),
    .A1(\Inst_bitbang.data[0] ),
    .S(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._093_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._195_  (.A(\Inst_bitbang._093_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._003_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._196_  (.A0(\Inst_bitbang.serial_data[1] ),
    .A1(\Inst_bitbang.data[1] ),
    .S(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._094_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._197_  (.A(\Inst_bitbang._094_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._004_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._198_  (.A0(\Inst_bitbang.serial_data[2] ),
    .A1(\Inst_bitbang.data[2] ),
    .S(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._095_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._199_  (.A(\Inst_bitbang._095_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._005_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._200_  (.A0(\Inst_bitbang.serial_data[3] ),
    .A1(\Inst_bitbang.data[3] ),
    .S(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._096_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._201_  (.A(\Inst_bitbang._096_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._006_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._202_  (.A0(\Inst_bitbang.serial_data[4] ),
    .A1(\Inst_bitbang.data[4] ),
    .S(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._097_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._203_  (.A(\Inst_bitbang._097_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._007_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._204_  (.A0(\Inst_bitbang.serial_data[5] ),
    .A1(\Inst_bitbang.data[5] ),
    .S(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._098_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._205_  (.A(\Inst_bitbang._098_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._008_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._206_  (.A0(\Inst_bitbang.serial_data[6] ),
    .A1(\Inst_bitbang.data[6] ),
    .S(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._099_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._207_  (.A(\Inst_bitbang._099_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._009_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._208_  (.A0(\Inst_bitbang.serial_data[7] ),
    .A1(\Inst_bitbang.data[7] ),
    .S(\Inst_bitbang._088_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._100_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._209_  (.A(\Inst_bitbang._100_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._010_ ));
 sky130_fd_sc_hd__buf_4 \Inst_bitbang._210_  (.A(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._101_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._211_  (.A0(\Inst_bitbang.serial_data[8] ),
    .A1(\Inst_bitbang.data[8] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._102_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._212_  (.A(\Inst_bitbang._102_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._011_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._213_  (.A0(\Inst_bitbang.serial_data[9] ),
    .A1(\Inst_bitbang.data[9] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._103_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._214_  (.A(\Inst_bitbang._103_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._012_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._215_  (.A0(\Inst_bitbang.serial_data[10] ),
    .A1(\Inst_bitbang.data[10] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._104_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._216_  (.A(\Inst_bitbang._104_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._013_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._217_  (.A0(\Inst_bitbang.serial_data[11] ),
    .A1(\Inst_bitbang.data[11] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._105_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._218_  (.A(\Inst_bitbang._105_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._014_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._219_  (.A0(\Inst_bitbang.serial_data[12] ),
    .A1(\Inst_bitbang.data[12] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._106_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._220_  (.A(\Inst_bitbang._106_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._015_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._221_  (.A0(\Inst_bitbang.serial_data[13] ),
    .A1(\Inst_bitbang.data[13] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._107_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._222_  (.A(\Inst_bitbang._107_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._016_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._223_  (.A0(\Inst_bitbang.serial_data[14] ),
    .A1(\Inst_bitbang.data[14] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._108_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._224_  (.A(\Inst_bitbang._108_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._017_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._225_  (.A0(\Inst_bitbang.serial_data[15] ),
    .A1(\Inst_bitbang.data[15] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._109_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._226_  (.A(\Inst_bitbang._109_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._018_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._227_  (.A0(\Inst_bitbang.serial_data[16] ),
    .A1(\Inst_bitbang.data[16] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._110_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._228_  (.A(\Inst_bitbang._110_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._019_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._229_  (.A0(\Inst_bitbang.serial_data[17] ),
    .A1(\Inst_bitbang.data[17] ),
    .S(\Inst_bitbang._101_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._111_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._230_  (.A(\Inst_bitbang._111_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._020_ ));
 sky130_fd_sc_hd__clkbuf_4 \Inst_bitbang._231_  (.A(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._112_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._232_  (.A0(\Inst_bitbang.serial_data[18] ),
    .A1(\Inst_bitbang.data[18] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._113_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._233_  (.A(\Inst_bitbang._113_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._021_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._234_  (.A0(\Inst_bitbang.serial_data[19] ),
    .A1(\Inst_bitbang.data[19] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._114_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._235_  (.A(\Inst_bitbang._114_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._022_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._236_  (.A0(\Inst_bitbang.serial_data[20] ),
    .A1(\Inst_bitbang.data[20] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._115_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._237_  (.A(\Inst_bitbang._115_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._023_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._238_  (.A0(\Inst_bitbang.serial_data[21] ),
    .A1(\Inst_bitbang.data[21] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._116_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._239_  (.A(\Inst_bitbang._116_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._024_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._240_  (.A0(\Inst_bitbang.serial_data[22] ),
    .A1(\Inst_bitbang.data[22] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._117_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._241_  (.A(\Inst_bitbang._117_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._025_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._242_  (.A0(\Inst_bitbang.serial_data[23] ),
    .A1(\Inst_bitbang.data[23] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._118_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._243_  (.A(\Inst_bitbang._118_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._026_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._244_  (.A0(\Inst_bitbang.serial_data[24] ),
    .A1(\Inst_bitbang.data[24] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._119_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._245_  (.A(\Inst_bitbang._119_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._027_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._246_  (.A0(\Inst_bitbang.serial_data[25] ),
    .A1(\Inst_bitbang.data[25] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._120_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._247_  (.A(\Inst_bitbang._120_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._028_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._248_  (.A0(\Inst_bitbang.serial_data[26] ),
    .A1(\Inst_bitbang.data[26] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._121_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._249_  (.A(\Inst_bitbang._121_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._029_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._250_  (.A0(\Inst_bitbang.serial_data[27] ),
    .A1(\Inst_bitbang.data[27] ),
    .S(\Inst_bitbang._112_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._122_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._251_  (.A(\Inst_bitbang._122_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._030_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._252_  (.A0(\Inst_bitbang.serial_data[28] ),
    .A1(\Inst_bitbang.data[28] ),
    .S(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._123_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._253_  (.A(\Inst_bitbang._123_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._031_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._254_  (.A0(\Inst_bitbang.serial_data[29] ),
    .A1(\Inst_bitbang.data[29] ),
    .S(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._124_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._255_  (.A(\Inst_bitbang._124_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._032_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._256_  (.A0(\Inst_bitbang.serial_data[30] ),
    .A1(\Inst_bitbang.data[30] ),
    .S(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._125_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._257_  (.A(\Inst_bitbang._125_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._033_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._258_  (.A0(\Inst_bitbang.serial_data[31] ),
    .A1(\Inst_bitbang.data[31] ),
    .S(\Inst_bitbang._087_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._126_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._259_  (.A(\Inst_bitbang._126_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._034_ ));
 sky130_fd_sc_hd__nand2b_4 \Inst_bitbang._260_  (.A_N(\Inst_bitbang.s_clk_sample[3] ),
    .B(\Inst_bitbang.s_clk_sample[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_bitbang._127_ ));
 sky130_fd_sc_hd__buf_4 \Inst_bitbang._261_  (.A(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._128_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._262_  (.A0(\Inst_bitbang.s_data_sample[3] ),
    .A1(\Inst_bitbang.serial_data[0] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._129_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._263_  (.A(\Inst_bitbang._129_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._035_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._264_  (.A0(\Inst_bitbang.serial_data[0] ),
    .A1(\Inst_bitbang.serial_data[1] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._130_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._265_  (.A(\Inst_bitbang._130_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._036_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._266_  (.A0(\Inst_bitbang.serial_data[1] ),
    .A1(\Inst_bitbang.serial_data[2] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._131_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._267_  (.A(\Inst_bitbang._131_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._037_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._268_  (.A0(\Inst_bitbang.serial_data[2] ),
    .A1(\Inst_bitbang.serial_data[3] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._132_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._269_  (.A(\Inst_bitbang._132_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._038_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._270_  (.A0(\Inst_bitbang.serial_data[3] ),
    .A1(\Inst_bitbang.serial_data[4] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._133_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._271_  (.A(\Inst_bitbang._133_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._039_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._272_  (.A0(\Inst_bitbang.serial_data[4] ),
    .A1(\Inst_bitbang.serial_data[5] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._134_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._273_  (.A(\Inst_bitbang._134_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._040_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._274_  (.A0(\Inst_bitbang.serial_data[5] ),
    .A1(\Inst_bitbang.serial_data[6] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._135_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._275_  (.A(\Inst_bitbang._135_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._041_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._276_  (.A0(\Inst_bitbang.serial_data[6] ),
    .A1(\Inst_bitbang.serial_data[7] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._136_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._277_  (.A(\Inst_bitbang._136_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._042_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._278_  (.A0(\Inst_bitbang.serial_data[7] ),
    .A1(\Inst_bitbang.serial_data[8] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._137_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._279_  (.A(\Inst_bitbang._137_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._043_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._280_  (.A0(\Inst_bitbang.serial_data[8] ),
    .A1(\Inst_bitbang.serial_data[9] ),
    .S(\Inst_bitbang._128_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._138_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._281_  (.A(\Inst_bitbang._138_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._044_ ));
 sky130_fd_sc_hd__clkbuf_4 \Inst_bitbang._282_  (.A(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._139_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._283_  (.A0(\Inst_bitbang.serial_data[9] ),
    .A1(\Inst_bitbang.serial_data[10] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._140_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._284_  (.A(\Inst_bitbang._140_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._045_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._285_  (.A0(\Inst_bitbang.serial_data[10] ),
    .A1(\Inst_bitbang.serial_data[11] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._141_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._286_  (.A(\Inst_bitbang._141_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._046_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._287_  (.A0(\Inst_bitbang.serial_data[11] ),
    .A1(\Inst_bitbang.serial_data[12] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._142_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._288_  (.A(\Inst_bitbang._142_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._047_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._289_  (.A0(\Inst_bitbang.serial_data[12] ),
    .A1(\Inst_bitbang.serial_data[13] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._143_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._290_  (.A(\Inst_bitbang._143_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._048_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._291_  (.A0(\Inst_bitbang.serial_data[13] ),
    .A1(\Inst_bitbang.serial_data[14] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._144_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._292_  (.A(\Inst_bitbang._144_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._049_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._293_  (.A0(\Inst_bitbang.serial_data[14] ),
    .A1(\Inst_bitbang.serial_data[15] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._145_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._294_  (.A(\Inst_bitbang._145_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._050_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._295_  (.A0(\Inst_bitbang.serial_data[15] ),
    .A1(\Inst_bitbang.serial_data[16] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._146_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._296_  (.A(\Inst_bitbang._146_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._051_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._297_  (.A0(\Inst_bitbang.serial_data[16] ),
    .A1(\Inst_bitbang.serial_data[17] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._147_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._298_  (.A(\Inst_bitbang._147_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._052_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._299_  (.A0(\Inst_bitbang.serial_data[17] ),
    .A1(\Inst_bitbang.serial_data[18] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._148_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._300_  (.A(\Inst_bitbang._148_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._053_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._301_  (.A0(\Inst_bitbang.serial_data[18] ),
    .A1(\Inst_bitbang.serial_data[19] ),
    .S(\Inst_bitbang._139_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._149_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._302_  (.A(\Inst_bitbang._149_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._054_ ));
 sky130_fd_sc_hd__clkbuf_4 \Inst_bitbang._303_  (.A(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._150_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._304_  (.A0(\Inst_bitbang.serial_data[19] ),
    .A1(\Inst_bitbang.serial_data[20] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._151_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._305_  (.A(\Inst_bitbang._151_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._055_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._306_  (.A0(\Inst_bitbang.serial_data[20] ),
    .A1(\Inst_bitbang.serial_data[21] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._152_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._307_  (.A(\Inst_bitbang._152_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._056_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._308_  (.A0(\Inst_bitbang.serial_data[21] ),
    .A1(\Inst_bitbang.serial_data[22] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._153_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._309_  (.A(\Inst_bitbang._153_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._057_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._310_  (.A0(\Inst_bitbang.serial_data[22] ),
    .A1(\Inst_bitbang.serial_data[23] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._154_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._311_  (.A(\Inst_bitbang._154_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._058_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._312_  (.A0(\Inst_bitbang.serial_data[23] ),
    .A1(\Inst_bitbang.serial_data[24] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._155_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._313_  (.A(\Inst_bitbang._155_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._059_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._314_  (.A0(\Inst_bitbang.serial_data[24] ),
    .A1(\Inst_bitbang.serial_data[25] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._156_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._315_  (.A(\Inst_bitbang._156_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._060_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._316_  (.A0(\Inst_bitbang.serial_data[25] ),
    .A1(\Inst_bitbang.serial_data[26] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._157_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._317_  (.A(\Inst_bitbang._157_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._061_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._318_  (.A0(\Inst_bitbang.serial_data[26] ),
    .A1(\Inst_bitbang.serial_data[27] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._158_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._319_  (.A(\Inst_bitbang._158_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._062_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._320_  (.A0(\Inst_bitbang.serial_data[27] ),
    .A1(\Inst_bitbang.serial_data[28] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._159_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._321_  (.A(\Inst_bitbang._159_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._063_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._322_  (.A0(\Inst_bitbang.serial_data[28] ),
    .A1(\Inst_bitbang.serial_data[29] ),
    .S(\Inst_bitbang._150_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._160_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._323_  (.A(\Inst_bitbang._160_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._064_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._324_  (.A0(\Inst_bitbang.serial_data[29] ),
    .A1(\Inst_bitbang.serial_data[30] ),
    .S(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._161_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._325_  (.A(\Inst_bitbang._161_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._065_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._326_  (.A0(\Inst_bitbang.serial_data[30] ),
    .A1(\Inst_bitbang.serial_data[31] ),
    .S(\Inst_bitbang._127_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._162_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._327_  (.A(\Inst_bitbang._162_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._066_ ));
 sky130_fd_sc_hd__nand2b_4 \Inst_bitbang._328_  (.A_N(\Inst_bitbang.s_clk_sample[2] ),
    .B(\Inst_bitbang.s_clk_sample[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_bitbang._163_ ));
 sky130_fd_sc_hd__clkbuf_4 \Inst_bitbang._329_  (.A(\Inst_bitbang._163_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._164_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._330_  (.A0(\Inst_bitbang.s_data_sample[3] ),
    .A1(\Inst_bitbang.serial_control[0] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._165_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._331_  (.A(\Inst_bitbang._165_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._067_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._332_  (.A0(\Inst_bitbang.serial_control[0] ),
    .A1(\Inst_bitbang.serial_control[1] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._166_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._333_  (.A(\Inst_bitbang._166_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._068_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._334_  (.A0(\Inst_bitbang.serial_control[1] ),
    .A1(\Inst_bitbang.serial_control[2] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._167_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._335_  (.A(\Inst_bitbang._167_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._069_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._336_  (.A0(\Inst_bitbang.serial_control[2] ),
    .A1(\Inst_bitbang.serial_control[3] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._168_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._337_  (.A(\Inst_bitbang._168_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._070_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._338_  (.A0(\Inst_bitbang.serial_control[3] ),
    .A1(\Inst_bitbang.serial_control[4] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._169_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._339_  (.A(\Inst_bitbang._169_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._071_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._340_  (.A0(\Inst_bitbang.serial_control[4] ),
    .A1(\Inst_bitbang.serial_control[5] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._170_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._341_  (.A(\Inst_bitbang._170_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._072_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._342_  (.A0(\Inst_bitbang.serial_control[5] ),
    .A1(\Inst_bitbang.serial_control[6] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._171_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._343_  (.A(\Inst_bitbang._171_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._073_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._344_  (.A0(\Inst_bitbang.serial_control[6] ),
    .A1(\Inst_bitbang.serial_control[7] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._172_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._345_  (.A(\Inst_bitbang._172_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._074_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._346_  (.A0(\Inst_bitbang.serial_control[7] ),
    .A1(\Inst_bitbang.serial_control[8] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._173_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._347_  (.A(\Inst_bitbang._173_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._075_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._348_  (.A0(\Inst_bitbang.serial_control[8] ),
    .A1(\Inst_bitbang.serial_control[9] ),
    .S(\Inst_bitbang._164_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._174_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._349_  (.A(\Inst_bitbang._174_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._076_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._350_  (.A0(\Inst_bitbang.serial_control[9] ),
    .A1(\Inst_bitbang.serial_control[10] ),
    .S(\Inst_bitbang._163_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._175_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._351_  (.A(\Inst_bitbang._175_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._077_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._352_  (.A0(\Inst_bitbang.serial_control[10] ),
    .A1(\Inst_bitbang.serial_control[11] ),
    .S(\Inst_bitbang._163_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._176_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._353_  (.A(\Inst_bitbang._176_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._078_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._354_  (.A0(\Inst_bitbang.serial_control[11] ),
    .A1(\Inst_bitbang.serial_control[12] ),
    .S(\Inst_bitbang._163_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._177_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._355_  (.A(\Inst_bitbang._177_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._079_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._356_  (.A0(\Inst_bitbang.serial_control[12] ),
    .A1(\Inst_bitbang.serial_control[13] ),
    .S(\Inst_bitbang._163_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._178_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._357_  (.A(\Inst_bitbang._178_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._080_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._358_  (.A0(\Inst_bitbang.serial_control[13] ),
    .A1(\Inst_bitbang.serial_control[14] ),
    .S(\Inst_bitbang._163_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._179_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._359_  (.A(\Inst_bitbang._179_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._081_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_bitbang._360_  (.A0(\Inst_bitbang.serial_control[14] ),
    .A1(\Inst_bitbang.serial_control[15] ),
    .S(\Inst_bitbang._163_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._180_ ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_bitbang._361_  (.A(\Inst_bitbang._180_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_bitbang._082_ ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._362_  (.CLK(net1),
    .D(\Inst_bitbang._001_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.strobe ));
 sky130_fd_sc_hd__dfrtp_4 \Inst_bitbang._363_  (.CLK(net1),
    .D(\Inst_bitbang._002_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.active ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._364_  (.CLK(net1),
    .D(\Inst_bitbang._000_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.local_strobe ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._365_  (.CLK(net1),
    .D(\Inst_bitbang.local_strobe ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.old_local_strobe ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._366_  (.CLK(net1),
    .D(\Inst_bitbang._003_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[0] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._367_  (.CLK(net1),
    .D(\Inst_bitbang._004_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[1] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._368_  (.CLK(net1),
    .D(\Inst_bitbang._005_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[2] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._369_  (.CLK(net1),
    .D(\Inst_bitbang._006_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[3] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._370_  (.CLK(net1),
    .D(\Inst_bitbang._007_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[4] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._371_  (.CLK(net1),
    .D(\Inst_bitbang._008_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[5] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._372_  (.CLK(net1),
    .D(\Inst_bitbang._009_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[6] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._373_  (.CLK(net1),
    .D(\Inst_bitbang._010_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[7] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._374_  (.CLK(net1),
    .D(\Inst_bitbang._011_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[8] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._375_  (.CLK(net1),
    .D(\Inst_bitbang._012_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[9] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._376_  (.CLK(net1),
    .D(\Inst_bitbang._013_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[10] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._377_  (.CLK(net1),
    .D(\Inst_bitbang._014_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[11] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._378_  (.CLK(net1),
    .D(\Inst_bitbang._015_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[12] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._379_  (.CLK(net1),
    .D(\Inst_bitbang._016_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[13] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._380_  (.CLK(net1),
    .D(\Inst_bitbang._017_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[14] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._381_  (.CLK(net1),
    .D(\Inst_bitbang._018_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[15] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._382_  (.CLK(net1),
    .D(\Inst_bitbang._019_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[16] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._383_  (.CLK(net1),
    .D(\Inst_bitbang._020_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[17] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._384_  (.CLK(net1),
    .D(\Inst_bitbang._021_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[18] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._385_  (.CLK(net1),
    .D(\Inst_bitbang._022_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[19] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._386_  (.CLK(net1),
    .D(\Inst_bitbang._023_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[20] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._387_  (.CLK(net1),
    .D(\Inst_bitbang._024_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[21] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._388_  (.CLK(net1),
    .D(\Inst_bitbang._025_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[22] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._389_  (.CLK(net1),
    .D(\Inst_bitbang._026_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[23] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._390_  (.CLK(net1),
    .D(\Inst_bitbang._027_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[24] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._391_  (.CLK(net1),
    .D(\Inst_bitbang._028_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[25] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._392_  (.CLK(net1),
    .D(\Inst_bitbang._029_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[26] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._393_  (.CLK(net1),
    .D(\Inst_bitbang._030_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[27] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._394_  (.CLK(net1),
    .D(\Inst_bitbang._031_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[28] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._395_  (.CLK(net1),
    .D(\Inst_bitbang._032_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[29] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._396_  (.CLK(net1),
    .D(\Inst_bitbang._033_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[30] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._397_  (.CLK(net1),
    .D(\Inst_bitbang._034_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.data[31] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._398_  (.CLK(net1),
    .D(\Inst_bitbang._035_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._399_  (.CLK(net1),
    .D(\Inst_bitbang._036_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._400_  (.CLK(net1),
    .D(\Inst_bitbang._037_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._401_  (.CLK(net1),
    .D(\Inst_bitbang._038_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._402_  (.CLK(net1),
    .D(\Inst_bitbang._039_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._403_  (.CLK(net1),
    .D(\Inst_bitbang._040_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._404_  (.CLK(net1),
    .D(\Inst_bitbang._041_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._405_  (.CLK(net1),
    .D(\Inst_bitbang._042_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._406_  (.CLK(net1),
    .D(\Inst_bitbang._043_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._407_  (.CLK(net1),
    .D(\Inst_bitbang._044_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._408_  (.CLK(net1),
    .D(\Inst_bitbang._045_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._409_  (.CLK(net1),
    .D(\Inst_bitbang._046_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._410_  (.CLK(net1),
    .D(\Inst_bitbang._047_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._411_  (.CLK(net1),
    .D(\Inst_bitbang._048_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._412_  (.CLK(net1),
    .D(\Inst_bitbang._049_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._413_  (.CLK(net1),
    .D(\Inst_bitbang._050_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._414_  (.CLK(net1),
    .D(\Inst_bitbang._051_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[16] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._415_  (.CLK(net1),
    .D(\Inst_bitbang._052_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[17] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._416_  (.CLK(net1),
    .D(\Inst_bitbang._053_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[18] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._417_  (.CLK(net1),
    .D(\Inst_bitbang._054_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[19] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._418_  (.CLK(net1),
    .D(\Inst_bitbang._055_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[20] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._419_  (.CLK(net1),
    .D(\Inst_bitbang._056_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[21] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._420_  (.CLK(net1),
    .D(\Inst_bitbang._057_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[22] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._421_  (.CLK(net1),
    .D(\Inst_bitbang._058_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[23] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._422_  (.CLK(net1),
    .D(\Inst_bitbang._059_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[24] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._423_  (.CLK(net1),
    .D(\Inst_bitbang._060_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[25] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._424_  (.CLK(net1),
    .D(\Inst_bitbang._061_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[26] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._425_  (.CLK(net1),
    .D(\Inst_bitbang._062_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[27] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._426_  (.CLK(net1),
    .D(\Inst_bitbang._063_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[28] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._427_  (.CLK(net1),
    .D(\Inst_bitbang._064_ ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[29] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._428_  (.CLK(net1),
    .D(\Inst_bitbang._065_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[30] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._429_  (.CLK(net1),
    .D(\Inst_bitbang._066_ ),
    .RESET_B(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_data[31] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._430_  (.CLK(net1),
    .D(net38),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.s_data_sample[0] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._431_  (.CLK(net1),
    .D(\Inst_bitbang.s_data_sample[0] ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.s_data_sample[1] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._432_  (.CLK(net1),
    .D(\Inst_bitbang.s_data_sample[1] ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.s_data_sample[2] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._433_  (.CLK(net1),
    .D(\Inst_bitbang.s_data_sample[2] ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.s_data_sample[3] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._434_  (.CLK(net1),
    .D(net37),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.s_clk_sample[0] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._435_  (.CLK(net1),
    .D(\Inst_bitbang.s_clk_sample[0] ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.s_clk_sample[1] ));
 sky130_fd_sc_hd__dfrtp_2 \Inst_bitbang._436_  (.CLK(net1),
    .D(\Inst_bitbang.s_clk_sample[1] ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.s_clk_sample[2] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._437_  (.CLK(net1),
    .D(\Inst_bitbang.s_clk_sample[2] ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.s_clk_sample[3] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._438_  (.CLK(net1),
    .D(\Inst_bitbang._067_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[0] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._439_  (.CLK(net1),
    .D(\Inst_bitbang._068_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[1] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._440_  (.CLK(net1),
    .D(\Inst_bitbang._069_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[2] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._441_  (.CLK(net1),
    .D(\Inst_bitbang._070_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[3] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._442_  (.CLK(net1),
    .D(\Inst_bitbang._071_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[4] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._443_  (.CLK(net1),
    .D(\Inst_bitbang._072_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[5] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._444_  (.CLK(net1),
    .D(\Inst_bitbang._073_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[6] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._445_  (.CLK(net1),
    .D(\Inst_bitbang._074_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[7] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._446_  (.CLK(net1),
    .D(\Inst_bitbang._075_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[8] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._447_  (.CLK(net1),
    .D(\Inst_bitbang._076_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[9] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._448_  (.CLK(net1),
    .D(\Inst_bitbang._077_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[10] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._449_  (.CLK(net1),
    .D(\Inst_bitbang._078_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[11] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._450_  (.CLK(net1),
    .D(\Inst_bitbang._079_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[12] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._451_  (.CLK(net1),
    .D(\Inst_bitbang._080_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[13] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._452_  (.CLK(net1),
    .D(\Inst_bitbang._081_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[14] ));
 sky130_fd_sc_hd__dfrtp_1 \Inst_bitbang._453_  (.CLK(net1),
    .D(\Inst_bitbang._082_ ),
    .RESET_B(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_bitbang.serial_control[15] ));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_4 _073_ (.A(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_000_));
 sky130_fd_sc_hd__clkbuf_4 _074_ (.A(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_001_));
 sky130_fd_sc_hd__or2_1 _075_ (.A(_000_),
    .B(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_002_));
 sky130_fd_sc_hd__buf_1 _076_ (.A(_002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.FSM_Reset ));
 sky130_fd_sc_hd__mux2_1 _077_ (.A0(net3),
    .A1(\Inst_bitbang.data[0] ),
    .S(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _078_ (.A0(_003_),
    .A1(\INST_config_UART.WriteData[0] ),
    .S(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_004_));
 sky130_fd_sc_hd__buf_2 _079_ (.A(_004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[0] ));
 sky130_fd_sc_hd__mux2_1 _080_ (.A0(net14),
    .A1(\Inst_bitbang.data[1] ),
    .S(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _081_ (.A0(_005_),
    .A1(\INST_config_UART.WriteData[1] ),
    .S(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_006_));
 sky130_fd_sc_hd__buf_2 _082_ (.A(_006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[1] ));
 sky130_fd_sc_hd__mux2_1 _083_ (.A0(net25),
    .A1(\Inst_bitbang.data[2] ),
    .S(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _084_ (.A0(_007_),
    .A1(\INST_config_UART.WriteData[2] ),
    .S(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_008_));
 sky130_fd_sc_hd__buf_2 _085_ (.A(_008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[2] ));
 sky130_fd_sc_hd__mux2_1 _086_ (.A0(net28),
    .A1(\Inst_bitbang.data[3] ),
    .S(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _087_ (.A0(_009_),
    .A1(\INST_config_UART.WriteData[3] ),
    .S(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_010_));
 sky130_fd_sc_hd__buf_2 _088_ (.A(_010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[3] ));
 sky130_fd_sc_hd__mux2_1 _089_ (.A0(net29),
    .A1(\Inst_bitbang.data[4] ),
    .S(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _090_ (.A0(_011_),
    .A1(\INST_config_UART.WriteData[4] ),
    .S(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_012_));
 sky130_fd_sc_hd__buf_2 _091_ (.A(_012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[4] ));
 sky130_fd_sc_hd__mux2_1 _092_ (.A0(net30),
    .A1(\Inst_bitbang.data[5] ),
    .S(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _093_ (.A0(_013_),
    .A1(\INST_config_UART.WriteData[5] ),
    .S(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_014_));
 sky130_fd_sc_hd__buf_2 _094_ (.A(_014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[5] ));
 sky130_fd_sc_hd__mux2_1 _095_ (.A0(net31),
    .A1(\Inst_bitbang.data[6] ),
    .S(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _096_ (.A0(_015_),
    .A1(\INST_config_UART.WriteData[6] ),
    .S(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_016_));
 sky130_fd_sc_hd__buf_2 _097_ (.A(_016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[6] ));
 sky130_fd_sc_hd__mux2_1 _098_ (.A0(net32),
    .A1(\Inst_bitbang.data[7] ),
    .S(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _099_ (.A0(_017_),
    .A1(\INST_config_UART.WriteData[7] ),
    .S(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_018_));
 sky130_fd_sc_hd__buf_2 _100_ (.A(_018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[7] ));
 sky130_fd_sc_hd__mux2_1 _101_ (.A0(net33),
    .A1(\Inst_bitbang.data[8] ),
    .S(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _102_ (.A0(_019_),
    .A1(\INST_config_UART.WriteData[8] ),
    .S(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_020_));
 sky130_fd_sc_hd__buf_2 _103_ (.A(_020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[8] ));
 sky130_fd_sc_hd__buf_4 _104_ (.A(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _105_ (.A0(net34),
    .A1(\Inst_bitbang.data[9] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_022_));
 sky130_fd_sc_hd__clkbuf_4 _106_ (.A(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _107_ (.A0(_022_),
    .A1(\INST_config_UART.WriteData[9] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_024_));
 sky130_fd_sc_hd__buf_2 _108_ (.A(_024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[9] ));
 sky130_fd_sc_hd__mux2_1 _109_ (.A0(net4),
    .A1(\Inst_bitbang.data[10] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _110_ (.A0(_025_),
    .A1(\INST_config_UART.WriteData[10] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_026_));
 sky130_fd_sc_hd__buf_2 _111_ (.A(_026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[10] ));
 sky130_fd_sc_hd__mux2_1 _112_ (.A0(net5),
    .A1(\Inst_bitbang.data[11] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _113_ (.A0(_027_),
    .A1(\INST_config_UART.WriteData[11] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_028_));
 sky130_fd_sc_hd__buf_2 _114_ (.A(_028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[11] ));
 sky130_fd_sc_hd__mux2_1 _115_ (.A0(net6),
    .A1(\Inst_bitbang.data[12] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _116_ (.A0(_029_),
    .A1(\INST_config_UART.WriteData[12] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_030_));
 sky130_fd_sc_hd__buf_2 _117_ (.A(_030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[12] ));
 sky130_fd_sc_hd__mux2_1 _118_ (.A0(net7),
    .A1(\Inst_bitbang.data[13] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _119_ (.A0(_031_),
    .A1(\INST_config_UART.WriteData[13] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_032_));
 sky130_fd_sc_hd__clkbuf_2 _120_ (.A(_032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[13] ));
 sky130_fd_sc_hd__mux2_1 _121_ (.A0(net8),
    .A1(\Inst_bitbang.data[14] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _122_ (.A0(_033_),
    .A1(\INST_config_UART.WriteData[14] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_034_));
 sky130_fd_sc_hd__buf_2 _123_ (.A(_034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[14] ));
 sky130_fd_sc_hd__mux2_1 _124_ (.A0(net9),
    .A1(\Inst_bitbang.data[15] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _125_ (.A0(_035_),
    .A1(\INST_config_UART.WriteData[15] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_036_));
 sky130_fd_sc_hd__clkbuf_2 _126_ (.A(_036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[15] ));
 sky130_fd_sc_hd__mux2_1 _127_ (.A0(net10),
    .A1(\Inst_bitbang.data[16] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _128_ (.A0(_037_),
    .A1(\INST_config_UART.WriteData[16] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_038_));
 sky130_fd_sc_hd__clkbuf_2 _129_ (.A(_038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[16] ));
 sky130_fd_sc_hd__mux2_1 _130_ (.A0(net11),
    .A1(\Inst_bitbang.data[17] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _131_ (.A0(_039_),
    .A1(\INST_config_UART.WriteData[17] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_040_));
 sky130_fd_sc_hd__clkbuf_2 _132_ (.A(_040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[17] ));
 sky130_fd_sc_hd__mux2_1 _133_ (.A0(net12),
    .A1(\Inst_bitbang.data[18] ),
    .S(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _134_ (.A0(_041_),
    .A1(\INST_config_UART.WriteData[18] ),
    .S(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_042_));
 sky130_fd_sc_hd__clkbuf_2 _135_ (.A(_042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[18] ));
 sky130_fd_sc_hd__clkbuf_4 _136_ (.A(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _137_ (.A0(net13),
    .A1(\Inst_bitbang.data[19] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_044_));
 sky130_fd_sc_hd__clkbuf_4 _138_ (.A(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _139_ (.A0(_044_),
    .A1(\INST_config_UART.WriteData[19] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_046_));
 sky130_fd_sc_hd__clkbuf_2 _140_ (.A(_046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[19] ));
 sky130_fd_sc_hd__mux2_1 _141_ (.A0(net15),
    .A1(\Inst_bitbang.data[20] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _142_ (.A0(_047_),
    .A1(\INST_config_UART.WriteData[20] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_2 _143_ (.A(_048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[20] ));
 sky130_fd_sc_hd__mux2_1 _144_ (.A0(net16),
    .A1(\Inst_bitbang.data[21] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _145_ (.A0(_049_),
    .A1(\INST_config_UART.WriteData[21] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_050_));
 sky130_fd_sc_hd__clkbuf_2 _146_ (.A(_050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[21] ));
 sky130_fd_sc_hd__mux2_1 _147_ (.A0(net17),
    .A1(\Inst_bitbang.data[22] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _148_ (.A0(_051_),
    .A1(\INST_config_UART.WriteData[22] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_052_));
 sky130_fd_sc_hd__clkbuf_2 _149_ (.A(_052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[22] ));
 sky130_fd_sc_hd__mux2_1 _150_ (.A0(net18),
    .A1(\Inst_bitbang.data[23] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _151_ (.A0(_053_),
    .A1(\INST_config_UART.WriteData[23] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_054_));
 sky130_fd_sc_hd__clkbuf_2 _152_ (.A(_054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[23] ));
 sky130_fd_sc_hd__mux2_1 _153_ (.A0(net19),
    .A1(\Inst_bitbang.data[24] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _154_ (.A0(_055_),
    .A1(\INST_config_UART.WriteData[24] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_056_));
 sky130_fd_sc_hd__clkbuf_2 _155_ (.A(_056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[24] ));
 sky130_fd_sc_hd__mux2_1 _156_ (.A0(net20),
    .A1(\Inst_bitbang.data[25] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _157_ (.A0(_057_),
    .A1(\INST_config_UART.WriteData[25] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_058_));
 sky130_fd_sc_hd__clkbuf_2 _158_ (.A(_058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[25] ));
 sky130_fd_sc_hd__mux2_1 _159_ (.A0(net21),
    .A1(\Inst_bitbang.data[26] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _160_ (.A0(_059_),
    .A1(\INST_config_UART.WriteData[26] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_060_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _161_ (.A(_060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[26] ));
 sky130_fd_sc_hd__mux2_1 _162_ (.A0(net22),
    .A1(\Inst_bitbang.data[27] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _163_ (.A0(_061_),
    .A1(\INST_config_UART.WriteData[27] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_062_));
 sky130_fd_sc_hd__buf_1 _164_ (.A(_062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[27] ));
 sky130_fd_sc_hd__mux2_1 _165_ (.A0(net23),
    .A1(\Inst_bitbang.data[28] ),
    .S(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _166_ (.A0(_063_),
    .A1(\INST_config_UART.WriteData[28] ),
    .S(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_064_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _167_ (.A(_064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[28] ));
 sky130_fd_sc_hd__mux2_1 _168_ (.A0(net24),
    .A1(\Inst_bitbang.data[29] ),
    .S(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _169_ (.A0(_065_),
    .A1(\INST_config_UART.WriteData[29] ),
    .S(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_066_));
 sky130_fd_sc_hd__buf_1 _170_ (.A(_066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[29] ));
 sky130_fd_sc_hd__mux2_1 _171_ (.A0(net26),
    .A1(\Inst_bitbang.data[30] ),
    .S(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _172_ (.A0(_067_),
    .A1(\INST_config_UART.WriteData[30] ),
    .S(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_068_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _173_ (.A(_068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[30] ));
 sky130_fd_sc_hd__mux2_1 _174_ (.A0(net27),
    .A1(\Inst_bitbang.data[31] ),
    .S(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _175_ (.A0(_069_),
    .A1(\INST_config_UART.WriteData[31] ),
    .S(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_070_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _176_ (.A(_070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\ConfigFSM_inst.WriteData[31] ));
 sky130_fd_sc_hd__mux2_1 _177_ (.A0(net35),
    .A1(\Inst_bitbang.strobe ),
    .S(\Inst_bitbang.active ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _178_ (.A0(_071_),
    .A1(\INST_config_UART.WriteStrobe ),
    .S(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_072_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _179_ (.A(_072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net72));
 sky130_fd_sc_hd__xor2_1 _180_ (.A(\Inst_bitbang.strobe ),
    .B(\INST_config_UART.ReceiveLED ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 _181_ (.A(\ConfigFSM_inst.WriteData[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 _182_ (.A(\ConfigFSM_inst.WriteData[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _183_ (.A(\ConfigFSM_inst.WriteData[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _184_ (.A(\ConfigFSM_inst.WriteData[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _185_ (.A(\ConfigFSM_inst.WriteData[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _186_ (.A(\ConfigFSM_inst.WriteData[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _187_ (.A(\ConfigFSM_inst.WriteData[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _188_ (.A(\ConfigFSM_inst.WriteData[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _189_ (.A(\ConfigFSM_inst.WriteData[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _190_ (.A(\ConfigFSM_inst.WriteData[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _191_ (.A(\ConfigFSM_inst.WriteData[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 _192_ (.A(\ConfigFSM_inst.WriteData[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _193_ (.A(\ConfigFSM_inst.WriteData[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 _194_ (.A(\ConfigFSM_inst.WriteData[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 _195_ (.A(\ConfigFSM_inst.WriteData[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 _196_ (.A(\ConfigFSM_inst.WriteData[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 _197_ (.A(\ConfigFSM_inst.WriteData[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 _198_ (.A(\ConfigFSM_inst.WriteData[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 _199_ (.A(\ConfigFSM_inst.WriteData[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _200_ (.A(\ConfigFSM_inst.WriteData[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _201_ (.A(\ConfigFSM_inst.WriteData[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _202_ (.A(\ConfigFSM_inst.WriteData[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _203_ (.A(\ConfigFSM_inst.WriteData[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _204_ (.A(\ConfigFSM_inst.WriteData[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _205_ (.A(\ConfigFSM_inst.WriteData[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _206_ (.A(\ConfigFSM_inst.WriteData[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 _207_ (.A(\ConfigFSM_inst.WriteData[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _208_ (.A(\ConfigFSM_inst.WriteData[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _209_ (.A(\ConfigFSM_inst.WriteData[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 _210_ (.A(\ConfigFSM_inst.WriteData[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _211_ (.A(\ConfigFSM_inst.WriteData[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _212_ (.A(\ConfigFSM_inst.WriteData[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _213_ (.A(\ConfigFSM_inst.FrameAddressRegister[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _214_ (.A(\ConfigFSM_inst.FrameAddressRegister[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _215_ (.A(\ConfigFSM_inst.FrameAddressRegister[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _216_ (.A(\ConfigFSM_inst.FrameAddressRegister[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _217_ (.A(\ConfigFSM_inst.FrameAddressRegister[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _218_ (.A(\ConfigFSM_inst.FrameAddressRegister[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _219_ (.A(\ConfigFSM_inst.FrameAddressRegister[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _220_ (.A(\ConfigFSM_inst.FrameAddressRegister[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _221_ (.A(\ConfigFSM_inst.FrameAddressRegister[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _222_ (.A(\ConfigFSM_inst.FrameAddressRegister[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _223_ (.A(\ConfigFSM_inst.FrameAddressRegister[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _224_ (.A(\ConfigFSM_inst.FrameAddressRegister[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _225_ (.A(\ConfigFSM_inst.FrameAddressRegister[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _226_ (.A(\ConfigFSM_inst.FrameAddressRegister[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _227_ (.A(\ConfigFSM_inst.FrameAddressRegister[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _228_ (.A(\ConfigFSM_inst.FrameAddressRegister[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _229_ (.A(\ConfigFSM_inst.FrameAddressRegister[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _230_ (.A(\ConfigFSM_inst.FrameAddressRegister[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _231_ (.A(\ConfigFSM_inst.FrameAddressRegister[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _232_ (.A(\ConfigFSM_inst.FrameAddressRegister[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net83));
 sky130_fd_sc_hd__buf_2 _233_ (.A(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[20]));
 sky130_fd_sc_hd__conb_1 _233__113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net113));
 sky130_fd_sc_hd__clkbuf_1 _234_ (.A(\ConfigFSM_inst.FrameAddressRegister[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _235_ (.A(\ConfigFSM_inst.FrameAddressRegister[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _236_ (.A(\ConfigFSM_inst.FrameAddressRegister[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _237_ (.A(\ConfigFSM_inst.FrameAddressRegister[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _238_ (.A(\ConfigFSM_inst.FrameAddressRegister[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _239_ (.A(\ConfigFSM_inst.FrameAddressRegister[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _240_ (.A(\ConfigFSM_inst.FrameAddressRegister[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _241_ (.A(\ConfigFSM_inst.FrameAddressRegister[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _242_ (.A(\ConfigFSM_inst.FrameAddressRegister[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _243_ (.A(\ConfigFSM_inst.FrameAddressRegister[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _244_ (.A(\ConfigFSM_inst.FrameAddressRegister[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(\ConfigFSM_inst.RowSelect[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 _246_ (.A(\ConfigFSM_inst.RowSelect[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 _247_ (.A(\ConfigFSM_inst.RowSelect[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 _248_ (.A(\ConfigFSM_inst.RowSelect[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 _249_ (.A(\ConfigFSM_inst.RowSelect[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_16 input1 (.A(CLK),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(SelfWriteData[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(SelfWriteData[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(SelfWriteData[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(SelfWriteData[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(SelfWriteData[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(SelfWriteData[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(SelfWriteData[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(SelfWriteData[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(SelfWriteData[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(SelfWriteData[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(Rx),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(SelfWriteData[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(SelfWriteData[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(SelfWriteData[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(SelfWriteData[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(SelfWriteData[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(SelfWriteData[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(SelfWriteData[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(SelfWriteData[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(SelfWriteData[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(SelfWriteData[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(SelfWriteData[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(SelfWriteData[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(SelfWriteData[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(SelfWriteData[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(SelfWriteData[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(SelfWriteData[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(SelfWriteStrobe),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_16 input36 (.A(resetn),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(s_clk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(s_data),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(SelfWriteData[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(SelfWriteData[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(SelfWriteData[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(SelfWriteData[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(SelfWriteData[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(SelfWriteData[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_16 load_slew111 (.A(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_16 load_slew112 (.A(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net112));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[6]));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[7]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[8]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[9]));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LongFrameStrobe));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ReceiveLED));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(RowSelect[0]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(RowSelect[1]));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(RowSelect[2]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(RowSelect[3]));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(RowSelect[4]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ComActive));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[0]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[10]));
 sky130_fd_sc_hd__clkbuf_4 output42 (.A(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[11]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[12]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[13]));
 sky130_fd_sc_hd__clkbuf_4 output45 (.A(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[14]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[15]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[16]));
 sky130_fd_sc_hd__clkbuf_4 output48 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[17]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[18]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[19]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[1]));
 sky130_fd_sc_hd__clkbuf_4 output52 (.A(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[20]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[21]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[22]));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[23]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[24]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[25]));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[26]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[27]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[28]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[29]));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[2]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[30]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[31]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[3]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[4]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[5]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[6]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[7]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[8]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteData[9]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(ConfigWriteStrobe));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[0]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[10]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[11]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[12]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[13]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[14]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[15]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[16]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[17]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[18]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[19]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[1]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[21]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[22]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[23]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[24]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[25]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[26]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[27]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[28]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[29]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[2]));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[30]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[31]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[3]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[4]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameAddressRegister[5]));
endmodule
