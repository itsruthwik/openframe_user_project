* NGSPICE file created from DSP.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt DSP Tile_X0Y0_E1BEG[0] Tile_X0Y0_E1BEG[1] Tile_X0Y0_E1BEG[2] Tile_X0Y0_E1BEG[3]
+ Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3] Tile_X0Y0_E2BEG[0]
+ Tile_X0Y0_E2BEG[1] Tile_X0Y0_E2BEG[2] Tile_X0Y0_E2BEG[3] Tile_X0Y0_E2BEG[4] Tile_X0Y0_E2BEG[5]
+ Tile_X0Y0_E2BEG[6] Tile_X0Y0_E2BEG[7] Tile_X0Y0_E2BEGb[0] Tile_X0Y0_E2BEGb[1] Tile_X0Y0_E2BEGb[2]
+ Tile_X0Y0_E2BEGb[3] Tile_X0Y0_E2BEGb[4] Tile_X0Y0_E2BEGb[5] Tile_X0Y0_E2BEGb[6]
+ Tile_X0Y0_E2BEGb[7] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6BEG[0] Tile_X0Y0_E6BEG[10] Tile_X0Y0_E6BEG[11]
+ Tile_X0Y0_E6BEG[1] Tile_X0Y0_E6BEG[2] Tile_X0Y0_E6BEG[3] Tile_X0Y0_E6BEG[4] Tile_X0Y0_E6BEG[5]
+ Tile_X0Y0_E6BEG[6] Tile_X0Y0_E6BEG[7] Tile_X0Y0_E6BEG[8] Tile_X0Y0_E6BEG[9] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3]
+ Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4BEG[0] Tile_X0Y0_EE4BEG[10] Tile_X0Y0_EE4BEG[11]
+ Tile_X0Y0_EE4BEG[12] Tile_X0Y0_EE4BEG[13] Tile_X0Y0_EE4BEG[14] Tile_X0Y0_EE4BEG[15]
+ Tile_X0Y0_EE4BEG[1] Tile_X0Y0_EE4BEG[2] Tile_X0Y0_EE4BEG[3] Tile_X0Y0_EE4BEG[4]
+ Tile_X0Y0_EE4BEG[5] Tile_X0Y0_EE4BEG[6] Tile_X0Y0_EE4BEG[7] Tile_X0Y0_EE4BEG[8]
+ Tile_X0Y0_EE4BEG[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_NN4BEG[0] Tile_X0Y0_NN4BEG[10] Tile_X0Y0_NN4BEG[11]
+ Tile_X0Y0_NN4BEG[12] Tile_X0Y0_NN4BEG[13] Tile_X0Y0_NN4BEG[14] Tile_X0Y0_NN4BEG[15]
+ Tile_X0Y0_NN4BEG[1] Tile_X0Y0_NN4BEG[2] Tile_X0Y0_NN4BEG[3] Tile_X0Y0_NN4BEG[4]
+ Tile_X0Y0_NN4BEG[5] Tile_X0Y0_NN4BEG[6] Tile_X0Y0_NN4BEG[7] Tile_X0Y0_NN4BEG[8]
+ Tile_X0Y0_NN4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3]
+ Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4]
+ Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1]
+ Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6]
+ Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12]
+ Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7]
+ Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_SS4END[0] Tile_X0Y0_SS4END[10] Tile_X0Y0_SS4END[11]
+ Tile_X0Y0_SS4END[12] Tile_X0Y0_SS4END[13] Tile_X0Y0_SS4END[14] Tile_X0Y0_SS4END[15]
+ Tile_X0Y0_SS4END[1] Tile_X0Y0_SS4END[2] Tile_X0Y0_SS4END[3] Tile_X0Y0_SS4END[4]
+ Tile_X0Y0_SS4END[5] Tile_X0Y0_SS4END[6] Tile_X0Y0_SS4END[7] Tile_X0Y0_SS4END[8]
+ Tile_X0Y0_SS4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[1] Tile_X0Y0_W1END[2] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4]
+ Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1]
+ Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5]
+ Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W2END[0] Tile_X0Y0_W2END[1] Tile_X0Y0_W2END[2]
+ Tile_X0Y0_W2END[3] Tile_X0Y0_W2END[4] Tile_X0Y0_W2END[5] Tile_X0Y0_W2END[6] Tile_X0Y0_W2END[7]
+ Tile_X0Y0_W2MID[0] Tile_X0Y0_W2MID[1] Tile_X0Y0_W2MID[2] Tile_X0Y0_W2MID[3] Tile_X0Y0_W2MID[4]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_W2MID[6] Tile_X0Y0_W2MID[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_W6END[0] Tile_X0Y0_W6END[10] Tile_X0Y0_W6END[11] Tile_X0Y0_W6END[1] Tile_X0Y0_W6END[2]
+ Tile_X0Y0_W6END[3] Tile_X0Y0_W6END[4] Tile_X0Y0_W6END[5] Tile_X0Y0_W6END[6] Tile_X0Y0_W6END[7]
+ Tile_X0Y0_W6END[8] Tile_X0Y0_W6END[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11]
+ Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15]
+ Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4]
+ Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8]
+ Tile_X0Y0_WW4BEG[9] Tile_X0Y0_WW4END[0] Tile_X0Y0_WW4END[10] Tile_X0Y0_WW4END[11]
+ Tile_X0Y0_WW4END[12] Tile_X0Y0_WW4END[13] Tile_X0Y0_WW4END[14] Tile_X0Y0_WW4END[15]
+ Tile_X0Y0_WW4END[1] Tile_X0Y0_WW4END[2] Tile_X0Y0_WW4END[3] Tile_X0Y0_WW4END[4]
+ Tile_X0Y0_WW4END[5] Tile_X0Y0_WW4END[6] Tile_X0Y0_WW4END[7] Tile_X0Y0_WW4END[8]
+ Tile_X0Y0_WW4END[9] Tile_X0Y1_E1BEG[0] Tile_X0Y1_E1BEG[1] Tile_X0Y1_E1BEG[2] Tile_X0Y1_E1BEG[3]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2BEG[0]
+ Tile_X0Y1_E2BEG[1] Tile_X0Y1_E2BEG[2] Tile_X0Y1_E2BEG[3] Tile_X0Y1_E2BEG[4] Tile_X0Y1_E2BEG[5]
+ Tile_X0Y1_E2BEG[6] Tile_X0Y1_E2BEG[7] Tile_X0Y1_E2BEGb[0] Tile_X0Y1_E2BEGb[1] Tile_X0Y1_E2BEGb[2]
+ Tile_X0Y1_E2BEGb[3] Tile_X0Y1_E2BEGb[4] Tile_X0Y1_E2BEGb[5] Tile_X0Y1_E2BEGb[6]
+ Tile_X0Y1_E2BEGb[7] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6BEG[0] Tile_X0Y1_E6BEG[10] Tile_X0Y1_E6BEG[11]
+ Tile_X0Y1_E6BEG[1] Tile_X0Y1_E6BEG[2] Tile_X0Y1_E6BEG[3] Tile_X0Y1_E6BEG[4] Tile_X0Y1_E6BEG[5]
+ Tile_X0Y1_E6BEG[6] Tile_X0Y1_E6BEG[7] Tile_X0Y1_E6BEG[8] Tile_X0Y1_E6BEG[9] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3]
+ Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_EE4BEG[0] Tile_X0Y1_EE4BEG[10] Tile_X0Y1_EE4BEG[11]
+ Tile_X0Y1_EE4BEG[12] Tile_X0Y1_EE4BEG[13] Tile_X0Y1_EE4BEG[14] Tile_X0Y1_EE4BEG[15]
+ Tile_X0Y1_EE4BEG[1] Tile_X0Y1_EE4BEG[2] Tile_X0Y1_EE4BEG[3] Tile_X0Y1_EE4BEG[4]
+ Tile_X0Y1_EE4BEG[5] Tile_X0Y1_EE4BEG[6] Tile_X0Y1_EE4BEG[7] Tile_X0Y1_EE4BEG[8]
+ Tile_X0Y1_EE4BEG[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_NN4END[0]
+ Tile_X0Y1_NN4END[10] Tile_X0Y1_NN4END[11] Tile_X0Y1_NN4END[12] Tile_X0Y1_NN4END[13]
+ Tile_X0Y1_NN4END[14] Tile_X0Y1_NN4END[15] Tile_X0Y1_NN4END[1] Tile_X0Y1_NN4END[2]
+ Tile_X0Y1_NN4END[3] Tile_X0Y1_NN4END[4] Tile_X0Y1_NN4END[5] Tile_X0Y1_NN4END[6]
+ Tile_X0Y1_NN4END[7] Tile_X0Y1_NN4END[8] Tile_X0Y1_NN4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1]
+ Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2]
+ Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7]
+ Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_SS4BEG[0] Tile_X0Y1_SS4BEG[10] Tile_X0Y1_SS4BEG[11]
+ Tile_X0Y1_SS4BEG[12] Tile_X0Y1_SS4BEG[13] Tile_X0Y1_SS4BEG[14] Tile_X0Y1_SS4BEG[15]
+ Tile_X0Y1_SS4BEG[1] Tile_X0Y1_SS4BEG[2] Tile_X0Y1_SS4BEG[3] Tile_X0Y1_SS4BEG[4]
+ Tile_X0Y1_SS4BEG[5] Tile_X0Y1_SS4BEG[6] Tile_X0Y1_SS4BEG[7] Tile_X0Y1_SS4BEG[8]
+ Tile_X0Y1_SS4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W1END[0] Tile_X0Y1_W1END[1] Tile_X0Y1_W1END[2] Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4]
+ Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1]
+ Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5]
+ Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W2END[0] Tile_X0Y1_W2END[1] Tile_X0Y1_W2END[2]
+ Tile_X0Y1_W2END[3] Tile_X0Y1_W2END[4] Tile_X0Y1_W2END[5] Tile_X0Y1_W2END[6] Tile_X0Y1_W2END[7]
+ Tile_X0Y1_W2MID[0] Tile_X0Y1_W2MID[1] Tile_X0Y1_W2MID[2] Tile_X0Y1_W2MID[3] Tile_X0Y1_W2MID[4]
+ Tile_X0Y1_W2MID[5] Tile_X0Y1_W2MID[6] Tile_X0Y1_W2MID[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_W6END[0] Tile_X0Y1_W6END[10] Tile_X0Y1_W6END[11] Tile_X0Y1_W6END[1] Tile_X0Y1_W6END[2]
+ Tile_X0Y1_W6END[3] Tile_X0Y1_W6END[4] Tile_X0Y1_W6END[5] Tile_X0Y1_W6END[6] Tile_X0Y1_W6END[7]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_W6END[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11]
+ Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15]
+ Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4]
+ Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8]
+ Tile_X0Y1_WW4BEG[9] Tile_X0Y1_WW4END[0] Tile_X0Y1_WW4END[10] Tile_X0Y1_WW4END[11]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_WW4END[13] Tile_X0Y1_WW4END[14] Tile_X0Y1_WW4END[15]
+ Tile_X0Y1_WW4END[1] Tile_X0Y1_WW4END[2] Tile_X0Y1_WW4END[3] Tile_X0Y1_WW4END[4]
+ Tile_X0Y1_WW4END[5] Tile_X0Y1_WW4END[6] Tile_X0Y1_WW4END[7] Tile_X0Y1_WW4END[8]
+ Tile_X0Y1_WW4END[9] VGND VPWR
Xclkbuf_2_2__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs VGND VGND VPWR
+ VPWR clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_100_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3155_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q VGND VGND VPWR
+ VPWR _0110_ sky130_fd_sc_hd__inv_2
X_2106_ _1106_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__inv_1
XFILLER_94_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3086_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR
+ VPWR _0041_ sky130_fd_sc_hd__inv_2
X_2037_ _1036_ _1037_ _1035_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o21ai_4
XFILLER_62_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3988_ _0886_ _0891_ _0885_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__o21a_1
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2939_ net972 net967 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4609_ net153 net1114 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_163_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4960_ net45 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_1
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4891_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 VGND VGND VPWR VPWR net242
+ sky130_fd_sc_hd__buf_4
X_3911_ _0117_ _0805_ _0817_ _0816_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__a22o_4
X_3842_ _0543_ net665 VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__or2_4
X_3773_ net58 net60 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q VGND
+ VGND VPWR VPWR _0691_ sky130_fd_sc_hd__mux2_1
X_2724_ _1647_ _1648_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 sky130_fd_sc_hd__mux2_1
XFILLER_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2655_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7
+ _1606_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR
+ VPWR _1607_ sky130_fd_sc_hd__a211o_1
XFILLER_145_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput401 net401 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[1] sky130_fd_sc_hd__buf_2
XFILLER_172_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput412 net412 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput423 net423 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput434 net434 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[8] sky130_fd_sc_hd__buf_2
X_2586_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[17\] net1064 VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__mux2_4
X_4325_ net1254 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput445 net445 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput478 net478 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput456 net456 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput467 net467 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput489 net489 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[14] sky130_fd_sc_hd__buf_2
X_4256_ net52 net1092 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3207_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q _0161_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__a21bo_1
X_4187_ net1253 net1108 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3138_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR
+ VPWR _0093_ sky130_fd_sc_hd__inv_2
XFILLER_103_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3069_ net186 VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__inv_2
XFILLER_42_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_124_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_177_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2440_ net203 net125 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__mux2_1
XFILLER_52_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2371_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q _1349_ _1351_
+ _1353_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__o22a_1
X_4110_ net1239 net1126 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_150_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5090_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 VGND VGND VPWR VPWR net441
+ sky130_fd_sc_hd__buf_1
X_4041_ net1232 net1143 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_142_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4943_ net1252 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__buf_2
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4874_ net1179 net1148 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_50_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_151_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3825_ _0737_ _0736_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3756_ _0674_ _0673_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A2 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_154_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2707_ net1255 net98 net86 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q VGND VGND VPWR VPWR
+ _1644_ sky130_fd_sc_hd__mux4_1
XFILLER_145_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3687_ net100 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__mux2_1
X_2638_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q _1587_ _1591_
+ _1581_ _1583_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7
+ sky130_fd_sc_hd__o32a_1
XFILLER_160_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput253 net253 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput242 net242 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[3] sky130_fd_sc_hd__buf_2
X_2569_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q _1526_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__a21bo_1
Xoutput286 net286 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[12] sky130_fd_sc_hd__buf_2
XFILLER_160_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput264 net264 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput275 net275 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_133_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput297 net297 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[22] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_160_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4308_ net35 net1076 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_141_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4239_ net41 net1091 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1940_ _0922_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q _0939_
+ _0942_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B1 sky130_fd_sc_hd__a22o_4
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3610_ net189 net65 net23 net101 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q VGND VGND VPWR VPWR
+ _0540_ sky130_fd_sc_hd__mux4_2
XFILLER_119_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4590_ net1183 net1120 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_12_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3541_ net1009 net1024 net723 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0476_ sky130_fd_sc_hd__mux4_2
XFILLER_142_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3472_ _0020_ net69 VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__nor2_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5211_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net553
+ sky130_fd_sc_hd__buf_4
X_2423_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q _1392_ _1402_
+ _1396_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C3 sky130_fd_sc_hd__a22o_4
XFILLER_142_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5142_ net1179 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__clkbuf_2
X_2354_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q _1337_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__o21ai_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5073_ Tile_X0Y0_WW4END[8] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_2
X_2285_ _1271_ _1194_ _1272_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__nor3_2
X_4024_ net1250 net1178 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4926_ Tile_X0Y0_EE4END[14] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4857_ net1195 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3808_ _0712_ _0713_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q
+ _0721_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q VGND VGND VPWR
+ VPWR _0722_ sky130_fd_sc_hd__a221o_1
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4788_ net1186 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3739_ _0653_ _0658_ net1061 _0636_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__a211o_4
XFILLER_109_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1220 net95 VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__buf_4
Xfanout1231 net46 VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__buf_4
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1242 net39 VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__buf_4
Xfanout1253 net28 VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__buf_4
XFILLER_78_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2070_ _1065_ _1066_ _1060_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__a21bo_1
XFILLER_93_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2972_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q _1840_ _1842_
+ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1923_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q _0926_ _0123_
+ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__a21o_1
X_4711_ net148 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4642_ net1205 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4573_ net158 net1122 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_151_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3524_ net1010 net724 net1025 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0459_ sky130_fd_sc_hd__mux4_1
X_3455_ net7 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q VGND VGND
+ VPWR VPWR _0396_ sky130_fd_sc_hd__nand2b_1
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2406_ _1079_ _1086_ _1085_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__a21o_1
XFILLER_130_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3386_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0332_ VGND VGND
+ VPWR VPWR _0333_ sky130_fd_sc_hd__nand2_1
XFILLER_69_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2337_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\] _1320_ net1057 VGND VGND VPWR VPWR
+ _1321_ sky130_fd_sc_hd__mux2_4
XFILLER_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5125_ Tile_X0Y1_EE4END[12] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkbuf_1
X_5056_ net112 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__buf_1
XFILLER_84_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2268_ net978 net997 net1019 net1014 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR
+ _1258_ sky130_fd_sc_hd__mux4_1
XFILLER_29_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4007_ net1229 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2199_ _1190_ _1191_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_83_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4909_ Tile_X0Y0_E6END[7] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3240_ _0187_ _0189_ _0192_ _0026_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q
+ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a221o_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3171_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q VGND VGND VPWR
+ VPWR _0126_ sky130_fd_sc_hd__inv_1
X_2122_ _0089_ _1122_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__or2_1
Xfanout1050 net1052 VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__buf_2
Xfanout1083 net1085 VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__clkbuf_2
Xfanout1072 net1077 VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__buf_2
XFILLER_86_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1061 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q VGND VGND
+ VPWR VPWR net1061 sky130_fd_sc_hd__buf_4
XFILLER_66_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1094 net1095 VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2053_ _1040_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__and2b_1
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2955_ net747 net733 net693 net709 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q VGND VGND VPWR VPWR
+ _1828_ sky130_fd_sc_hd__mux4_1
XFILLER_175_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1906_ _0740_ _0829_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__nor2_1
Xrebuffer118 Tile_X0Y1_DSP_bot.A0 VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer129 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 VGND VGND VPWR VPWR net746
+ sky130_fd_sc_hd__dlygate4sd1_1
X_2886_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 _1327_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q
+ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4625_ net1190 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4556_ net1181 net1129 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3507_ net76 net112 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q VGND
+ VGND VPWR VPWR _0444_ sky130_fd_sc_hd__mux2_1
XFILLER_143_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4487_ net1211 net1173 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_106_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3438_ _0376_ _0046_ _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__o21ai_4
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3369_ _0314_ _0315_ _0316_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q VGND VGND VPWR VPWR
+ _0317_ sky130_fd_sc_hd__a221o_1
XFILLER_66_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5108_ Tile_X0Y1_E6END[5] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_2
XFILLER_57_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5039_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 VGND VGND VPWR VPWR net390
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput120 Tile_X0Y1_E1END[1] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_4
Xinput153 Tile_X0Y1_FrameData[18] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_2
Xinput131 Tile_X0Y1_E2MID[0] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xinput142 Tile_X0Y1_EE4END[1] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput164 Tile_X0Y1_FrameData[29] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_4
Xinput175 Tile_X0Y1_N1END[2] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_4
Xinput186 Tile_X0Y1_N2MID[1] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_4
XFILLER_56_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput197 Tile_X0Y1_N4END[4] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_4
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2740_ net740 _0704_ _0733_ _0253_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _1661_ sky130_fd_sc_hd__mux4_1
XFILLER_82_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2671_ net1012 net1048 net1027 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR
+ _1617_ sky130_fd_sc_hd__mux4_1
XFILLER_157_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4410_ net1252 net1152 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_117_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput605 net605 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[14] sky130_fd_sc_hd__buf_4
XFILLER_172_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4341_ net1247 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_125_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4272_ net40 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3223_ net971 net727 net707 net977 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0177_ sky130_fd_sc_hd__mux4_2
XFILLER_140_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3154_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q VGND VGND VPWR
+ VPWR _0109_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_19_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2105_ _0845_ _0848_ _1104_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__nor3b_1
X_3085_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q VGND VGND VPWR
+ VPWR _0040_ sky130_fd_sc_hd__inv_2
X_2036_ _1034_ _1033_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__xnor2_4
XFILLER_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3987_ _0887_ _0890_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2938_ net1217 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_157_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2869_ _1760_ _1761_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 sky130_fd_sc_hd__mux2_1
XFILLER_163_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4608_ net154 net1114 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4539_ net1197 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4890_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 VGND VGND VPWR VPWR net241
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_83_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3910_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q VGND VGND VPWR VPWR
+ _0817_ sky130_fd_sc_hd__o21a_1
XFILLER_149_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3841_ _0752_ _0750_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__nor2_4
X_3772_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q _0689_ _0687_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q VGND VGND VPWR VPWR
+ _0690_ sky130_fd_sc_hd__a211o_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2723_ net1006 _0704_ _0733_ _1498_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR
+ _1648_ sky130_fd_sc_hd__mux4_1
XFILLER_157_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2654_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q _1186_ VGND VGND
+ VPWR VPWR _1606_ sky130_fd_sc_hd__nor2_1
XFILLER_145_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput402 net402 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[2] sky130_fd_sc_hd__buf_2
XFILLER_160_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput413 net413 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput424 net424 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[13] sky130_fd_sc_hd__buf_6
Xoutput435 net435 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[9] sky130_fd_sc_hd__buf_2
X_2585_ _1541_ _1523_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ sky130_fd_sc_hd__mux2_4
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4324_ net1243 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput446 net446 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[6] sky130_fd_sc_hd__buf_8
Xoutput468 net468 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput457 net457 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[10] sky130_fd_sc_hd__buf_2
Xoutput479 net479 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[5] sky130_fd_sc_hd__buf_2
X_4255_ net1224 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3206_ net1036 net1006 net1031 net1054 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0161_ sky130_fd_sc_hd__mux4_1
X_4186_ net1252 net1108 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3137_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q VGND VGND VPWR
+ VPWR _0092_ sky130_fd_sc_hd__inv_2
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3068_ net189 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__inv_1
XFILLER_179_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2019_ _0995_ _1018_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_177_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2370_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q _1352_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__a21bo_1
XFILLER_110_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4040_ net1231 net1143 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4942_ net1253 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4873_ net1213 net1153 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_50_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3824_ net205 net63 net7 net99 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q VGND VGND VPWR VPWR
+ _0737_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_15_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3755_ _0662_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q _0663_
+ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__o21ai_2
X_2706_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q _1640_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_154_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3686_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q _0610_ VGND VGND
+ VPWR VPWR _0611_ sky130_fd_sc_hd__and2b_1
X_2637_ _0142_ _1590_ _1589_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q
+ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__o211a_1
XFILLER_145_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput243 net243 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[4] sky130_fd_sc_hd__buf_2
X_2568_ net1042 net1033 net1037 net1021 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q VGND VGND VPWR VPWR
+ _1526_ sky130_fd_sc_hd__mux4_1
XFILLER_160_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput265 net265 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput276 net276 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput254 net254 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput298 net298 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput287 net287 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[13] sky130_fd_sc_hd__buf_2
XFILLER_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4307_ net1245 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2499_ _1469_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 sky130_fd_sc_hd__mux2_4
X_4238_ net42 net1091 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4169_ net1232 net1108 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3540_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0458_ _0470_
+ _0472_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__o32a_1
XFILLER_127_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5210_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR net567
+ sky130_fd_sc_hd__buf_6
X_3471_ _0399_ _0406_ _0409_ _0020_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__o211a_1
XFILLER_89_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2422_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q _1401_ VGND VGND
+ VPWR VPWR _1402_ sky130_fd_sc_hd__nor2_1
XFILLER_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5141_ net1180 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__clkbuf_2
X_2353_ _1336_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__inv_1
X_5072_ Tile_X0Y0_WW4END[7] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__buf_2
X_4023_ net1249 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2284_ _1094_ _0994_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__xor2_1
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4925_ Tile_X0Y0_EE4END[13] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4856_ net1193 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3807_ net111 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__mux2_1
X_1999_ _0784_ _0575_ _0574_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__and3_4
XFILLER_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4787_ net1214 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3738_ _0653_ _0658_ _0636_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X
+ sky130_fd_sc_hd__a21o_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3669_ _0594_ _0595_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q
+ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__mux2_1
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1232 net45 VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__clkbuf_4
Xfanout1221 net56 VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__buf_4
XFILLER_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1210 net149 VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1254 net27 VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__buf_4
Xfanout1243 net38 VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__buf_4
XFILLER_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2971_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q _0662_ _1841_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q VGND VGND VPWR VPWR
+ _1842_ sky130_fd_sc_hd__a211o_1
XFILLER_91_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1922_ net1019 net1015 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__mux2_1
X_4710_ net1210 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4641_ net1204 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4572_ net159 net1122 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3523_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q _0457_ VGND VGND
+ VPWR VPWR _0458_ sky130_fd_sc_hd__and2b_1
X_3454_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q net104 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q
+ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__o21ai_2
XFILLER_6_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2405_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\] _1384_ net1057 VGND VGND VPWR VPWR
+ _1385_ sky130_fd_sc_hd__mux2_1
XFILLER_130_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3385_ net100 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux2_1
XFILLER_69_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2336_ Tile_X0Y1_DSP_bot.C8 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[8\] net1063 VGND
+ VGND VPWR VPWR _1320_ sky130_fd_sc_hd__mux2_2
XFILLER_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5124_ Tile_X0Y1_EE4END[11] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkbuf_1
X_5055_ net111 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__buf_1
X_2267_ net973 net968 net987 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR
+ _1257_ sky130_fd_sc_hd__mux4_1
XFILLER_84_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4006_ net1228 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2198_ _1191_ _1190_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_83_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4908_ Tile_X0Y0_E6END[6] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4839_ net148 net1157 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_153_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_180_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1040 net1041 VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__buf_6
X_3170_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q VGND VGND VPWR
+ VPWR _0125_ sky130_fd_sc_hd__inv_2
X_2121_ _1120_ _1121_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q
+ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__mux2_1
Xfanout1051 net1052 VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__buf_2
Xfanout1073 net1074 VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__buf_2
XFILLER_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1062 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q VGND VGND
+ VPWR VPWR net1062 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1084 net1085 VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__buf_2
XFILLER_120_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2052_ _1041_ _1049_ _1052_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__a21o_1
Xfanout1095 net1096 VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2954_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q _1824_ _1826_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q VGND VGND VPWR VPWR
+ _1827_ sky130_fd_sc_hd__o211a_1
XFILLER_175_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer108 _0174_ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_20_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2885_ net1017 net1003 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q
+ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__mux2_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4624_ net1185 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4555_ net171 net1129 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_128_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3506_ _0425_ _0044_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q
+ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__mux2_1
XFILLER_143_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4486_ net1210 net1173 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_103_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3437_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q _0379_ VGND VGND
+ VPWR VPWR _0380_ sky130_fd_sc_hd__or2_1
X_3368_ net988 net993 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2319_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q _0557_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q
+ _1304_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__a211o_1
X_5107_ Tile_X0Y1_E6END[4] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__buf_1
XFILLER_181_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3299_ net94 net1219 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
XFILLER_111_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5038_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 VGND VGND VPWR VPWR net389
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput110 Tile_X0Y0_W2MID[5] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput154 Tile_X0Y1_FrameData[19] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_2
Xinput121 Tile_X0Y1_E1END[2] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
Xinput132 Tile_X0Y1_E2MID[1] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput143 Tile_X0Y1_EE4END[2] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
Xinput165 Tile_X0Y1_FrameData[2] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
Xinput187 Tile_X0Y1_N2MID[2] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_4
Xinput176 Tile_X0Y1_N1END[3] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput198 Tile_X0Y1_N4END[5] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_4
XFILLER_63_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2670_ _1616_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 sky130_fd_sc_hd__mux2_4
XFILLER_75_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput606 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR
+ Tile_X0Y1_WW4BEG[15] sky130_fd_sc_hd__buf_6
X_4340_ net1246 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4271_ net1240 net1084 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_125_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3222_ _0031_ _0175_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__nor2_2
XFILLER_100_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3153_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR
+ VPWR _0108_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2104_ _0845_ _0848_ _1104_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__o21ba_4
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3084_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q VGND VGND VPWR
+ VPWR _0039_ sky130_fd_sc_hd__inv_2
X_2035_ _1029_ _1030_ _1031_ _1023_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3986_ _0832_ _0888_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2937_ net212 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q VGND
+ VGND VPWR VPWR _1811_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_157_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4607_ net1201 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2868_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 _1327_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q
+ VGND VGND VPWR VPWR _1761_ sky130_fd_sc_hd__mux2_1
XFILLER_163_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2799_ _0243_ net94 net2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q VGND VGND VPWR VPWR
+ _1711_ sky130_fd_sc_hd__mux4_1
XFILLER_116_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4538_ net1196 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_171_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4469_ net1188 net1173 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3840_ _0580_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__nand2_1
X_3771_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__inv_1
X_2722_ net619 net1258 net1220 net1026 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q VGND VGND VPWR VPWR
+ _1647_ sky130_fd_sc_hd__mux4_1
XFILLER_145_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2653_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q _1601_ _1605_
+ _1595_ _1597_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7
+ sky130_fd_sc_hd__o32a_1
XFILLER_145_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput414 net414 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput425 net425 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput403 net403 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[3] sky130_fd_sc_hd__buf_2
X_2584_ _1536_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q _1538_
+ _1540_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__o22a_1
XFILLER_153_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4323_ net1230 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput458 net458 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[11] sky130_fd_sc_hd__buf_6
Xoutput436 net436 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput447 net447 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[7] sky130_fd_sc_hd__buf_6
Xoutput469 net469 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[10] sky130_fd_sc_hd__buf_2
XFILLER_113_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4254_ net1223 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3205_ _0085_ _0159_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__and2_1
X_4185_ net1251 net1110 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3136_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR
+ VPWR _0091_ sky130_fd_sc_hd__inv_2
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3067_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q VGND VGND VPWR
+ VPWR _0022_ sky130_fd_sc_hd__inv_2
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2018_ _1018_ _0995_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__and2b_1
XFILLER_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3969_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q _0870_ _0874_
+ _0865_ _0866_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6
+ sky130_fd_sc_hd__o32a_4
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4941_ net1221 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_2
XFILLER_177_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4872_ net1212 net1153 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3823_ net25 net79 net104 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q VGND VGND VPWR VPWR
+ _0736_ sky130_fd_sc_hd__mux4_1
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3754_ _0672_ _0671_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__mux2_4
X_2705_ _0068_ _1641_ VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_154_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3685_ net64 net80 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q VGND
+ VGND VPWR VPWR _0610_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2636_ net85 net115 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__mux2_1
XFILLER_133_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput244 net244 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[5] sky130_fd_sc_hd__buf_6
XFILLER_133_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2567_ _0098_ _1524_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__and2_1
XFILLER_160_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput266 net266 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[9] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput255 net255 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput277 net277 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput299 net299 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput288 net288 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[14] sky130_fd_sc_hd__buf_2
X_4306_ net1244 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2498_ _1450_ _1370_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__xor2_1
XFILLER_59_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4237_ net1238 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4168_ net46 net1108 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_74_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4099_ net1230 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3119_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q VGND VGND VPWR
+ VPWR _0074_ sky130_fd_sc_hd__inv_2
XFILLER_130_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap616 _1273_ VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__clkbuf_2
XFILLER_182_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3470_ _0399_ _0406_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__o21ai_4
X_2421_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q _1400_ _1398_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q VGND VGND VPWR VPWR
+ _1401_ sky130_fd_sc_hd__o211a_1
XFILLER_142_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5140_ net1181 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__buf_4
X_2352_ net186 net132 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__mux2_1
XFILLER_150_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5071_ Tile_X0Y0_WW4END[6] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkbuf_2
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2283_ net1063 Tile_X0Y1_DSP_bot.C9 _1270_ net1057 VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__o211a_1
X_4022_ net1248 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4924_ Tile_X0Y0_EE4END[12] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4855_ net1192 net1148 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3806_ _0717_ _0715_ _0720_ _0067_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3
+ sky130_fd_sc_hd__a22o_4
X_4786_ net1202 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_109_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3737_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q _0657_ _0655_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q VGND VGND VPWR VPWR
+ _0658_ sky130_fd_sc_hd__a31oi_4
X_1998_ _0677_ _0575_ _0574_ _0998_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__a31oi_4
XFILLER_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3668_ net71 net215 net83 net229 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q VGND VGND VPWR VPWR
+ _0595_ sky130_fd_sc_hd__mux4_1
X_2619_ net1012 net1048 net1027 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR
+ _1573_ sky130_fd_sc_hd__mux4_1
XFILLER_121_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3599_ _0528_ _0527_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ _0522_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__a211o_1
XFILLER_114_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1222 net55 VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__clkbuf_4
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1200 net157 VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__buf_4
XFILLER_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1211 net148 VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__buf_4
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1233 net1234 VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__buf_4
Xfanout1255 net22 VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__clkbuf_4
Xfanout1244 net37 VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_77_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2970_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q net734 VGND
+ VGND VPWR VPWR _1841_ sky130_fd_sc_hd__nor2_1
X_1921_ _0121_ net998 _0924_ _0122_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__o211a_1
XFILLER_42_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4640_ net1203 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4571_ net1197 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3522_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 net13 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q
+ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_139_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3453_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q _0329_ _0334_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q _0338_ VGND VGND VPWR
+ VPWR _0394_ sky130_fd_sc_hd__o311a_4
XFILLER_170_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2404_ Tile_X0Y1_DSP_bot.C4 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[4\] net1063 VGND
+ VGND VPWR VPWR _1384_ sky130_fd_sc_hd__mux2_1
XFILLER_130_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3384_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__inv_1
X_5123_ Tile_X0Y1_EE4END[10] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__buf_1
X_2335_ _1306_ _1303_ _1319_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C8 sky130_fd_sc_hd__o22a_4
XFILLER_69_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5054_ net110 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__buf_1
XFILLER_84_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2266_ _0127_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 VGND VGND VPWR
+ VPWR _1256_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_162_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2197_ _0954_ _1095_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__xnor2_1
X_4005_ _0906_ _0907_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__xor2_1
XFILLER_84_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_148_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4907_ Tile_X0Y0_E6END[5] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4838_ net149 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_138_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4769_ net1204 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_157_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1030 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 VGND VGND VPWR VPWR
+ net1030 sky130_fd_sc_hd__buf_2
X_2120_ net1042 net1033 net1007 net1054 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q VGND VGND VPWR VPWR
+ _1121_ sky130_fd_sc_hd__mux4_1
Xfanout1052 net1053 VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__buf_2
Xfanout1041 net1044 VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__buf_8
XFILLER_120_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1074 net1077 VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__buf_1
Xfanout1063 net1064 VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1085 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__clkbuf_2
Xfanout1096 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__clkbuf_2
X_2051_ _1051_ _1050_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__and2b_1
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2953_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q _1825_ VGND
+ VGND VPWR VPWR _1826_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2884_ net995 _0216_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 _0230_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_30_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer109 net746 VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__clkbuf_2
XFILLER_175_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4623_ net1184 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_175_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4554_ net172 net1129 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3505_ _0441_ _0440_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q
+ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux2_1
XFILLER_143_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4485_ net1209 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3436_ _0377_ _0378_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q
+ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux2_1
X_3367_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q net974 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__o21ba_1
X_2318_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4
+ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__nor2_1
X_5106_ Tile_X0Y1_E6END[3] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__buf_1
X_3298_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q _0248_ VGND VGND
+ VPWR VPWR _0249_ sky130_fd_sc_hd__or2_1
X_5037_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net388
+ sky130_fd_sc_hd__buf_1
XFILLER_174_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2249_ _1238_ _1239_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q
+ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__mux2_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput100 Tile_X0Y0_W2END[3] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_2
Xinput111 Tile_X0Y0_W2MID[6] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
XFILLER_163_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput122 Tile_X0Y1_E1END[3] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_1
Xinput133 Tile_X0Y1_E2MID[2] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xinput144 Tile_X0Y1_EE4END[3] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_1
XFILLER_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput155 Tile_X0Y1_FrameData[1] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xinput166 Tile_X0Y1_FrameData[3] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_2
Xinput177 Tile_X0Y1_N2END[0] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput199 Tile_X0Y1_N4END[6] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_4
Xinput188 Tile_X0Y1_N2MID[3] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput607 net607 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_125_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4270_ net1239 net1084 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3221_ net981 net995 net1017 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0175_ sky130_fd_sc_hd__mux4_2
XFILLER_140_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3152_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q VGND VGND VPWR
+ VPWR _0107_ sky130_fd_sc_hd__inv_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2103_ _1103_ _0661_ net722 _1102_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__o31ai_2
X_3083_ net228 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
XFILLER_94_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2034_ _1033_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__nand2_4
XFILLER_54_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3985_ _0576_ _0729_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__nor2_1
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2936_ _1806_ _1809_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q
+ _1810_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3
+ sky130_fd_sc_hd__o22a_4
XFILLER_148_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2867_ net747 _1361_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q
+ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__mux2_1
XFILLER_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4606_ net1200 net1114 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_163_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2798_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q _1709_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__a21bo_1
XFILLER_89_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4537_ net1195 net1131 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4468_ net1186 net1173 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3419_ net981 net996 net1016 net1015 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0363_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_168_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4399_ net1240 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3770_ net2 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q VGND
+ VGND VPWR VPWR _0688_ sky130_fd_sc_hd__mux2_1
X_2721_ net708 _0322_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 _0346_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2652_ _0140_ _1604_ _1603_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q
+ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__o211a_1
XFILLER_160_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput415 net415 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput426 net426 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[15] sky130_fd_sc_hd__buf_6
Xoutput404 net404 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[4] sky130_fd_sc_hd__buf_2
X_2583_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q _1539_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q
+ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__a21bo_1
XFILLER_160_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_112_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4322_ net1227 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput437 net437 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput448 net448 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput459 net459 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[1] sky130_fd_sc_hd__buf_2
X_4253_ net1222 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3204_ net1011 net1046 net1026 net1050 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0159_ sky130_fd_sc_hd__mux4_1
X_4184_ net1250 net1110 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3135_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q VGND VGND VPWR
+ VPWR _0090_ sky130_fd_sc_hd__inv_1
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3066_ net139 VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__inv_1
X_2017_ _1016_ _1017_ _1015_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_53_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3968_ _0095_ _0873_ _0872_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q
+ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__o211a_1
XFILLER_10_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2919_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q _0662_ _1795_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _1796_ sky130_fd_sc_hd__a211o_1
XFILLER_148_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3899_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q _0806_ VGND VGND
+ VPWR VPWR _0807_ sky130_fd_sc_hd__or2_4
XFILLER_128_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_177_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4940_ net1222 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4871_ net1211 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3822_ _0734_ _0733_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3753_ net181 net73 net141 net217 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q VGND VGND VPWR VPWR
+ _0672_ sky130_fd_sc_hd__mux4_2
X_2704_ net1036 net1006 net1031 net1054 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _1641_ sky130_fd_sc_hd__mux4_1
X_3684_ _0606_ _0607_ _0608_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR VPWR
+ _0609_ sky130_fd_sc_hd__a221o_1
X_2635_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q _1588_ VGND VGND
+ VPWR VPWR _1589_ sky130_fd_sc_hd__or2_1
XFILLER_145_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_120_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2566_ net1011 net1047 net1026 net1052 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR
+ _1524_ sky130_fd_sc_hd__mux4_1
X_4305_ net1242 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_160_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput256 net256 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[10] sky130_fd_sc_hd__buf_2
Xoutput267 net267 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_126_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput289 net289 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput278 net278 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_141_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2497_ _1468_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 sky130_fd_sc_hd__mux2_4
X_4236_ net1237 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4167_ net1229 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3118_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q VGND VGND VPWR
+ VPWR _0073_ sky130_fd_sc_hd__inv_2
XFILLER_67_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4098_ net1227 net1133 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3049_ net963 _1467_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__and2b_1
XFILLER_90_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2420_ _1399_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__inv_1
XFILLER_89_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2351_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net222 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__mux2_4
X_5070_ Tile_X0Y0_WW4END[5] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkbuf_2
X_2282_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[9\] net1064 VGND VGND VPWR VPWR _1270_
+ sky130_fd_sc_hd__nand2b_1
X_4021_ net1247 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4923_ Tile_X0Y0_EE4END[11] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4854_ net1191 net1148 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_165_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3805_ _0718_ _0719_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q
+ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__mux2_1
X_1997_ _0450_ _0785_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__nor2_1
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4785_ net1190 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_158_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3736_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q _0656_ VGND VGND
+ VPWR VPWR _0657_ sky130_fd_sc_hd__nand2_1
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3667_ net173 net179 net125 net1216 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0594_ sky130_fd_sc_hd__mux4_1
X_2618_ _0145_ _1571_ _1570_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q
+ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__o211a_1
XFILLER_133_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3598_ _0527_ _0528_ _0522_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__a21o_4
X_2549_ net206 net66 net10 net102 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q VGND VGND VPWR VPWR
+ _1509_ sky130_fd_sc_hd__mux4_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4219_ net28 net1100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_85_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5199_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net541
+ sky130_fd_sc_hd__buf_1
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1223 net54 VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__buf_4
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1201 net156 VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__buf_4
Xfanout1212 net147 VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__buf_4
Xfanout1234 Tile_X0Y0_FrameData[27] VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__clkbuf_2
Xfanout1245 net36 VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__clkbuf_4
Xfanout1256 net21 VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__buf_2
XFILLER_78_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1920_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q net983 VGND VGND
+ VPWR VPWR _0924_ sky130_fd_sc_hd__or2_1
X_4570_ net1196 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_155_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3521_ _0456_ _0453_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 sky130_fd_sc_hd__mux2_4
X_3452_ _0357_ _0358_ _0392_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q VGND VGND VPWR VPWR
+ _0393_ sky130_fd_sc_hd__a221o_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3383_ net1255 net64 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__mux2_1
XFILLER_103_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2403_ _1374_ _1380_ _1383_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C4 sky130_fd_sc_hd__a22o_1
XFILLER_111_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2334_ _1307_ _1318_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q
+ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__mux2_1
XFILLER_69_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5122_ Tile_X0Y1_EE4END[9] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_110_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5053_ net109 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__buf_1
XFILLER_84_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2265_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q _1253_ _1255_
+ _1248_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7
+ sky130_fd_sc_hd__o31ai_2
XTAP_TAPCELL_ROW_162_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2196_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\] _1189_ net1058 VGND VGND VPWR VPWR
+ _1190_ sky130_fd_sc_hd__mux2_4
X_4004_ _0906_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__nor2_1
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4906_ Tile_X0Y0_E6END[4] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4837_ net1209 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_153_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4768_ net1203 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3719_ _0243_ net190 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux2_2
X_4699_ net160 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_136_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_180_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1031 net1033 VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__buf_2
Xfanout1020 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 VGND VGND VPWR VPWR net1020
+ sky130_fd_sc_hd__buf_12
Xfanout1042 net1044 VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__buf_2
Xfanout1053 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 VGND VGND VPWR VPWR
+ net1053 sky130_fd_sc_hd__buf_8
Xfanout1064 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q VGND VGND
+ VPWR VPWR net1064 sky130_fd_sc_hd__buf_4
XFILLER_86_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1075 net1076 VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__clkbuf_2
X_2050_ _1049_ _1041_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__xnor2_2
Xfanout1097 net1098 VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__clkbuf_2
Xfanout1086 net1089 VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__buf_2
XFILLER_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_179_Right_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2952_ _1410_ _1349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__mux2_1
XFILLER_175_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2883_ _1763_ _1765_ _1768_ _0153_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4622_ net1183 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4553_ net146 net1129 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3504_ net208 net67 net11 net103 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q VGND VGND VPWR VPWR
+ _0441_ sky130_fd_sc_hd__mux4_1
XFILLER_128_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4484_ net1208 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3435_ net72 net216 net84 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q VGND VGND VPWR VPWR
+ _0378_ sky130_fd_sc_hd__mux4_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3366_ _0055_ net968 VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__or2_1
X_3297_ net58 net66 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q VGND
+ VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
XFILLER_111_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2317_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6
+ _1302_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q VGND VGND VPWR
+ VPWR _1303_ sky130_fd_sc_hd__o211a_1
X_5105_ Tile_X0Y1_E6END[2] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5036_ clknet_1_0__leaf_Tile_X0Y1_UserCLK VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__buf_2
X_2248_ net979 net998 net984 net1002 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q VGND VGND VPWR VPWR
+ _1239_ sky130_fd_sc_hd__mux4_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2179_ net200 net8 net100 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q VGND VGND VPWR VPWR
+ _1175_ sky130_fd_sc_hd__mux4_2
XFILLER_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput101 Tile_X0Y0_W2END[4] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_4
Xinput112 Tile_X0Y0_W2MID[7] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput145 Tile_X0Y1_FrameData[0] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput134 Tile_X0Y1_E2MID[3] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput123 Tile_X0Y1_E2END[0] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_1
Xinput156 Tile_X0Y1_FrameData[20] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_2
Xinput167 Tile_X0Y1_FrameData[4] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_2
Xinput178 Tile_X0Y1_N2END[1] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 Tile_X0Y1_N2MID[4] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_4
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput608 net608 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_125_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_176_Left_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3220_ _0170_ _0171_ _0172_ _0035_ _0029_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a221o_1
XFILLER_100_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3151_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q VGND VGND VPWR
+ VPWR _0106_ sky130_fd_sc_hd__inv_2
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2102_ _0492_ _0620_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__or2_1
X_3082_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR
+ VPWR _0037_ sky130_fd_sc_hd__inv_2
X_2033_ _1011_ _1006_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__xor2_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3984_ _0450_ _0729_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__nor2_1
XFILLER_148_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2935_ net174 net120 _0529_ net984 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _1810_ sky130_fd_sc_hd__mux4_2
XFILLER_148_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2866_ net715 _0216_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 _0230_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_157_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4605_ net1199 net1114 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2797_ _1512_ _0489_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q
+ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__mux2_1
XFILLER_116_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4536_ net1193 net1131 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_171_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4467_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3418_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q _0361_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a21bo_1
X_4398_ net1239 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_168_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3349_ _0296_ _0297_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q
+ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5019_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net361
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2720_ net695 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net965 _0278_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 sky130_fd_sc_hd__mux4_1
X_2651_ net93 net1220 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__mux2_1
XFILLER_157_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput416 net416 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput405 net405 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[5] sky130_fd_sc_hd__buf_2
X_2582_ net70 net106 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q
+ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__mux2_1
XFILLER_153_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput427 net427 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4321_ net1226 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput438 net438 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput449 net449 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[1] sky130_fd_sc_hd__buf_2
X_4252_ net1221 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3203_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR _0158_
+ sky130_fd_sc_hd__inv_1
X_4183_ net32 net1110 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3134_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q VGND VGND VPWR
+ VPWR _0089_ sky130_fd_sc_hd__inv_1
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3065_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q VGND VGND VPWR
+ VPWR _0020_ sky130_fd_sc_hd__inv_2
X_2016_ _1013_ _1014_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__xnor2_2
XFILLER_35_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3967_ net94 net1219 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__mux2_1
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2918_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q net733 VGND
+ VGND VPWR VPWR _1795_ sky130_fd_sc_hd__nor2_1
XFILLER_163_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3898_ net974 net970 net989 net994 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0806_ sky130_fd_sc_hd__mux4_2
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2849_ net179 net1215 net194 net743 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A sky130_fd_sc_hd__mux4_1
XFILLER_151_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4519_ net1211 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4870_ net1210 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3821_ net15 net107 net71 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q VGND VGND VPWR VPWR
+ _0734_ sky130_fd_sc_hd__mux4_1
XFILLER_177_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3752_ net194 net230 net1215 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q
+ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__mux4_2
X_2703_ net1046 net1026 net1050 net1042 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _1640_ sky130_fd_sc_hd__mux4_1
X_3683_ net8 net1255 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q VGND
+ VGND VPWR VPWR _0608_ sky130_fd_sc_hd__mux2_1
X_2634_ net57 net59 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q VGND
+ VGND VPWR VPWR _1588_ sky130_fd_sc_hd__mux2_1
XFILLER_160_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput235 net235 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[0] sky130_fd_sc_hd__buf_2
X_2565_ _1522_ _0278_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q
+ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__mux2_1
XFILLER_99_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4304_ net1241 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_160_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput257 net257 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[11] sky130_fd_sc_hd__buf_6
Xoutput268 net268 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput246 net246 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_99_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput279 net279 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2496_ _1407_ _1448_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__xor2_1
X_4235_ net1236 net1091 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_165_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4166_ net1228 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3117_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q VGND VGND VPWR
+ VPWR _0072_ sky130_fd_sc_hd__inv_2
XFILLER_67_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4097_ net1226 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3048_ net963 _1468_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__and2b_1
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4999_ net694 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_6
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2350_ _1332_ _1331_ _1333_ _0136_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__a221o_1
XFILLER_96_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2281_ _1242_ _0128_ _1269_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C9 sky130_fd_sc_hd__o21ba_4
X_4020_ net1246 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_8_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4922_ Tile_X0Y0_EE4END[10] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4853_ net1189 net1148 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3804_ net1256 net65 net101 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0719_ sky130_fd_sc_hd__mux4_1
X_1996_ _0601_ _0829_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__nor2_1
X_4784_ net1185 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3735_ net74 net110 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q
+ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__mux2_1
XFILLER_173_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3666_ _0590_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q
+ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_171_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2617_ net61 net93 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q VGND
+ VGND VPWR VPWR _1571_ sky130_fd_sc_hd__mux2_1
X_3597_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q net1035 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q
+ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__o21ba_1
X_2548_ net22 net78 net118 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR
+ _1508_ sky130_fd_sc_hd__mux4_1
XFILLER_141_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4218_ net29 net1100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2479_ _1454_ _1453_ _1324_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__a21o_1
X_5198_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net540
+ sky130_fd_sc_hd__clkbuf_1
X_4149_ net34 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload0 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_4
XFILLER_166_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1202 net155 VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__clkbuf_4
Xfanout1213 net146 VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__buf_4
Xfanout1246 net35 VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__buf_4
Xfanout1224 net53 VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__buf_4
XFILLER_132_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1235 net1236 VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__buf_4
XFILLER_120_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1257 net4 VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_85_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3520_ _0454_ _0455_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q
+ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__mux2_1
XFILLER_170_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3451_ net75 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q
+ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux2_1
XFILLER_6_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3382_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0325_ _0326_
+ _0328_ _0043_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__o311a_4
X_2402_ _1382_ _1381_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__mux2_1
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2333_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q VGND VGND VPWR VPWR
+ _1318_ sky130_fd_sc_hd__mux2_1
X_5121_ Tile_X0Y1_EE4END[8] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_110_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5052_ net108 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_2
X_2264_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q _1254_ VGND VGND
+ VPWR VPWR _1255_ sky130_fd_sc_hd__nor2_1
X_2195_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[10\] net1064 VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__mux2_4
X_4003_ _0881_ _0882_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4905_ Tile_X0Y0_E6END[3] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_1
XFILLER_33_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4836_ net1208 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_23_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1979_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\] net1061 VGND VGND VPWR VPWR _0980_
+ sky130_fd_sc_hd__nand2b_1
X_4767_ net1201 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3718_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q _0639_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a21bo_1
XFILLER_146_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4698_ net161 net1089 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3649_ _0574_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__nand2_1
XFILLER_161_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_89_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1021 net1023 VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__clkbuf_4
Xfanout1010 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 VGND VGND VPWR VPWR
+ net1010 sky130_fd_sc_hd__buf_8
XFILLER_105_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1032 net1033 VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__buf_2
Xfanout1054 net1056 VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__clkbuf_4
Xfanout1043 net1044 VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__buf_2
Xfanout1065 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q VGND VGND
+ VPWR VPWR net1065 sky130_fd_sc_hd__clkbuf_4
Xfanout1076 net1077 VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1098 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__clkbuf_2
Xfanout1087 net1089 VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__buf_2
XFILLER_66_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2951_ _0662_ _0819_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__mux2_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2882_ _1766_ _1767_ _0152_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__mux2_1
X_4621_ net1182 net1112 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4552_ net147 net1129 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3503_ net8 net117 net88 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q VGND VGND VPWR VPWR
+ _0440_ sky130_fd_sc_hd__mux4_1
XFILLER_128_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4483_ net1206 net1174 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3434_ net174 net180 net126 net1215 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0377_ sky130_fd_sc_hd__mux4_1
XFILLER_143_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3365_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q _0312_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q
+ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__a21bo_1
X_3296_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q _0244_ _0246_
+ _0085_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__o211a_1
X_5104_ net138 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_1
X_2316_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q _1301_ VGND VGND
+ VPWR VPWR _1302_ sky130_fd_sc_hd__nand2_1
X_5035_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 VGND VGND VPWR VPWR net377
+ sky130_fd_sc_hd__buf_4
XFILLER_111_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2247_ net973 net968 net987 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR
+ _1238_ sky130_fd_sc_hd__mux4_1
XFILLER_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2178_ _1172_ _1173_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nand2b_4
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4819_ net1214 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_181_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput102 Tile_X0Y0_W2END[5] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_163_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput113 Tile_X0Y0_W6END[0] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput135 Tile_X0Y1_E2MID[4] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xinput124 Tile_X0Y1_E2END[1] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput157 Tile_X0Y1_FrameData[21] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_2
Xinput146 Tile_X0Y1_FrameData[10] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_2
Xinput168 Tile_X0Y1_FrameData[5] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_2
XFILLER_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 Tile_X0Y1_N2END[2] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput609 net609 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3150_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q VGND VGND VPWR
+ VPWR _0105_ sky130_fd_sc_hd__inv_1
X_2101_ net722 _0620_ _0661_ _0492_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__o22ai_2
X_3081_ net185 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_1
X_2032_ _1022_ _1032_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__nor2_8
XFILLER_94_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3983_ _0543_ _0829_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__or2_1
XFILLER_148_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2934_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q _1808_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q
+ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__o21ai_1
XFILLER_148_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2865_ _1755_ _1756_ _1759_ _0151_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4604_ net1198 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2796_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q _1149_ _1707_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q VGND VGND VPWR VPWR
+ _1708_ sky130_fd_sc_hd__a211oi_1
XFILLER_116_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4535_ net1192 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4466_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3417_ net1042 net1033 net1037 net1054 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q VGND VGND VPWR VPWR
+ _0361_ sky130_fd_sc_hd__mux4_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4397_ net1238 net1152 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3348_ net1216 net73 net217 net229 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0297_ sky130_fd_sc_hd__mux4_1
XFILLER_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3279_ net194 net90 net217 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q VGND VGND VPWR VPWR
+ _0230_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5018_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 VGND VGND VPWR VPWR net360
+ sky130_fd_sc_hd__buf_1
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2650_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q _1602_ VGND VGND
+ VPWR VPWR _1603_ sky130_fd_sc_hd__or2_1
XFILLER_172_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput417 net417 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput406 net406 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[6] sky130_fd_sc_hd__buf_2
X_2581_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q _1537_ VGND VGND
+ VPWR VPWR _1538_ sky130_fd_sc_hd__and2b_1
XFILLER_153_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput428 net428 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[2] sky130_fd_sc_hd__buf_2
X_4320_ net1225 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput439 net439 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4251_ net1253 net1091 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3202_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q VGND VGND VPWR
+ VPWR _0157_ sky130_fd_sc_hd__inv_1
X_4182_ net33 net1110 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3133_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q VGND VGND VPWR
+ VPWR _0088_ sky130_fd_sc_hd__inv_2
XFILLER_121_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3064_ net964 _1611_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__and2b_1
XFILLER_103_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2015_ _1007_ _1010_ _1008_ _1009_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3966_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q _0871_ VGND VGND
+ VPWR VPWR _0872_ sky130_fd_sc_hd__or2_1
XFILLER_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2917_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q _1793_ VGND
+ VGND VPWR VPWR _1794_ sky130_fd_sc_hd__nand2_1
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3897_ net189 net135 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q
+ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__mux2_1
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2848_ net1025 _0407_ _0468_ _0398_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 sky130_fd_sc_hd__mux4_1
X_2779_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q _1694_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q
+ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4518_ net1210 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_104_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4449_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C1 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3820_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net16 net72 net108 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q VGND VGND VPWR VPWR
+ _0733_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_25_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3751_ _0667_ _0666_ _0670_ _0105_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1
+ sky130_fd_sc_hd__a22o_4
XFILLER_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2702_ net1053 _0407_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 _0398_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3682_ _0042_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__a21oi_1
X_2633_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q _1584_ _1586_
+ _0143_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__o211a_1
XFILLER_145_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2564_ net186 net62 net26 net98 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q VGND VGND VPWR VPWR
+ _1522_ sky130_fd_sc_hd__mux4_2
X_4303_ net1240 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_153_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput258 net258 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput247 net247 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput236 net236 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[1] sky130_fd_sc_hd__buf_4
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput269 net269 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_141_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2495_ _1467_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 sky130_fd_sc_hd__mux2_4
XFILLER_59_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4234_ net1233 net1091 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4165_ net1254 net1116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3116_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q VGND VGND VPWR
+ VPWR _0071_ sky130_fd_sc_hd__inv_1
X_4096_ net1225 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3047_ net963 _1464_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__and2b_1
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4998_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 VGND VGND VPWR VPWR net349
+ sky130_fd_sc_hd__buf_6
XFILLER_23_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3949_ _0852_ _0853_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2280_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q _1244_ _1256_
+ _1268_ _0128_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__o221a_1
XFILLER_150_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4921_ Tile_X0Y0_EE4END[9] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_1
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4852_ net1187 net1148 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3803_ net189 net197 net1258 net9 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0718_ sky130_fd_sc_hd__mux4_1
XFILLER_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1995_ _0957_ _0961_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__xor2_2
X_4783_ net1184 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_158_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_109_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3734_ _0060_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q
+ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__a211o_1
XFILLER_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3665_ _0591_ _0100_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__or2_4
X_2616_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q _1569_ VGND VGND
+ VPWR VPWR _1570_ sky130_fd_sc_hd__or2_4
XFILLER_133_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3596_ _0524_ _0523_ _0525_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ _0076_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a221o_1
X_2547_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\]
+ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__and2_1
XFILLER_114_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2478_ _1323_ _1321_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__xor2_2
X_4217_ net1251 net1101 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5197_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net539
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4148_ net35 net1117 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4079_ net1240 net1135 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload1 clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_6
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1203 net154 VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__buf_4
Xfanout1214 net145 VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__clkbuf_4
Xfanout1247 net34 VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__buf_4
Xfanout1225 net52 VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__buf_4
Xfanout1236 Tile_X0Y0_FrameData[26] VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__clkbuf_2
Xfanout1258 net3 VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3450_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q _0391_ _0387_
+ _0360_ _0362_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6
+ sky130_fd_sc_hd__o32a_4
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3381_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0327_ VGND VGND
+ VPWR VPWR _0328_ sky130_fd_sc_hd__nand2_1
X_2401_ net184 net130 net76 net231 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q VGND VGND VPWR VPWR
+ _1382_ sky130_fd_sc_hd__mux4_1
XFILLER_170_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2332_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q _1315_ _1317_
+ _1311_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ sky130_fd_sc_hd__o31ai_4
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5120_ Tile_X0Y1_EE4END[7] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__buf_1
XFILLER_123_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5051_ net107 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_110_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4002_ _0786_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__nand2_1
XFILLER_84_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2263_ net173 net177 net119 net123 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q VGND VGND VPWR VPWR
+ _1254_ sky130_fd_sc_hd__mux4_1
X_2194_ _1188_ _1177_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ sky130_fd_sc_hd__mux2_4
XFILLER_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4904_ Tile_X0Y0_E6END[2] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_1
XFILLER_33_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4835_ net1206 net1156 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4766_ net1200 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3717_ net1036 net1008 net1032 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0639_ sky130_fd_sc_hd__mux4_1
X_1978_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q _0969_ _0979_
+ _0973_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B0 sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_31_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4697_ net1195 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3648_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\] net1062 VGND VGND VPWR VPWR _0575_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3579_ _0077_ _0510_ _0509_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__o211a_1
XFILLER_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5249_ Tile_X0Y1_WW4END[4] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1011 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 VGND VGND VPWR VPWR
+ net1011 sky130_fd_sc_hd__clkbuf_4
Xfanout1022 net676 VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__buf_8
XFILLER_126_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1000 net1001 VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__buf_8
Xfanout1055 net1056 VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__buf_2
Xfanout1033 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 VGND VGND VPWR VPWR
+ net1033 sky130_fd_sc_hd__buf_2
Xfanout1044 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 VGND VGND VPWR VPWR
+ net1044 sky130_fd_sc_hd__buf_8
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1066 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q VGND VGND
+ VPWR VPWR net1066 sky130_fd_sc_hd__clkbuf_4
Xfanout1077 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1088 net1089 VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1099 net1102 VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__buf_2
XFILLER_19_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2950_ _0155_ _1814_ _1819_ _1823_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0
+ sky130_fd_sc_hd__a31o_1
X_2881_ net202 net1217 net124 net1215 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _1767_ sky130_fd_sc_hd__mux4_1
X_4620_ net1181 net1112 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4551_ net1211 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3502_ _0434_ _0436_ _0439_ _0071_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2
+ sky130_fd_sc_hd__a22o_1
X_4482_ net1205 net1174 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3433_ _0374_ _0375_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q
+ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux2_4
X_3364_ net1019 net1014 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__mux2_1
X_5103_ net137 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_2
X_3295_ _0084_ _0245_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__or2_1
X_2315_ _1301_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6
+ sky130_fd_sc_hd__inv_4
X_5034_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 VGND VGND VPWR VPWR net376
+ sky130_fd_sc_hd__buf_1
X_2246_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q _1236_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__o21ba_1
X_2177_ _1170_ _1171_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__nand2b_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4818_ net1202 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_31_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4749_ net1182 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput114 Tile_X0Y0_W6END[1] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_4
Xinput103 Tile_X0Y0_W2END[6] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput136 Tile_X0Y1_E2MID[5] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
Xinput125 Tile_X0Y1_E2END[2] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_2
XFILLER_48_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput158 Tile_X0Y1_FrameData[22] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_2
Xinput147 Tile_X0Y1_FrameData[11] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
Xinput169 Tile_X0Y1_FrameData[6] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_2
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2100_ _0854_ _0857_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__nor2_1
XFILLER_94_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3080_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q VGND VGND VPWR
+ VPWR _0035_ sky130_fd_sc_hd__inv_2
XFILLER_39_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2031_ _1023_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_109_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3982_ _0883_ _0884_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__xnor2_1
X_2933_ _1807_ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__inv_1
XFILLER_148_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2864_ _1757_ _1758_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q
+ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__mux2_1
XFILLER_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2795_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q net1054 VGND
+ VGND VPWR VPWR _1707_ sky130_fd_sc_hd__nor2_1
X_4603_ net1197 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4534_ net1191 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4465_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3416_ _0092_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__and2_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4396_ net1237 net1152 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3347_ net181 net1218 net193 net127 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q VGND VGND VPWR VPWR
+ _0296_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_168_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5017_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 VGND VGND VPWR VPWR net359
+ sky130_fd_sc_hd__buf_1
XFILLER_45_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3278_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR _0229_
+ sky130_fd_sc_hd__inv_2
X_2229_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q _1217_ _1221_
+ _1212_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 sky130_fd_sc_hd__a31o_1
XFILLER_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput407 net407 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[7] sky130_fd_sc_hd__buf_2
X_2580_ net690 net14 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q
+ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__mux2_1
XFILLER_153_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput418 net418 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput429 net429 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4250_ net1252 net1091 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4181_ net1247 net1108 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3201_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q VGND VGND VPWR
+ VPWR _0156_ sky130_fd_sc_hd__inv_1
X_3132_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR
+ VPWR _0087_ sky130_fd_sc_hd__inv_2
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3063_ net964 _1614_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__and2b_1
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2014_ _1014_ _1013_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__and2b_1
X_3965_ net60 net68 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q VGND
+ VGND VPWR VPWR _0871_ sky130_fd_sc_hd__mux2_1
XFILLER_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2916_ _0818_ _1437_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q
+ VGND VGND VPWR VPWR _1793_ sky130_fd_sc_hd__mux2_1
X_3896_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q _0803_ VGND VGND
+ VPWR VPWR _0804_ sky130_fd_sc_hd__and2_4
X_2847_ _1747_ _1752_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1
+ sky130_fd_sc_hd__or2_1
XFILLER_148_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2778_ _1693_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__inv_1
XFILLER_151_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4517_ net1209 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4448_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C0 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4379_ net28 net1162 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3750_ _0668_ _0669_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q
+ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__mux2_1
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2701_ net186 net113 net197 net695 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 sky130_fd_sc_hd__mux4_1
X_3681_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q _0243_ VGND VGND
+ VPWR VPWR _0606_ sky130_fd_sc_hd__or2_1
X_2632_ _0142_ _1585_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__or2_1
XFILLER_145_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2563_ _1502_ _1517_ _1518_ _1516_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__o31a_1
X_4302_ net1239 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_160_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput259 net259 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput248 net248 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput237 net237 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_126_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4233_ net45 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_113_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2494_ _1389_ _1449_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__xnor2_2
XFILLER_4_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4164_ net1243 net1116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3115_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q VGND VGND VPWR
+ VPWR _0070_ sky130_fd_sc_hd__inv_2
X_4095_ net1224 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3046_ net963 _1615_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_124_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4997_ net666 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__buf_6
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3948_ _0852_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__nor2_2
XFILLER_176_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3879_ _0601_ _0709_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__or2_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4920_ Tile_X0Y0_EE4END[8] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_63_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4851_ net1214 net1156 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3802_ _0716_ _0066_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__o21a_1
X_1994_ _0990_ _0991_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__xor2_1
XFILLER_60_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4782_ net168 net1072 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3733_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q net710 VGND VGND
+ VPWR VPWR _0654_ sky130_fd_sc_hd__nor2_2
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3664_ net982 net996 net1018 net1001 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0591_ sky130_fd_sc_hd__mux4_2
X_2615_ net57 net59 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q VGND
+ VGND VPWR VPWR _1569_ sky130_fd_sc_hd__mux2_2
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3595_ _0524_ _0523_ _0525_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__a22o_4
X_2546_ _1115_ _1480_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q
+ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__a21bo_2
X_2477_ _1452_ _1344_ _1343_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__a21o_1
X_5196_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net538
+ sky130_fd_sc_hd__buf_6
X_4216_ net1250 net1101 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4147_ net1245 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4078_ net1239 net1135 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_141_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3029_ net707 net743 net716 net980 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q VGND VGND VPWR VPWR
+ _1892_ sky130_fd_sc_hd__mux4_1
XFILLER_36_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_174_Right_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload2 clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinv_2
XFILLER_166_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1204 net153 VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__buf_4
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput590 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 VGND VGND VPWR VPWR
+ Tile_X0Y1_W6BEG[11] sky130_fd_sc_hd__buf_6
Xfanout1237 net44 VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__buf_4
Xfanout1226 net51 VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__buf_4
XFILLER_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1215 net140 VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__buf_2
Xfanout1248 net33 VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__buf_4
XFILLER_93_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2400_ net196 net84 net141 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q VGND VGND VPWR VPWR
+ _1381_ sky130_fd_sc_hd__mux4_1
XFILLER_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3380_ net200 net8 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q VGND
+ VGND VPWR VPWR _0327_ sky130_fd_sc_hd__mux2_1
XFILLER_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2331_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q _1316_ VGND VGND
+ VPWR VPWR _1317_ sky130_fd_sc_hd__nor2_1
X_5050_ net106 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_2
X_2262_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q _1250_ _1252_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR VPWR
+ _1253_ sky130_fd_sc_hd__o211a_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4001_ _0709_ _0878_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__nor2_1
XFILLER_84_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2193_ _1187_ _0526_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__mux2_1
XFILLER_84_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4903_ net20 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4834_ net152 net1156 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_178_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4765_ net1199 net1070 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3716_ _0088_ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__and2_1
XFILLER_146_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1977_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q _0978_ VGND VGND
+ VPWR VPWR _0979_ sky130_fd_sc_hd__nor2_1
X_4696_ net1193 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3647_ _0569_ _0568_ _0573_ net1061 VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__a211o_4
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3578_ net1034 net736 net1029 net676 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _0510_ sky130_fd_sc_hd__mux4_2
X_2529_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q _1491_ VGND VGND
+ VPWR VPWR _1492_ sky130_fd_sc_hd__or2_1
XFILLER_161_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5179_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR net530
+ sky130_fd_sc_hd__buf_2
XFILLER_68_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1012 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 VGND VGND VPWR VPWR
+ net1012 sky130_fd_sc_hd__buf_2
XFILLER_105_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1001 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 VGND VGND VPWR VPWR net1001
+ sky130_fd_sc_hd__buf_12
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1023 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 VGND VGND VPWR VPWR
+ net1023 sky130_fd_sc_hd__buf_8
Xfanout1056 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 VGND VGND VPWR VPWR
+ net1056 sky130_fd_sc_hd__buf_8
Xfanout1045 net1048 VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__buf_8
Xfanout1034 net1035 VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__buf_8
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1089 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__clkbuf_2
Xfanout1067 net212 VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__clkbuf_4
Xfanout1078 net1081 VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__buf_2
XFILLER_74_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ net70 net82 net214 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _1766_ sky130_fd_sc_hd__mux4_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4550_ net1210 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3501_ _0437_ _0438_ _0070_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__mux2_1
XFILLER_128_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4481_ net1204 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3432_ net980 net995 net1016 net1013 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0375_ sky130_fd_sc_hd__mux4_1
XFILLER_143_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3363_ _0055_ net997 _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__o21a_1
XFILLER_97_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5102_ net136 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_1
X_3294_ net2 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q VGND
+ VGND VPWR VPWR _0245_ sky130_fd_sc_hd__mux2_1
X_2314_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q _1300_ _1298_
+ _1292_ _1293_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__o32a_4
X_5033_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 VGND VGND VPWR VPWR net375
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_111_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2245_ net173 net177 net119 net123 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR
+ _1236_ sky130_fd_sc_hd__mux4_1
XFILLER_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2176_ _1171_ _1170_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__and2b_1
XFILLER_65_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4817_ net1190 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_178_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4748_ net1181 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4679_ net148 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput115 Tile_X0Y0_WW4END[0] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
Xinput104 Tile_X0Y0_W2END[7] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_2
Xinput126 Tile_X0Y1_E2END[3] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput159 Tile_X0Y1_FrameData[23] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_2
Xinput148 Tile_X0Y1_FrameData[12] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_2
Xinput137 Tile_X0Y1_E2MID[6] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_2
XFILLER_56_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_136_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2030_ _1030_ _1029_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_145_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3981_ _0883_ _0884_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__or2_1
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2932_ net1015 _1410_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q
+ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__mux2_4
XFILLER_148_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2863_ net1215 net214 net70 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q VGND VGND VPWR VPWR
+ _1758_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_154_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2794_ _1703_ _1706_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 sky130_fd_sc_hd__mux2_1
X_4602_ net1196 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4533_ net1189 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_156_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4464_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3415_ net1011 net1046 net1026 net1052 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR VPWR
+ _0359_ sky130_fd_sc_hd__mux4_1
XFILLER_171_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4395_ net1235 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3346_ _0293_ _0294_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q
+ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_168_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_163_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5016_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net358
+ sky130_fd_sc_hd__buf_1
X_3277_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q _0224_ _0228_
+ _0222_ _0220_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ sky130_fd_sc_hd__o32a_4
X_2228_ _1218_ _1219_ _1220_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q VGND VGND VPWR VPWR
+ _1221_ sky130_fd_sc_hd__a221o_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ _1154_ _1155_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__xor2_2
XFILLER_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_172_Left_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_181_Left_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput408 net408 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_153_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput419 net419 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_153_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4180_ net1246 net1108 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3200_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q VGND VGND VPWR
+ VPWR _0155_ sky130_fd_sc_hd__inv_1
X_3131_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR
+ VPWR _0086_ sky130_fd_sc_hd__inv_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3062_ net964 _1548_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__and2b_1
X_2013_ _0965_ _0986_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__xnor2_2
XFILLER_90_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3964_ _0867_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q _0869_
+ _0096_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__o211a_1
XFILLER_50_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2915_ _1791_ _1792_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 sky130_fd_sc_hd__mux2_1
X_3895_ _0802_ _0801_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q
+ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__mux2_4
X_2846_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q _1748_ _1751_
+ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__o21a_1
XFILLER_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2777_ net1028 net1051 net1043 net1038 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q VGND VGND VPWR VPWR
+ _1693_ sky130_fd_sc_hd__mux4_1
XFILLER_163_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4516_ net1208 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4447_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_4378_ net29 net1162 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3329_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q _0260_ _0276_
+ _0275_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q VGND VGND VPWR
+ VPWR _0279_ sky130_fd_sc_hd__o221a_4
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2700_ net185 net200 net114 net1006 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 sky130_fd_sc_hd__mux4_1
X_3680_ _0062_ _0604_ _0603_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q
+ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__o211a_1
X_2631_ net1 net5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q VGND
+ VGND VPWR VPWR _1585_ sky130_fd_sc_hd__mux2_1
XFILLER_160_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2562_ _1520_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 sky130_fd_sc_hd__mux2_4
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4301_ net43 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput249 net249 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput238 net238 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_99_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4232_ net1231 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2493_ _1466_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 sky130_fd_sc_hd__mux2_2
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4163_ net1230 net1116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3114_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q VGND VGND VPWR
+ VPWR _0069_ sky130_fd_sc_hd__inv_1
X_4094_ net1223 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3045_ net963 _1466_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__and2b_1
XFILLER_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4996_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 VGND VGND VPWR VPWR net347
+ sky130_fd_sc_hd__buf_6
XFILLER_23_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3947_ _0493_ _0761_ _0760_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__o21a_1
XFILLER_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3878_ _0620_ _0785_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__nor2_1
XFILLER_31_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2829_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q _1734_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q
+ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__o21ai_1
XFILLER_136_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4850_ net1202 net1157 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_160_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3801_ net1035 net736 net695 net1023 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0716_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_71_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1993_ _0955_ _0992_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__xnor2_2
X_4781_ net169 net1072 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_158_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3732_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q _0649_ _0650_
+ _0651_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q VGND VGND VPWR
+ VPWR _0653_ sky130_fd_sc_hd__a221o_1
XFILLER_173_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3663_ net972 net986 net990 net976 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0590_ sky130_fd_sc_hd__mux4_2
XFILLER_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2614_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q _1565_ _1567_
+ _0146_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__o211a_1
XFILLER_133_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3594_ net76 net112 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q
+ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__mux2_1
X_2545_ _1505_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 sky130_fd_sc_hd__mux2_4
XFILLER_126_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2476_ _1451_ _1359_ _1358_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__a21o_1
X_5195_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net537
+ sky130_fd_sc_hd__buf_4
X_4215_ net1249 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4146_ net1244 net1117 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4077_ net43 net1135 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3028_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q _1890_ VGND VGND
+ VPWR VPWR _1891_ sky130_fd_sc_hd__nor2_1
XFILLER_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4979_ Tile_X0Y1_FrameStrobe[15] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_1
XFILLER_149_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1205 net152 VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__clkbuf_4
Xoutput580 net580 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_182_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1238 net43 VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__buf_4
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1227 net50 VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__buf_4
Xoutput591 net591 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[1] sky130_fd_sc_hd__buf_2
Xfanout1216 net139 VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1249 net32 VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_77_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2330_ net176 net184 net1217 net130 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR VPWR
+ _1316_ sky130_fd_sc_hd__mux4_1
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2261_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q _1251_ VGND VGND
+ VPWR VPWR _1252_ sky130_fd_sc_hd__nand2_1
XFILLER_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4000_ _0897_ _0898_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__xnor2_1
X_2192_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 net19 net111 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q
+ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__mux4_1
XFILLER_92_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4902_ net19 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__buf_1
XFILLER_52_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4833_ net153 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1976_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q _0977_ _0975_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q VGND VGND VPWR VPWR
+ _0978_ sky130_fd_sc_hd__o211a_1
X_4764_ net159 net1070 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3715_ net1011 net1046 net1027 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0637_ sky130_fd_sc_hd__mux4_1
XFILLER_146_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4695_ net1192 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3646_ _0568_ _0569_ _0573_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B3 sky130_fd_sc_hd__a21o_1
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3577_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q _0508_ VGND VGND
+ VPWR VPWR _0509_ sky130_fd_sc_hd__or2_4
X_2528_ net58 net60 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q VGND
+ VGND VPWR VPWR _1491_ sky130_fd_sc_hd__mux2_1
X_5247_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 VGND VGND VPWR VPWR net589
+ sky130_fd_sc_hd__buf_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2459_ net196 net126 net216 net658 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q VGND VGND VPWR VPWR
+ _1436_ sky130_fd_sc_hd__mux4_1
XFILLER_152_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5178_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 VGND VGND VPWR VPWR net529
+ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_180_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4129_ net1226 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1002 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 VGND VGND VPWR VPWR net1002
+ sky130_fd_sc_hd__clkbuf_2
Xfanout1013 net1015 VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__buf_8
Xfanout1046 net1047 VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__clkbuf_4
Xfanout1024 net1025 VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__buf_8
Xfanout1035 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 VGND VGND VPWR VPWR
+ net1035 sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_58_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1057 _0099_ VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__clkbuf_4
Xfanout1068 net211 VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__buf_4
XFILLER_59_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1079 net1081 VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__buf_2
XFILLER_74_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3500_ net188 net200 net2 net8 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0438_ sky130_fd_sc_hd__mux4_1
XFILLER_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4480_ net1203 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3431_ net971 net728 net991 net975 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0374_ sky130_fd_sc_hd__mux4_1
X_3362_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q net978 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__o21ba_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2313_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q _1299_ VGND VGND
+ VPWR VPWR _1300_ sky130_fd_sc_hd__nor2_1
X_5101_ net135 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_1
X_3293_ _0243_ net190 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_1
X_5032_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 VGND VGND VPWR VPWR net374
+ sky130_fd_sc_hd__buf_1
XFILLER_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2244_ _0133_ _1232_ _1234_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__a21o_1
XFILLER_122_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2175_ _0903_ _1096_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__xnor2_2
XFILLER_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4816_ net166 net1164 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1959_ _0960_ _0958_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__xnor2_2
X_4747_ net1180 net1079 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4678_ net149 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3629_ _0548_ _0550_ _0106_ _0556_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__a211o_1
XFILLER_134_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput116 Tile_X0Y0_WW4END[1] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput105 Tile_X0Y0_W2MID[0] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput127 Tile_X0Y1_E2END[4] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput149 Tile_X0Y1_FrameData[13] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_2
Xinput138 Tile_X0Y1_E2MID[7] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
XFILLER_56_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3980_ _0788_ _0789_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2931_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q _1349_ _1805_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _1806_ sky130_fd_sc_hd__o211a_1
XFILLER_148_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4601_ net1195 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2862_ net176 net178 net194 net142 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _1757_ sky130_fd_sc_hd__mux4_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2793_ _1704_ _1705_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__mux2_1
XFILLER_156_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4532_ net1187 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4463_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3414_ _0083_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q
+ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__a21oi_1
XFILLER_116_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4394_ net1233 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3345_ net980 net995 net1016 net1013 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0294_ sky130_fd_sc_hd__mux4_1
X_3276_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q _0225_ _0226_
+ _0227_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q VGND VGND VPWR
+ VPWR _0228_ sky130_fd_sc_hd__o221a_1
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2227_ net987 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__mux2_1
X_5015_ Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_6
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ _1154_ _1155_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__and2_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2089_ _1055_ _1089_ _1054_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput409 net409 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[10] sky130_fd_sc_hd__buf_2
XFILLER_99_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3130_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q VGND VGND VPWR
+ VPWR _0085_ sky130_fd_sc_hd__inv_2
XFILLER_79_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3061_ net964 _1520_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ _0996_ _1005_ _1012_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__a21o_1
XFILLER_90_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3963_ _0095_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__or2_1
XFILLER_35_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3894_ net181 net127 net91 net217 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q VGND VGND VPWR VPWR
+ _0802_ sky130_fd_sc_hd__mux4_2
X_2914_ net998 _0767_ _0940_ _1382_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q VGND VGND VPWR VPWR
+ _1792_ sky130_fd_sc_hd__mux4_1
X_2845_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q _1750_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q
+ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2776_ net1258 net1012 net1220 net1047 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q VGND VGND VPWR VPWR
+ _1692_ sky130_fd_sc_hd__mux4_1
XFILLER_163_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4515_ net1206 net1140 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4446_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\] sky130_fd_sc_hd__dfxtp_1
X_4377_ net30 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_104_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3328_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkinv_2
X_3259_ _0211_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q _0210_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q VGND VGND VPWR VPWR
+ _0212_ sky130_fd_sc_hd__o211a_1
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2630_ _0199_ net185 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__mux2_1
XFILLER_159_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2561_ _1517_ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__xnor2_1
Xclone90 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 VGND VGND VPWR VPWR net707
+ sky130_fd_sc_hd__buf_6
X_4300_ net1237 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_160_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput239 net239 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_126_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2492_ _1443_ _1465_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__nor2_1
XFILLER_153_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4231_ net1229 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4162_ net1227 net1116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3113_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q VGND VGND VPWR
+ VPWR _0068_ sky130_fd_sc_hd__inv_2
X_4093_ net1222 net1133 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3044_ _1898_ _1905_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4995_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 VGND VGND VPWR VPWR net346
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_90_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3946_ _0849_ _0850_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__xor2_1
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3877_ _0659_ _0660_ _0784_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__and3_1
X_2828_ net1044 net1036 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__mux2_1
X_2759_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q _1675_ _1674_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q VGND VGND VPWR VPWR
+ _1676_ sky130_fd_sc_hd__o211a_1
XFILLER_117_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4429_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0017_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3800_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q _0714_ VGND VGND
+ VPWR VPWR _0715_ sky130_fd_sc_hd__or2_4
X_4780_ net170 net1070 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_158_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3731_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q _0649_ _0650_
+ _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__a22o_2
X_1992_ _0992_ _0955_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_71_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3662_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q _0582_ _0584_
+ _0587_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__o32a_1
X_2613_ _0145_ _1566_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__or2_4
X_3593_ _0044_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2544_ _1504_ _1479_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__xnor2_2
XFILLER_141_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2475_ _1370_ _1450_ _1369_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__a21o_1
X_5263_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net605
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5194_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net551
+ sky130_fd_sc_hd__buf_4
X_4214_ net1248 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4145_ net1242 net1117 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4076_ net44 net1135 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_55_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3027_ net1218 net1068 net971 net691 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR
+ _1890_ sky130_fd_sc_hd__mux4_1
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4978_ Tile_X0Y1_FrameStrobe[14] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3929_ _0793_ _0834_ _0792_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__o21ba_4
XFILLER_164_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput570 net570 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput581 net581 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[1] sky130_fd_sc_hd__buf_2
Xfanout1228 net49 VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__buf_4
XFILLER_105_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1206 net1207 VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__buf_4
Xfanout1217 net122 VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__clkbuf_4
Xoutput592 net592 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[2] sky130_fd_sc_hd__buf_2
Xfanout1239 net42 VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__buf_4
XFILLER_115_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2260_ net209 net211 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__mux2_1
XFILLER_69_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2191_ _1186_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_162_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4901_ net18 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4832_ net1203 net1156 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1975_ _0976_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__inv_1
X_4763_ net160 net1070 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3714_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q _0635_ VGND VGND
+ VPWR VPWR _0636_ sky130_fd_sc_hd__and2_1
X_4694_ net1191 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_132_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3645_ _0110_ _0570_ _0572_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q
+ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__o211a_1
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3576_ net1045 net750 net713 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _0508_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_93_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2527_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q _1487_ _1489_
+ _0094_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__o211a_1
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5246_ Tile_X0Y1_W6END[11] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__clkbuf_2
X_2458_ _1434_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5177_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 VGND VGND VPWR VPWR net528
+ sky130_fd_sc_hd__buf_4
X_2389_ _1368_ _1367_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__xnor2_4
X_4128_ net1225 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4059_ net1253 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1003 _1361_ VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__clkbuf_4
Xfanout1047 net1048 VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__buf_2
Xfanout1036 net1038 VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__clkbuf_4
Xfanout1025 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 VGND VGND VPWR VPWR
+ net1025 sky130_fd_sc_hd__buf_8
XFILLER_120_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1014 net1015 VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1058 _0099_ VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__buf_4
Xfanout1069 net1070 VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__buf_2
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3430_ net204 net231 net84 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q VGND VGND VPWR VPWR
+ _0373_ sky130_fd_sc_hd__mux4_2
XFILLER_143_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3361_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q _0308_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q
+ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__o21ba_1
XFILLER_97_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2312_ net176 net184 net1217 net130 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR
+ _1299_ sky130_fd_sc_hd__mux4_1
X_5100_ net134 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_2
XFILLER_151_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3292_ net663 _0218_ _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a21o_4
X_5031_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__buf_4
X_2243_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q _1233_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q
+ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__a21bo_1
X_2174_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\] _1169_ net1058 VGND VGND VPWR VPWR
+ _1170_ sky130_fd_sc_hd__mux2_1
XFILLER_178_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4815_ net1184 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_178_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1958_ _0912_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__xor2_2
X_4746_ net1179 net1079 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4677_ net1209 net1096 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3628_ _0548_ _0550_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__a21oi_4
XFILLER_163_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3559_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ net1060 _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__o21ai_4
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput117 Tile_X0Y0_WW4END[2] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
Xinput106 Tile_X0Y0_W2MID[1] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput128 Tile_X0Y1_E2END[5] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_2
Xinput139 Tile_X0Y1_E6END[0] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlymetal6s2s_1
X_5229_ net221 VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__buf_1
XFILLER_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2930_ _0860_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q VGND
+ VGND VPWR VPWR _1805_ sky130_fd_sc_hd__nand2b_1
XFILLER_148_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4600_ net1193 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2861_ _0150_ _1753_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_41_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2792_ net965 _0615_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__mux2_1
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4531_ net1214 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_156_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4462_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3413_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6
+ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__or2_1
XFILLER_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4393_ net1232 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3344_ net971 net728 net985 net975 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0293_ sky130_fd_sc_hd__mux4_1
XFILLER_97_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3275_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q net233 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a21bo_1
X_2226_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q net973 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__o21ba_1
X_5014_ Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__buf_4
XFILLER_26_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ _1097_ _1099_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__xnor2_2
XFILLER_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2088_ _1070_ _1088_ _1069_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_179_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4729_ net162 net1081 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_181_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_86_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_95_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3060_ net964 _1505_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__and2b_1
XFILLER_121_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2011_ _1011_ _1006_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__nor2_1
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3962_ net1257 net12 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__mux2_1
XFILLER_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3893_ net202 net142 net82 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q VGND VGND VPWR VPWR
+ _0801_ sky130_fd_sc_hd__mux4_2
X_2913_ net175 net1218 _0302_ net989 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q VGND VGND VPWR VPWR
+ _1791_ sky130_fd_sc_hd__mux4_1
X_2844_ _1749_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__inv_1
XFILLER_148_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2775_ _1687_ _1689_ _1690_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q VGND VGND VPWR VPWR
+ _1691_ sky130_fd_sc_hd__o221a_1
X_4514_ net1205 net1140 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4445_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4376_ net1250 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3327_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q _0260_ _0275_
+ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__o22a_1
XFILLER_112_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3258_ net1009 net1045 net1024 net1049 net617 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux4_2
X_3189_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR
+ VPWR _0144_ sky130_fd_sc_hd__inv_1
X_2209_ net175 net121 net183 net129 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q VGND VGND VPWR VPWR
+ _1203_ sky130_fd_sc_hd__mux4_1
XFILLER_81_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2560_ _1502_ _1518_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__nor2_2
XFILLER_126_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone91 net1010 VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__buf_8
XFILLER_153_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2491_ _1081_ _1442_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__nor2_1
XFILLER_126_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4230_ net1228 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_99_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4161_ net1226 net1118 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3112_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q VGND VGND VPWR
+ VPWR _0067_ sky130_fd_sc_hd__inv_1
X_4092_ net1221 net1133 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3043_ _1899_ _1900_ _1904_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q
+ VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4994_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 VGND VGND VPWR VPWR net345
+ sky130_fd_sc_hd__buf_1
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3945_ _0849_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__and2b_1
XFILLER_176_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3876_ _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__clkinv_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2827_ _1733_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__inv_1
XFILLER_136_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2758_ net740 net1032 net1022 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q VGND VGND VPWR VPWR
+ _1675_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_96_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2689_ _0047_ _1633_ _1632_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__o211a_1
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4428_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0016_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4359_ net48 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_169_Left_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_178_Left_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout990 net991 VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__buf_2
XFILLER_64_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _0080_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q
+ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__a21oi_1
X_1991_ _0990_ _0991_ _0989_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_71_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3661_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q _0585_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q
+ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__a21bo_1
XFILLER_173_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2612_ net1 net5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q VGND
+ VGND VPWR VPWR _1566_ sky130_fd_sc_hd__mux2_2
X_3592_ _0417_ _0415_ _0424_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q
+ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_171_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2543_ _1502_ _1503_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__and2b_1
XFILLER_126_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2474_ _1388_ _1449_ _1387_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__o21bai_4
XTAP_TAPCELL_ROW_130_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5193_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net550
+ sky130_fd_sc_hd__buf_4
X_4213_ net1247 net1101 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4144_ net1241 net1117 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4075_ net1235 net1135 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3026_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q _1888_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q
+ VGND VGND VPWR VPWR _1889_ sky130_fd_sc_hd__o21ai_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4977_ Tile_X0Y1_FrameStrobe[13] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_1
XFILLER_149_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3928_ _0830_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__xnor2_4
XFILLER_166_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3859_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q _0768_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__o21a_1
XFILLER_166_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput571 net571 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput560 net560 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[2] sky130_fd_sc_hd__buf_2
Xfanout1229 net48 VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__buf_4
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1207 Tile_X0Y1_FrameData[16] VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__clkbuf_2
Xfanout1218 net121 VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__buf_4
Xoutput582 net582 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput593 net593 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_115_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2190_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q _1179_ _1181_
+ _1185_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__a31o_1
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4900_ net17 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_1
XFILLER_18_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4831_ net1201 net1156 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_178_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1974_ net192 net138 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q
+ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__mux2_1
X_4762_ net1196 net1070 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3713_ _0634_ _0633_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__mux2_1
X_4693_ net1188 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3644_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q _0571_ VGND VGND
+ VPWR VPWR _0572_ sky130_fd_sc_hd__or2_1
XFILLER_161_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3575_ _0079_ _0506_ _0505_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__o211a_1
X_2526_ _0093_ _1488_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__or2_1
XFILLER_114_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2457_ _1073_ _1081_ _1433_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__a21o_1
X_5245_ Tile_X0Y1_W6END[10] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__clkbuf_2
XFILLER_152_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5176_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 VGND VGND VPWR VPWR net527
+ sky130_fd_sc_hd__buf_6
X_2388_ _1368_ _1367_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__and2b_1
X_4127_ net1224 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4058_ net1252 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_43_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3009_ net974 net969 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__mux2_1
XFILLER_101_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1004 net1005 VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__buf_8
XFILLER_105_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1037 net1038 VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__clkbuf_2
Xfanout1026 net1028 VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__buf_2
Xoutput390 net390 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[2] sky130_fd_sc_hd__buf_2
Xfanout1015 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 VGND VGND VPWR VPWR net1015
+ sky130_fd_sc_hd__buf_12
Xfanout1048 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 VGND VGND VPWR VPWR
+ net1048 sky130_fd_sc_hd__buf_12
XFILLER_86_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1059 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q VGND VGND
+ VPWR VPWR net1059 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_106_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3360_ net175 net1218 net183 net129 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR VPWR
+ _0308_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_115_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2311_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q _1297_ _1295_
+ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__and3_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3291_ _0040_ _0230_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q
+ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__o211a_4
X_5030_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_4
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2242_ net69 net209 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__mux2_1
X_2173_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[11\] net1064 VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__mux2_1
XFILLER_111_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4814_ net1183 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4745_ net146 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1957_ _0676_ _0450_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__nor2_4
XFILLER_174_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4676_ net1208 net1096 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3627_ _0554_ _0552_ _0555_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q VGND VGND VPWR VPWR
+ _0556_ sky130_fd_sc_hd__o221a_4
XFILLER_134_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3558_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\] net1060 VGND VGND VPWR VPWR _0491_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_163_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2509_ _1474_ _1457_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__nor2_2
XFILLER_142_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput118 Tile_X0Y0_WW4END[3] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
Xinput107 Tile_X0Y0_W2MID[2] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
X_3489_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q _0427_ VGND VGND
+ VPWR VPWR _0428_ sky130_fd_sc_hd__nand2_1
X_5228_ net220 VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__buf_1
Xinput129 Tile_X0Y1_E2END[6] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_2
X_5159_ net162 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2860_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q _1754_ VGND VGND
+ VPWR VPWR _1755_ sky130_fd_sc_hd__or2_1
XFILLER_175_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2791_ net676 net623 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4530_ net1202 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4461_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_123_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3412_ _0354_ _0356_ _0258_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6
+ sky130_fd_sc_hd__a21o_2
XFILLER_171_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4392_ net1231 net1151 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3343_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q VGND VGND VPWR VPWR
+ _0292_ sky130_fd_sc_hd__o21ai_4
X_3274_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q net217 VGND VGND
+ VPWR VPWR _0226_ sky130_fd_sc_hd__and2b_1
XFILLER_97_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2225_ net968 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q VGND VGND
+ VPWR VPWR _1218_ sky130_fd_sc_hd__nand2b_1
X_5013_ Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_127_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\] _1153_ net1058 VGND VGND VPWR VPWR
+ _1154_ sky130_fd_sc_hd__mux2_4
XFILLER_93_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_132_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2087_ _1085_ _1086_ _1079_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_179_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2989_ _0818_ _1408_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q
+ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__mux2_1
XFILLER_147_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4728_ net1193 net1081 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_141_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4659_ net1214 net1105 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_150_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2010_ _1010_ _1007_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__xnor2_4
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3961_ net673 net192 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__mux2_1
XFILLER_90_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2912_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q _1785_ _1790_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A sky130_fd_sc_hd__o21a_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3892_ _0797_ _0795_ _0800_ _0119_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ sky130_fd_sc_hd__a22o_4
XFILLER_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2843_ net1026 net1050 net1042 net1036 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q VGND VGND VPWR VPWR
+ _1749_ sky130_fd_sc_hd__mux4_1
X_2774_ net1007 net1032 net1021 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q VGND VGND VPWR VPWR
+ _1690_ sky130_fd_sc_hd__mux4_1
XFILLER_163_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4513_ net1204 net1140 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_174_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4444_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4375_ net1249 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3326_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q net97 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q
+ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__o21ai_1
XFILLER_112_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3257_ _0207_ _0208_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ _0209_ _0037_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3188_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q VGND VGND VPWR
+ VPWR _0143_ sky130_fd_sc_hd__inv_2
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2208_ _0410_ _0302_ net75 net1068 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ _1202_ sky130_fd_sc_hd__mux4_2
X_2139_ net207 net6 net62 net98 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q VGND VGND VPWR VPWR
+ _1139_ sky130_fd_sc_hd__mux4_2
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone92 net1015 VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__clkbuf_1
XFILLER_153_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2490_ _1464_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 sky130_fd_sc_hd__mux2_4
XFILLER_57_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4160_ net1225 net1118 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3111_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q VGND VGND VPWR
+ VPWR _0066_ sky130_fd_sc_hd__inv_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4091_ net28 net1133 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_66_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3042_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 _1895_ _1902_ _1903_ VGND
+ VGND VPWR VPWR _1904_ sky130_fd_sc_hd__a211o_1
XFILLER_48_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4993_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 VGND VGND VPWR VPWR net344
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_90_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3944_ _0743_ _0755_ _0757_ _0754_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3875_ Tile_X0Y1_DSP_bot.A1 Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\] net1060 VGND
+ VGND VPWR VPWR _0784_ sky130_fd_sc_hd__mux2_4
X_2826_ net1026 net1050 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__mux2_1
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2757_ _1673_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q VGND
+ VGND VPWR VPWR _1674_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_135_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2688_ net1037 net1007 net1031 net1021 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _1633_ sky130_fd_sc_hd__mux4_1
X_4427_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0015_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4358_ net49 net1160 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3309_ net205 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q VGND VGND
+ VPWR VPWR _0259_ sky130_fd_sc_hd__or2_1
X_4289_ net1226 net1083 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout980 net981 VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__buf_12
Xfanout991 net994 VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__buf_8
XFILLER_37_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1990_ _0987_ _0988_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__xor2_1
XFILLER_158_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3660_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q _0586_ VGND VGND
+ VPWR VPWR _0587_ sky130_fd_sc_hd__and2b_1
X_2611_ net744 net185 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__mux2_1
X_3591_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q
+ _0521_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q VGND VGND VPWR
+ VPWR _0522_ sky130_fd_sc_hd__o211a_4
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2542_ _1115_ _1480_ _1501_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__a21o_1
XFILLER_126_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5261_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR net603
+ sky130_fd_sc_hd__buf_1
X_4212_ net1246 net1101 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2473_ _1407_ _1448_ _1406_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__o21a_4
X_5192_ Tile_X0Y0_S4END[15] VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_130_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4143_ net41 net1117 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_122_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4074_ net1233 net1135 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3025_ net995 net1016 net714 net709 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR
+ _1888_ sky130_fd_sc_hd__mux4_1
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4976_ net1151 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3927_ _0577_ _0831_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3858_ _0113_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__or2_1
XFILLER_164_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2809_ net618 net1219 net60 net1050 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q VGND VGND VPWR VPWR
+ _1719_ sky130_fd_sc_hd__mux4_1
X_3789_ _0703_ _0704_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q
+ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__mux2_4
XFILLER_105_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput572 net572 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput550 net550 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput561 net561 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[3] sky130_fd_sc_hd__buf_2
Xfanout1219 net96 VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__clkbuf_4
Xfanout1208 net151 VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__buf_4
Xoutput583 net583 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput594 net594 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_115_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_1__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs VGND VGND VPWR
+ VPWR clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_61_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4830_ net1200 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_178_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1973_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q _0974_ VGND VGND
+ VPWR VPWR _0975_ sky130_fd_sc_hd__nand2_1
X_4761_ net162 net1070 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3712_ net189 net9 net87 net101 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q VGND VGND VPWR VPWR
+ _0634_ sky130_fd_sc_hd__mux4_2
X_4692_ net1186 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3643_ net177 net69 net142 net213 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q VGND VGND VPWR VPWR
+ _0571_ sky130_fd_sc_hd__mux4_2
XFILLER_146_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3574_ net984 net998 net1020 net1001 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0506_ sky130_fd_sc_hd__mux4_1
X_2525_ net1257 net12 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__mux2_1
XFILLER_114_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2456_ net624 _0944_ _0981_ _0785_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__o22a_1
X_5244_ Tile_X0Y1_W6END[9] VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__clkbuf_2
X_5175_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR net526
+ sky130_fd_sc_hd__clkbuf_2
X_4126_ net1223 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2387_ _1088_ _1070_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__xnor2_4
XFILLER_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4057_ net1251 net1144 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_45_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3008_ net122 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__o21ba_1
XFILLER_24_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4959_ net1233 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_2
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput380 net380 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1027 net1028 VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__buf_2
Xfanout1038 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 VGND VGND VPWR VPWR
+ net1038 sky130_fd_sc_hd__buf_2
Xfanout1005 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 VGND VGND VPWR VPWR
+ net1005 sky130_fd_sc_hd__buf_8
XFILLER_126_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput391 net391 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_105_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1016 net1017 VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__buf_6
Xfanout1049 net1053 VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__buf_8
XFILLER_59_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2310_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q _1296_ VGND VGND
+ VPWR VPWR _1297_ sky130_fd_sc_hd__nand2_1
X_3290_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q _0240_ VGND VGND
+ VPWR VPWR _0241_ sky130_fd_sc_hd__or2_4
X_2241_ _0410_ _0302_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__mux2_1
XFILLER_2_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2172_ _1168_ _1166_ _1158_ _1167_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X sky130_fd_sc_hd__mux4_2
XFILLER_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4813_ net1182 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_44_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1956_ net662 _0829_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__nor2_1
XFILLER_21_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4744_ net1212 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4675_ net1206 net1096 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3626_ net974 net970 net989 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR
+ _0555_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3557_ _0475_ _0490_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ sky130_fd_sc_hd__mux2_4
XFILLER_163_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2508_ _1274_ _1456_ _1193_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__a21oi_1
Xinput108 Tile_X0Y0_W2MID[3] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlymetal6s2s_1
X_3488_ net76 net112 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q
+ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux2_1
XFILLER_102_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput119 Tile_X0Y1_E1END[0] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_4
X_2439_ net83 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__mux2_1
X_5158_ net161 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__buf_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4109_ net1238 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5089_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 VGND VGND VPWR VPWR net440
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2790_ _0199_ net93 net1 net1041 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q VGND VGND VPWR VPWR
+ _1703_ sky130_fd_sc_hd__mux4_1
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4460_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4391_ net48 net1151 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3411_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q _0355_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__o21ba_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3342_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q _0287_ _0291_
+ _0283_ _0281_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1
+ sky130_fd_sc_hd__o32a_4
X_3273_ net73 net81 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q VGND
+ VGND VPWR VPWR _0225_ sky130_fd_sc_hd__mux2_1
XFILLER_97_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2224_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q _1215_ _1216_
+ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__a21o_1
X_5012_ Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_6
XFILLER_38_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2155_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[12\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q
+ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__mux2_2
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2086_ _1079_ _1085_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__nand3_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2988_ _1855_ _1854_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 sky130_fd_sc_hd__mux2_1
XFILLER_159_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1939_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q _0941_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q
+ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__a21oi_2
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4727_ net1192 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4658_ net155 net1105 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput90 Tile_X0Y0_SS4END[5] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_4
XFILLER_162_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3609_ net198 net114 net1255 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__mux4_1
XFILLER_162_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4589_ net169 net1120 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_107_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3960_ _0096_ _0863_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q
+ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__a21bo_1
XFILLER_90_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2911_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q _1786_ _1789_
+ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__a21o_1
X_3891_ _0798_ _0799_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q
+ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__mux2_1
X_2842_ net1258 net1011 net1220 net1046 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q VGND VGND VPWR VPWR
+ _1748_ sky130_fd_sc_hd__mux4_1
XFILLER_148_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2773_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q _1688_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q
+ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__a21bo_1
XFILLER_129_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4512_ net1203 net1140 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_174_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4443_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.B3 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4374_ net1248 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3325_ _0273_ _0271_ _0052_ _0266_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__a211oi_4
XFILLER_112_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3256_ net1004 net1023 net617 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
X_2207_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q _1196_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_69_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3187_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR
+ VPWR _0142_ sky130_fd_sc_hd__inv_2
X_2138_ net26 net116 net77 _0468_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q VGND VGND VPWR VPWR
+ _1138_ sky130_fd_sc_hd__mux4_2
X_2069_ _1068_ _1056_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__xor2_4
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3110_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q VGND VGND VPWR
+ VPWR _0065_ sky130_fd_sc_hd__inv_1
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4090_ net29 net1133 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3041_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q VGND VGND VPWR VPWR
+ _1903_ sky130_fd_sc_hd__and3b_1
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4992_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 VGND VGND VPWR VPWR net343
+ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_74_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3943_ _0847_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__or2_4
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3874_ _0783_ _0781_ _0767_ _0782_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.A1 sky130_fd_sc_hd__mux4_2
XFILLER_176_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2825_ _1729_ _1730_ _1731_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q VGND VGND VPWR VPWR
+ _1732_ sky130_fd_sc_hd__a221o_1
XFILLER_176_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2756_ _0733_ net622 _0704_ net965 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q VGND VGND VPWR VPWR
+ _1673_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_135_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2687_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q _1631_ VGND VGND
+ VPWR VPWR _1632_ sky130_fd_sc_hd__or2_1
XFILLER_155_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4426_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0014_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ net1254 net1169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4288_ net52 net1083 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3308_ _0075_ _0257_ _0256_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__o211a_1
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3239_ _0189_ _0187_ _0192_ _0026_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ sky130_fd_sc_hd__a22o_4
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout970 net726 VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__buf_6
Xfanout992 net993 VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__buf_2
Xfanout981 net982 VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__buf_8
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2610_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q VGND VGND VPWR VPWR
+ _1564_ sky130_fd_sc_hd__mux2_1
X_3590_ _0076_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_11_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2541_ _1115_ _1480_ _1501_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__and3_4
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5260_ Tile_X0Y1_WW4END[15] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__clkbuf_2
X_2472_ _1414_ _1415_ _1447_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__a21boi_4
X_4211_ net1245 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5191_ Tile_X0Y0_S4END[14] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__buf_6
XFILLER_141_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4142_ net42 net1117 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_130_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4073_ net1232 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3024_ _1884_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q _1886_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q VGND VGND VPWR VPWR
+ _1887_ sky130_fd_sc_hd__o211a_1
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4975_ net1160 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_1
X_3926_ _0576_ _0740_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__nor2_1
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_178_Right_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3857_ net982 net996 net1018 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0769_ sky130_fd_sc_hd__mux4_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2808_ net1031 net721 _0652_ _1147_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q VGND VGND VPWR VPWR
+ _1718_ sky130_fd_sc_hd__mux4_1
XFILLER_149_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3788_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net16 net72 net108 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q VGND VGND VPWR VPWR
+ _0704_ sky130_fd_sc_hd__mux4_2
X_2739_ net621 net59 net1258 net1027 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _1660_ sky130_fd_sc_hd__mux4_1
XFILLER_117_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput551 net551 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput540 net540 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput562 net562 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[4] sky130_fd_sc_hd__buf_2
X_4409_ net1251 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput573 net573 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput584 net584 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput595 net595 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[5] sky130_fd_sc_hd__buf_2
Xfanout1209 net150 VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__buf_4
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1972_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 net228 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q
+ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__mux2_4
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4760_ net1194 net1070 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3711_ net206 net24 net78 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q VGND VGND VPWR VPWR
+ _0633_ sky130_fd_sc_hd__mux4_1
X_4691_ net1214 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3642_ net193 net89 net229 net706 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q VGND VGND VPWR VPWR
+ _0570_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_132_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3573_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q _0504_ VGND VGND
+ VPWR VPWR _0505_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2524_ net675 net192 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__mux2_1
XFILLER_114_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5243_ Tile_X0Y1_W6END[8] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__clkbuf_2
X_2455_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\] _1431_ net1057 VGND VGND VPWR VPWR
+ _1432_ sky130_fd_sc_hd__mux2_4
X_5174_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR net525
+ sky130_fd_sc_hd__buf_4
XFILLER_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2386_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\] _1366_ net1057 VGND VGND VPWR VPWR
+ _1367_ sky130_fd_sc_hd__mux2_4
X_4125_ net1222 net1124 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4056_ net1250 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3007_ net1067 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q VGND
+ VGND VPWR VPWR _1871_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_82_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4958_ net1235 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4889_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 VGND VGND VPWR VPWR net240
+ sky130_fd_sc_hd__clkbuf_2
X_3909_ _0815_ _0813_ _0115_ _0809_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput370 net370 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput381 net381 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[4] sky130_fd_sc_hd__buf_2
Xfanout1006 net1007 VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__buf_6
Xfanout1028 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 VGND VGND VPWR VPWR
+ net1028 sky130_fd_sc_hd__buf_2
XFILLER_120_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput392 net392 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1017 net1020 VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__buf_4
Xfanout1039 net1041 VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__buf_2
XFILLER_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2240_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q _1229_ _1231_
+ _1227_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ sky130_fd_sc_hd__a31o_4
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2171_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net15 net71 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q
+ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__mux4_1
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4812_ net1181 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1955_ _0906_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_1_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4743_ net1211 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4674_ net1205 net1096 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3625_ _0553_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q
+ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__a21bo_1
XFILLER_134_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3556_ _0489_ _0488_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux2_4
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2507_ net977 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 net1003 _1327_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 sky130_fd_sc_hd__mux4_2
Xinput109 Tile_X0Y0_W2MID[4] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
X_3487_ _0425_ _0044_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q
+ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
XFILLER_102_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5226_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 VGND VGND VPWR VPWR net577
+ sky130_fd_sc_hd__buf_4
XFILLER_102_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2438_ _1415_ _1414_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__xnor2_2
X_5157_ net160 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__buf_1
X_2369_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net226 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__mux2_4
XFILLER_56_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4108_ net1237 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5088_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 VGND VGND VPWR VPWR net439
+ sky130_fd_sc_hd__buf_1
X_4039_ net1229 net1144 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4390_ net49 net1151 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3410_ net176 net184 net1217 net130 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR VPWR
+ _0355_ sky130_fd_sc_hd__mux4_1
XFILLER_7_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3341_ _0057_ _0290_ _0289_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q
+ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__o211a_1
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3272_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q _0223_ VGND VGND
+ VPWR VPWR _0224_ sky130_fd_sc_hd__and2b_1
X_5011_ Tile_X0Y1_N4END[15] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_1
XFILLER_97_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2223_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q _1214_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q
+ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__o21ai_1
X_2154_ _1152_ _1148_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_127_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2085_ _1067_ _1071_ _1078_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_46_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2987_ net175 net1068 _0302_ net988 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q VGND VGND VPWR VPWR
+ _1855_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4726_ net1191 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1938_ _0940_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__inv_2
XFILLER_162_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4657_ net1190 net1105 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput91 Tile_X0Y0_SS4END[6] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_4
Xinput80 Tile_X0Y0_S4END[3] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3608_ _0537_ _0322_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q
+ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__mux2_4
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4588_ net170 net1120 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3539_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q _0473_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_55_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5209_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net566
+ sky130_fd_sc_hd__buf_6
XFILLER_123_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2910_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q _1788_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q
+ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__o21ai_1
XFILLER_176_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3890_ net72 net216 net84 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q VGND VGND VPWR VPWR
+ _0799_ sky130_fd_sc_hd__mux4_1
X_2841_ _1743_ _1745_ _1746_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q VGND VGND VPWR VPWR
+ _1747_ sky130_fd_sc_hd__o221a_1
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2772_ _1150_ _1512_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__mux2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4511_ net1201 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_174_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_91_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4442_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.B2 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4373_ net1247 net1160 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3324_ _0271_ _0273_ _0266_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a21o_1
XFILLER_112_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3255_ net617 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__o21ba_1
XFILLER_85_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2206_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q _1197_ _1198_
+ _1199_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q VGND VGND VPWR
+ VPWR _1200_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_69_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q VGND VGND VPWR
+ VPWR _0141_ sky130_fd_sc_hd__inv_2
X_2137_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q _1136_ VGND VGND
+ VPWR VPWR _1137_ sky130_fd_sc_hd__nor2_1
X_2068_ _1056_ _1068_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__nor2_1
XFILLER_41_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4709_ net150 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_Tile_X0Y1_UserCLK_regs Tile_X0Y1_UserCLK_regs VGND VGND VPWR VPWR clknet_0_Tile_X0Y1_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3040_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ _1901_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q VGND VGND VPWR
+ VPWR _1902_ sky130_fd_sc_hd__o211a_1
XFILLER_48_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4991_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 VGND VGND VPWR VPWR net342
+ sky130_fd_sc_hd__buf_4
XFILLER_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3942_ _0842_ _0846_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__nor2_1
XFILLER_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3873_ net133 net223 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__mux4_2
XFILLER_176_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2824_ net1011 net1046 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2755_ _1669_ _1671_ _1672_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_135_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2686_ net1046 net1026 net1050 net1042 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _1631_ sky130_fd_sc_hd__mux4_1
XFILLER_132_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4425_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0013_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_4356_ net1243 net1169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3307_ net979 net1019 net984 net1002 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q VGND VGND VPWR VPWR
+ _0257_ sky130_fd_sc_hd__mux4_1
XFILLER_48_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4287_ net1224 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_104_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3238_ _0190_ _0191_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q
+ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
XFILLER_39_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3169_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q VGND VGND VPWR
+ VPWR _0124_ sky130_fd_sc_hd__inv_1
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_138_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_147_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout993 net994 VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__clkbuf_2
Xfanout971 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 VGND VGND VPWR VPWR net971
+ sky130_fd_sc_hd__buf_4
Xfanout982 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 VGND VGND VPWR VPWR net982
+ sky130_fd_sc_hd__buf_8
XFILLER_64_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2540_ _1500_ net1058 _1482_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__a21oi_2
XFILLER_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2471_ _1416_ _1446_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__or2_4
X_4210_ net1244 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5190_ Tile_X0Y0_S4END[13] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__buf_6
X_4141_ net43 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_130_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4072_ net1231 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_182_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3023_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q _1885_ VGND VGND
+ VPWR VPWR _1886_ sky130_fd_sc_hd__nand2_1
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4974_ net1169 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_141_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3925_ _0450_ _0740_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__nor2_1
XFILLER_51_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3856_ net972 net986 net990 net976 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0768_ sky130_fd_sc_hd__mux4_1
XFILLER_166_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2807_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q _1712_ _1717_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 sky130_fd_sc_hd__o21ba_1
X_3787_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net107 net15 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q
+ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__mux4_2
XFILLER_164_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2738_ _1656_ _1658_ _1659_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 sky130_fd_sc_hd__o22a_1
XFILLER_117_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4408_ net31 net1151 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2669_ _1453_ _1454_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__xor2_1
XFILLER_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput530 net530 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput552 net552 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput541 net541 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput563 net563 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput574 net574 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput585 net585 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput596 net596 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[6] sky130_fd_sc_hd__buf_2
X_4339_ net1245 net1169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1971_ _0970_ _0971_ _0972_ _0126_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__a221o_1
X_3710_ _0632_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2
+ sky130_fd_sc_hd__clkinv_2
XFILLER_81_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4690_ net1202 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3641_ _0110_ _0196_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q
+ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__o21ba_1
X_3572_ net974 net970 net989 net994 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0504_ sky130_fd_sc_hd__mux4_1
X_2523_ _1485_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q
+ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__a21bo_1
XFILLER_114_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5242_ Tile_X0Y1_W6END[7] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__clkbuf_2
X_2454_ Tile_X0Y1_DSP_bot.C1 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[1\] net1063 VGND
+ VGND VPWR VPWR _1431_ sky130_fd_sc_hd__mux2_2
XFILLER_102_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5173_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR net524
+ sky130_fd_sc_hd__buf_6
X_2385_ Tile_X0Y1_DSP_bot.C5 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[5\] net1063 VGND
+ VGND VPWR VPWR _1366_ sky130_fd_sc_hd__mux2_2
X_4124_ net1221 net1124 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput1 Tile_X0Y0_E1END[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_6
XFILLER_68_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4055_ net1249 net1144 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_39_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3006_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q _1865_ _1870_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 sky130_fd_sc_hd__o21a_1
XFILLER_91_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4957_ net1237 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_2
XFILLER_61_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4888_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 VGND VGND VPWR VPWR net239
+ sky130_fd_sc_hd__buf_2
X_3908_ _0813_ _0815_ _0809_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ sky130_fd_sc_hd__a21o_1
XFILLER_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3839_ _0578_ _0579_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__or2_1
XFILLER_117_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput371 net371 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput360 net360 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput382 net382 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[5] sky130_fd_sc_hd__buf_2
Xfanout1007 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 VGND VGND VPWR VPWR
+ net1007 sky130_fd_sc_hd__buf_8
Xfanout1029 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 VGND VGND VPWR VPWR
+ net1029 sky130_fd_sc_hd__buf_8
Xoutput393 net393 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_105_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1018 net1020 VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__buf_8
XFILLER_59_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2170_ net207 net79 net7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q VGND VGND VPWR VPWR
+ _1167_ sky130_fd_sc_hd__mux4_1
XFILLER_65_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4811_ net1180 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1954_ _0709_ _0785_ net624 _0661_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__o22ai_2
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4742_ net1210 net1079 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4673_ net1204 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3624_ net734 net1015 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__mux2_2
XFILLER_174_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3555_ net185 net5 net61 net118 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q VGND VGND VPWR VPWR
+ _0489_ sky130_fd_sc_hd__mux4_2
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3486_ _0425_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7
+ sky130_fd_sc_hd__inv_1
X_2506_ _1473_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 sky130_fd_sc_hd__mux2_4
XFILLER_142_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2437_ _1083_ _1082_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__xor2_4
X_5225_ net217 VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_102_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5156_ net159 VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__buf_1
X_2368_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q _1350_ VGND VGND
+ VPWR VPWR _1351_ sky130_fd_sc_hd__and2b_1
XFILLER_56_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4107_ net1235 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2299_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1284_ _1286_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q VGND VGND VPWR VPWR
+ _1287_ sky130_fd_sc_hd__o211a_1
X_5087_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 VGND VGND VPWR VPWR net438
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4038_ net49 net1143 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_111_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3340_ net99 net118 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q VGND
+ VGND VPWR VPWR _0290_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5010_ Tile_X0Y1_N4END[14] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_1
XFILLER_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3271_ net181 net127 net1218 net1216 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q VGND VGND VPWR VPWR
+ _0223_ sky130_fd_sc_hd__mux4_1
X_2222_ net997 net693 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__mux2_1
X_2153_ _1150_ _1151_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__mux2_4
Xclone130 net999 VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2084_ _1080_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__and2_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2986_ _1852_ _1853_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q
+ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__mux2_1
XFILLER_159_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1937_ net188 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net224
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q
+ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__mux4_2
X_4725_ net1188 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4656_ net1185 net1105 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput81 Tile_X0Y0_S4END[4] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_4
Xinput70 Tile_X0Y0_S2MID[1] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_8
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3607_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 net109 net17 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q
+ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__mux4_2
X_4587_ net1180 net1120 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput92 Tile_X0Y0_SS4END[7] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_4
XFILLER_162_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3538_ net70 net106 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q VGND
+ VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
XFILLER_115_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3469_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q _0408_ VGND VGND
+ VPWR VPWR _0409_ sky130_fd_sc_hd__nand2b_1
XFILLER_88_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5208_ Tile_X0Y0_SS4END[15] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__buf_6
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5139_ net1182 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_4
XFILLER_123_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2840_ net1006 net1031 net1021 net1054 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q VGND VGND VPWR VPWR
+ _1746_ sky130_fd_sc_hd__mux4_1
XFILLER_92_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2771_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q _1686_ VGND
+ VGND VPWR VPWR _1687_ sky130_fd_sc_hd__and2b_1
XFILLER_156_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4510_ net1200 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4441_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.B1 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4372_ net1246 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3323_ _0054_ _0272_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__o21ba_1
XFILLER_152_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3254_ net1034 net617 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__nand2b_1
XFILLER_85_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2205_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q net693 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_69_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR
+ VPWR _0140_ sky130_fd_sc_hd__inv_2
Xfanout1190 net165 VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__clkbuf_4
X_2136_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q _1133_ _1135_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q VGND VGND VPWR VPWR
+ _1136_ sky130_fd_sc_hd__o211a_1
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2067_ _1067_ _1065_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__and2_4
XFILLER_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2969_ _0818_ _1391_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__mux2_1
X_4708_ net151 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4639_ net156 net1105 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4990_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 VGND VGND VPWR VPWR net341
+ sky130_fd_sc_hd__clkbuf_2
X_3941_ _0842_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__and2_1
XFILLER_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3872_ net143 net83 net220 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q VGND VGND VPWR VPWR
+ _0782_ sky130_fd_sc_hd__mux4_2
XFILLER_176_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2823_ net1257 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_14_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2754_ _0243_ net58 net2 net1038 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q VGND VGND VPWR VPWR
+ _1672_ sky130_fd_sc_hd__mux4_1
XFILLER_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2685_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q _1629_ _1628_
+ _0047_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__a211o_1
X_4424_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0012_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4355_ net1230 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3306_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q _0255_ VGND VGND
+ VPWR VPWR _0256_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4286_ net1223 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3237_ net79 net87 net99 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0191_ sky130_fd_sc_hd__mux4_1
XFILLER_104_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3168_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q VGND VGND VPWR
+ VPWR _0123_ sky130_fd_sc_hd__inv_2
XFILLER_73_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2119_ net1011 net1046 net1028 net1052 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR
+ _1120_ sky130_fd_sc_hd__mux4_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3099_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR
+ VPWR _0054_ sky130_fd_sc_hd__inv_2
XFILLER_120_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout983 net984 VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__buf_2
Xfanout972 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 VGND VGND VPWR VPWR net972
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout994 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 VGND VGND VPWR VPWR net994
+ sky130_fd_sc_hd__buf_12
XFILLER_161_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2470_ _1432_ _1435_ _1445_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__a21oi_2
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4140_ net44 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_130_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4071_ net1229 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_182_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3022_ _1410_ _1349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__mux2_1
XFILLER_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4973_ net1077 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_62_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3924_ _0492_ _0829_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__or2_4
X_3855_ net188 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net224
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q
+ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__mux4_2
XFILLER_164_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2806_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q _1716_ _1714_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q VGND VGND VPWR VPWR
+ _1717_ sky130_fd_sc_hd__o211a_1
X_3786_ _0702_ _0699_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 sky130_fd_sc_hd__mux2_4
XFILLER_164_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2737_ _0243_ net94 net2 net1037 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q VGND VGND VPWR VPWR
+ _1659_ sky130_fd_sc_hd__mux4_1
XFILLER_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput520 net520 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[0] sky130_fd_sc_hd__buf_2
X_2668_ _1615_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 sky130_fd_sc_hd__mux2_4
X_4407_ net1249 net1152 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput531 net531 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput542 net542 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput553 net553 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[10] sky130_fd_sc_hd__buf_2
X_2599_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6
+ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__nand2_1
Xoutput564 net564 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput575 net575 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput586 net586 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[6] sky130_fd_sc_hd__buf_2
X_4338_ net37 net1169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput597 net597 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_115_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4269_ net1238 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1970_ net137 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__mux2_1
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3640_ _0559_ _0558_ _0567_ _0109_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q
+ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__a221o_1
X_3571_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q _0501_ _0503_
+ _0496_ _0497_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ sky130_fd_sc_hd__o32a_4
X_2522_ net1043 net1032 net1038 net1022 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q VGND VGND VPWR VPWR
+ _1485_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_93_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5241_ Tile_X0Y1_W6END[6] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_2
X_2453_ _1430_ _1428_ _1423_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C1 sky130_fd_sc_hd__a21oi_2
XFILLER_114_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5172_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR net523
+ sky130_fd_sc_hd__buf_1
X_2384_ _1362_ _1365_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C5 sky130_fd_sc_hd__mux2_4
XFILLER_110_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4123_ net1253 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput2 Tile_X0Y0_E1END[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
X_4054_ net1248 net1144 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_166_Left_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3005_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q _1866_ _1869_
+ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__a21o_1
XFILLER_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4956_ net1238 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_2
XFILLER_177_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4887_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 VGND VGND VPWR VPWR net238
+ sky130_fd_sc_hd__buf_1
X_3907_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q _0814_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__o21ba_1
XFILLER_177_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_175_Left_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3838_ _0748_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__nand2b_4
X_3769_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q _0686_ VGND VGND
+ VPWR VPWR _0687_ sky130_fd_sc_hd__nor2_1
XFILLER_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput361 net361 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput350 net350 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[3] sky130_fd_sc_hd__buf_2
XFILLER_105_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput372 net372 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput383 net383 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[6] sky130_fd_sc_hd__buf_2
Xfanout1008 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 VGND VGND VPWR VPWR
+ net1008 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput394 net394 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1019 net1020 VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__buf_2
XFILLER_113_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4810_ net1179 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_178_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1953_ _0946_ _0950_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__xnor2_2
X_4741_ net150 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_14_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4672_ net1203 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3623_ _0107_ net998 _0551_ _0108_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__o211a_1
XFILLER_174_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3554_ net197 net1256 net77 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q
+ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux4_2
X_3485_ _0415_ _0417_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__a21oi_2
X_2505_ _1455_ _1472_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__xor2_1
XFILLER_102_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5224_ net216 VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__buf_1
X_2436_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\] _1413_ net1057 VGND VGND VPWR VPWR
+ _1414_ sky130_fd_sc_hd__mux2_4
X_5155_ net158 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__buf_1
XFILLER_29_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2367_ net190 net136 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__mux2_1
XFILLER_56_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4106_ net1234 net1126 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2298_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1285_ VGND VGND
+ VPWR VPWR _1286_ sky130_fd_sc_hd__nand2_1
X_5086_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 VGND VGND VPWR VPWR net437
+ sky130_fd_sc_hd__buf_1
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4037_ net27 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4939_ net54 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_2
XFILLER_177_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _0221_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a21bo_1
X_2221_ _1213_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__inv_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone120 net1035 VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__buf_6
X_2152_ net710 net74 net18 net110 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q VGND VGND VPWR VPWR
+ _1151_ sky130_fd_sc_hd__mux4_2
XFILLER_93_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2083_ _1082_ _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__nor2_1
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4724_ net1186 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2985_ _0940_ _1347_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__mux2_1
XFILLER_159_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1936_ _0937_ _0936_ _0938_ _0124_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__a221o_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4655_ net1184 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput82 Tile_X0Y0_S4END[5] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_4
Xinput71 Tile_X0Y0_S2MID[2] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_4
Xinput60 Tile_X0Y0_S1END[3] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
X_3606_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 VGND VGND VPWR VPWR _0536_
+ sky130_fd_sc_hd__inv_1
X_4586_ net1179 net1120 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput93 Tile_X0Y0_W1END[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
X_3537_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q _0471_ VGND VGND
+ VPWR VPWR _0472_ sky130_fd_sc_hd__and2b_1
XFILLER_130_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3468_ net1039 _0407_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q
+ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux2_1
XFILLER_88_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5207_ Tile_X0Y0_SS4END[14] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__buf_6
X_3399_ _0343_ _0344_ _0064_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__mux2_1
X_2419_ net186 net132 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q
+ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__mux2_1
XFILLER_123_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5138_ net1183 VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__buf_2
XFILLER_29_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5069_ Tile_X0Y0_WW4END[4] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkbuf_2
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2770_ net721 _0652_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__mux2_1
XFILLER_129_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4440_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.B0 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4371_ net36 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3322_ net58 net66 net60 net94 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q VGND VGND VPWR VPWR
+ _0272_ sky130_fd_sc_hd__mux4_1
XFILLER_112_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3253_ _0037_ _0205_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q
+ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__o21ba_1
X_3184_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q VGND VGND VPWR
+ VPWR _0139_ sky130_fd_sc_hd__inv_1
XFILLER_112_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2204_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q net734 VGND VGND
+ VPWR VPWR _1198_ sky130_fd_sc_hd__and2b_1
X_2135_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q _1134_ VGND VGND
+ VPWR VPWR _1135_ sky130_fd_sc_hd__nand2_1
Xfanout1180 net171 VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__buf_4
Xfanout1191 net164 VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2066_ _1060_ _1065_ _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nand3b_4
XTAP_TAPCELL_ROW_144_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2968_ net176 net1217 net1067 net994 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q VGND VGND VPWR VPWR
+ _1839_ sky130_fd_sc_hd__mux4_1
XFILLER_147_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1919_ net973 net968 net987 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR
+ _0923_ sky130_fd_sc_hd__mux4_2
X_4707_ net1206 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2899_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q _1777_ _1779_
+ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__a21bo_1
X_4638_ net157 net1105 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4569_ net1195 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_9_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone41 _0298_ _0295_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__mux2_4
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone74 net704 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkbuf_1
XFILLER_175_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3940_ _0844_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__or2_1
XFILLER_90_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3871_ net201 net71 net125 net215 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q VGND VGND VPWR VPWR
+ _0781_ sky130_fd_sc_hd__mux4_2
XFILLER_176_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2822_ net1219 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q VGND
+ VGND VPWR VPWR _1729_ sky130_fd_sc_hd__nand2b_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2753_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q _1670_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2684_ net98 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q VGND
+ VGND VPWR VPWR _1629_ sky130_fd_sc_hd__mux2_1
XFILLER_144_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4423_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs _0011_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4354_ net1227 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3305_ net973 net968 net988 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR VPWR
+ _0255_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_6_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4285_ net1222 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3236_ net207 net1 net25 net1256 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0190_ sky130_fd_sc_hd__mux4_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3167_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR
+ VPWR _0122_ sky130_fd_sc_hd__inv_2
XFILLER_39_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3098_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR
+ VPWR _0053_ sky130_fd_sc_hd__inv_2
X_2118_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\]
+ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__nand2_1
XFILLER_81_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ _1046_ _1048_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__nand2_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout973 net974 VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__buf_2
Xfanout995 net999 VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__buf_2
Xfanout984 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 VGND VGND VPWR VPWR net984
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_79_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4070_ net1228 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3021_ _0662_ _0819_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _1884_ sky130_fd_sc_hd__mux2_2
XFILLER_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4972_ net1084 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3923_ _0827_ _0828_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__nand2_8
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3854_ _0765_ _0580_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__xnor2_2
X_2805_ _1715_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__inv_1
X_3785_ _0701_ _0700_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q
+ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__mux2_1
X_2736_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q _1657_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__a21bo_1
XFILLER_117_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput510 net510 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[4] sky130_fd_sc_hd__buf_2
X_2667_ _1443_ _1444_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__xnor2_2
XFILLER_105_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4406_ net1248 net1152 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput521 net521 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput532 net532 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput543 net543 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput554 net554 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[11] sky130_fd_sc_hd__buf_6
X_2598_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q VGND VGND VPWR VPWR
+ _1553_ sky130_fd_sc_hd__mux2_4
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_97_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput576 net576 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput565 net565 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput587 net587 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[7] sky130_fd_sc_hd__buf_2
X_4337_ net39 net1170 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput598 net598 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[8] sky130_fd_sc_hd__buf_2
X_4268_ net1237 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3219_ _0171_ _0170_ _0172_ _0035_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a22o_4
X_4199_ net1229 net1101 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_85_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3570_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q _0502_ VGND VGND
+ VPWR VPWR _0503_ sky130_fd_sc_hd__and2b_1
X_2521_ _0094_ _1483_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__and2_1
XFILLER_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5240_ Tile_X0Y1_W6END[5] VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2452_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q
+ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__a21oi_1
X_5171_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR net522
+ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2383_ _1364_ _1363_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__mux2_4
XFILLER_122_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4122_ net1252 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4053_ net1247 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 Tile_X0Y0_E1END[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_39_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3004_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q _1868_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q
+ VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__o21ai_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4955_ net42 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_1
XFILLER_101_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3906_ net174 net182 net120 net128 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0814_ sky130_fd_sc_hd__mux4_1
XFILLER_51_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4886_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 VGND VGND VPWR VPWR net237
+ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_22_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3837_ _0681_ _0732_ _0747_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__or3b_1
X_3768_ _0243_ net190 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__mux2_1
X_2719_ net1004 _0526_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 _0520_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_150_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3699_ net1010 net724 net1053 net1041 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0622_ sky130_fd_sc_hd__mux4_1
XFILLER_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput351 net351 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[4] sky130_fd_sc_hd__buf_6
Xoutput362 net362 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput340 net340 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_160_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput384 net384 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput373 net373 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[11] sky130_fd_sc_hd__buf_2
Xfanout1009 net1010 VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__buf_8
XFILLER_120_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput395 net395 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1952_ _0952_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__nor2_1
X_4740_ net151 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_14_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4671_ net156 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3622_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q net984 VGND VGND
+ VPWR VPWR _0551_ sky130_fd_sc_hd__or2_1
XFILLER_174_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3553_ _0051_ _0483_ _0487_ _0479_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1
+ sky130_fd_sc_hd__a31o_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2504_ _1273_ _1275_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__nor2_2
X_3484_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q _0423_ _0422_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q VGND VGND VPWR VPWR
+ _0424_ sky130_fd_sc_hd__o211a_1
X_5223_ net705 VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__buf_1
X_2435_ Tile_X0Y1_DSP_bot.C2 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[2\] net1063 VGND
+ VGND VPWR VPWR _1413_ sky130_fd_sc_hd__mux2_4
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5154_ net1200 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkbuf_2
X_4105_ net1232 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2366_ net135 net225 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q
+ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__mux4_2
XFILLER_110_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2297_ net1019 net1014 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__mux2_1
X_5085_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 VGND VGND VPWR VPWR net436
+ sky130_fd_sc_hd__buf_1
XFILLER_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4036_ net38 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_16_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ net53 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4869_ net1209 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ net979 net984 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__mux2_1
XFILLER_87_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2151_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 net109 net73 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q
+ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_49_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2082_ _1075_ _1044_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__xnor2_4
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2984_ net997 _0767_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__mux2_1
X_4723_ net145 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1935_ net187 net133 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q
+ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4654_ net1183 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput72 Tile_X0Y0_S2MID[3] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_8
Xinput61 Tile_X0Y0_S2END[0] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_2
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput50 Tile_X0Y0_FrameData[3] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
X_3605_ _0535_ _0533_ _0507_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4
+ sky130_fd_sc_hd__a21o_4
X_4585_ net1213 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput83 Tile_X0Y0_S4END[6] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput94 Tile_X0Y0_W1END[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_4
X_3536_ net689 net14 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q VGND
+ VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_1
XFILLER_115_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5206_ Tile_X0Y0_SS4END[13] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__buf_6
XFILLER_130_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3467_ net689 net70 net14 net106 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q VGND VGND VPWR VPWR
+ _0407_ sky130_fd_sc_hd__mux4_2
X_3398_ net187 net1 net199 net7 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q VGND VGND VPWR VPWR
+ _0344_ sky130_fd_sc_hd__mux4_1
XFILLER_130_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2418_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q _1397_ VGND VGND
+ VPWR VPWR _1398_ sky130_fd_sc_hd__nand2_1
XFILLER_96_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5137_ net1184 VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_24_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2349_ net185 net131 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__mux2_1
X_5068_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 VGND VGND VPWR VPWR net410
+ sky130_fd_sc_hd__buf_4
XFILLER_123_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4019_ net1245 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_123_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4370_ net37 net1160 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3321_ _0267_ _0053_ _0268_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__a31o_4
XFILLER_152_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3252_ net57 net61 net93 net1220 net617 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__mux4_1
XFILLER_85_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2203_ net979 net998 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__mux2_1
X_3183_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q VGND VGND VPWR
+ VPWR _0138_ sky130_fd_sc_hd__inv_1
X_2134_ net70 net106 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q
+ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__mux2_1
Xfanout1170 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__buf_2
XFILLER_78_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1181 net170 VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__buf_4
Xfanout1192 net163 VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__clkbuf_4
XFILLER_81_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2065_ _1049_ _1064_ _1063_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__o21bai_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2967_ _1835_ _1838_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 sky130_fd_sc_hd__mux2_1
XFILLER_147_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4706_ net1205 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1918_ _0921_ _0173_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2898_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q _0662_ _1778_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR
+ _1779_ sky130_fd_sc_hd__a211o_1
XFILLER_162_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4637_ net1199 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4568_ net1193 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4499_ net145 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3519_ net1215 net214 net90 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q VGND VGND VPWR VPWR
+ _0455_ sky130_fd_sc_hd__mux4_1
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_108_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone75 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 VGND VGND VPWR VPWR net692
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone97 net1001 VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__buf_8
XFILLER_175_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3870_ _0780_ _0777_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 sky130_fd_sc_hd__mux2_4
XFILLER_176_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2821_ _1725_ _1727_ _1728_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_14_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2752_ _1512_ _0710_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q
+ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__mux2_1
XFILLER_129_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2683_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q _1627_ VGND VGND
+ VPWR VPWR _1628_ sky130_fd_sc_hd__and2b_1
X_4422_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs _0010_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4353_ net1226 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3304_ _0253_ _0252_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q
+ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
X_4284_ net1221 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3235_ _0025_ _0188_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__o21a_1
XFILLER_58_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3166_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q VGND VGND VPWR
+ VPWR _0121_ sky130_fd_sc_hd__inv_2
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2117_ _0432_ _1116_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__xor2_1
X_3097_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q VGND VGND VPWR
+ VPWR _0052_ sky130_fd_sc_hd__inv_2
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2048_ _1042_ _1047_ _1048_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__and3_4
XFILLER_54_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3999_ _0901_ _0902_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nor2_1
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout974 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 VGND VGND VPWR VPWR net974
+ sky130_fd_sc_hd__buf_2
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout985 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 VGND VGND VPWR VPWR net985
+ sky130_fd_sc_hd__buf_8
Xfanout963 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr VGND VGND VPWR VPWR net963
+ sky130_fd_sc_hd__buf_2
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net999 VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__buf_8
XFILLER_45_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3020_ _0157_ _1874_ _1879_ _1883_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0
+ sky130_fd_sc_hd__a31o_1
XFILLER_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4971_ net1091 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3922_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\] net1062 VGND VGND VPWR VPWR _0828_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3853_ _0764_ _0763_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__nor2_2
XFILLER_149_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2804_ net740 _0733_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q
+ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__mux2_1
XFILLER_157_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3784_ net180 net196 net120 net126 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0701_ sky130_fd_sc_hd__mux4_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2735_ _1512_ _0737_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q
+ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__mux2_1
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2666_ _1614_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 sky130_fd_sc_hd__mux2_4
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput500 net500 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput511 net511 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[5] sky130_fd_sc_hd__buf_2
XFILLER_132_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4405_ net1247 net1152 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput522 net522 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput533 net533 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput544 net544 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[2] sky130_fd_sc_hd__buf_2
X_2597_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q _1551_ _1550_
+ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__o21a_1
X_4336_ net1241 net1169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput566 net566 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[8] sky130_fd_sc_hd__buf_4
Xoutput555 net555 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput577 net577 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[5] sky130_fd_sc_hd__buf_6
XFILLER_115_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput588 net588 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput599 net599 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[9] sky130_fd_sc_hd__buf_2
X_4267_ net1235 net1084 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4198_ net1228 net1101 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3218_ net195 net125 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q
+ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
X_3149_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q VGND VGND VPWR
+ VPWR _0104_ sky130_fd_sc_hd__inv_1
XFILLER_27_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2520_ net1012 net1047 net1027 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR VPWR
+ _1483_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_93_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2451_ net188 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net224
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q
+ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__mux4_2
X_5170_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 VGND VGND VPWR VPWR net521
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2382_ net180 net126 net89 net216 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q VGND VGND VPWR VPWR
+ _1364_ sky130_fd_sc_hd__mux4_1
X_4121_ net1251 net1124 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4052_ net35 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput4 Tile_X0Y0_E1END[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_3003_ _1867_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__inv_1
XFILLER_91_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4954_ net1240 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3905_ _0811_ _0810_ _0812_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ _0116_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__a221o_1
XFILLER_177_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4885_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 VGND VGND VPWR VPWR net236
+ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_22_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3836_ _0681_ _0732_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__o21ba_4
X_3767_ _0684_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q VGND VGND
+ VPWR VPWR _0685_ sky130_fd_sc_hd__nand2_2
XFILLER_145_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2718_ net737 _0407_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 _0398_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3698_ _0601_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__nor2_4
Xoutput330 net330 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput341 net341 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput352 net352 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[5] sky130_fd_sc_hd__buf_2
X_2649_ net57 net61 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q VGND
+ VGND VPWR VPWR _1602_ sky130_fd_sc_hd__mux2_1
XFILLER_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput385 net385 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput363 net363 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput374 net374 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput396 net396 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_86_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4319_ net1224 net1076 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1951_ _0904_ _0951_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__and2b_1
XFILLER_14_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4670_ net157 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3621_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q _0549_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__o21ba_1
XFILLER_174_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3552_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q _0486_ _0485_
+ _0050_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__a211o_1
XFILLER_127_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2503_ _1471_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 sky130_fd_sc_hd__mux2_4
X_3483_ net973 net968 net987 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR VPWR
+ _0423_ sky130_fd_sc_hd__mux4_1
XFILLER_130_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5222_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR net573
+ sky130_fd_sc_hd__buf_1
X_2434_ _1412_ _1409_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C2 sky130_fd_sc_hd__mux2_4
XFILLER_142_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5153_ net1201 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkbuf_2
X_2365_ _1347_ _1346_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__mux2_4
X_4104_ net1231 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5084_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR net426
+ sky130_fd_sc_hd__buf_2
XFILLER_110_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2296_ _1283_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__inv_1
XFILLER_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4035_ net1230 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4937_ net1225 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_2
X_4868_ net1208 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_177_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3819_ _0730_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__nor2_1
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4799_ net156 net1166 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2150_ _0536_ _0081_ _0030_ _0158_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q VGND VGND VPWR VPWR
+ _1149_ sky130_fd_sc_hd__mux4_2
Xclone133 net1025 VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__buf_6
XFILLER_93_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2081_ _1073_ _1081_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__nand2_4
XFILLER_179_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2983_ _1848_ _1851_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 sky130_fd_sc_hd__mux2_1
X_4722_ net1202 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1934_ net223 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q
+ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__o21a_1
XFILLER_159_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput40 Tile_X0Y0_FrameData[21] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
XFILLER_147_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4653_ net1182 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput62 Tile_X0Y0_S2END[1] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
Xinput73 Tile_X0Y0_S2MID[4] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_4
XFILLER_174_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput51 Tile_X0Y0_FrameData[4] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
X_3604_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q _0534_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__o21ba_1
X_4584_ net1212 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput84 Tile_X0Y0_S4END[7] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_4
XFILLER_162_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput95 Tile_X0Y0_W1END[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
X_3535_ net69 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q
+ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__o211a_1
XFILLER_115_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3466_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q VGND VGND VPWR VPWR
+ _0406_ sky130_fd_sc_hd__o21ai_4
XFILLER_170_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5205_ Tile_X0Y0_SS4END[12] VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__buf_6
XFILLER_115_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2417_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net222 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q
+ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3397_ net21 net99 net63 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q VGND VGND VPWR VPWR
+ _0343_ sky130_fd_sc_hd__mux4_1
XFILLER_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5136_ net1185 VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_2
X_2348_ net221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q
+ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__o21a_1
X_5067_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 VGND VGND VPWR VPWR net409
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_123_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2279_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR
+ _1268_ sky130_fd_sc_hd__o21ai_1
XFILLER_177_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4018_ net1244 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3320_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q _0269_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q
+ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a21o_1
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3251_ _0201_ _0200_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__a21o_1
XFILLER_85_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2202_ _1195_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__inv_1
X_3182_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR
+ VPWR _0137_ sky130_fd_sc_hd__inv_1
Xfanout1160 net1161 VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2133_ _1132_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__inv_1
Xfanout1182 net169 VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__buf_4
Xfanout1171 net1173 VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__clkbuf_2
Xfanout1193 net1194 VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__clkbuf_4
X_2064_ _1049_ _1064_ _1063_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_144_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2966_ _1836_ _1837_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q
+ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__mux2_1
X_4705_ net1204 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_60_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1917_ net179 net125 net71 net233 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q VGND VGND VPWR VPWR
+ _0921_ sky130_fd_sc_hd__mux4_2
X_2897_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q net733 VGND
+ VGND VPWR VPWR _1778_ sky130_fd_sc_hd__nor2_1
XFILLER_147_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4636_ net1198 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4567_ net1192 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4498_ net155 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3518_ net178 net194 net1217 net124 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _0454_ sky130_fd_sc_hd__mux4_1
X_3449_ _0091_ _0390_ _0389_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q
+ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__o211a_1
XFILLER_103_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5119_ Tile_X0Y1_EE4END[6] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone76 net742 VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__clkbuf_1
XFILLER_175_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone98 net981 VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__buf_6
XFILLER_175_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput230 Tile_X0Y1_W6END[1] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2820_ _0243_ net94 net58 net1037 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q VGND VGND VPWR VPWR
+ _1728_ sky130_fd_sc_hd__mux4_1
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2751_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q _1149_ _1668_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q VGND VGND VPWR VPWR
+ _1669_ sky130_fd_sc_hd__a211oi_1
XFILLER_129_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2682_ net62 net78 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q VGND
+ VGND VPWR VPWR _1627_ sky130_fd_sc_hd__mux2_1
XFILLER_129_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4421_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs _0009_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4352_ net1225 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3303_ net192 net68 net12 net115 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q VGND VGND VPWR VPWR
+ _0253_ sky130_fd_sc_hd__mux4_2
X_4283_ net28 net1083 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3234_ net1034 net1004 net1029 net1023 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0188_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_146_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3165_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q VGND VGND VPWR
+ VPWR _0120_ sky130_fd_sc_hd__inv_2
XFILLER_39_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2116_ _1116_ _0432_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__nand2b_4
X_3096_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q VGND VGND VPWR
+ VPWR _0051_ sky130_fd_sc_hd__inv_1
XFILLER_81_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2047_ _1043_ _1045_ _1046_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__nand3_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3998_ _0899_ _0900_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__nor2_1
XFILLER_13_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2949_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q _1822_ _1821_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q VGND VGND VPWR VPWR
+ _1823_ sky130_fd_sc_hd__o211a_1
XFILLER_175_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4619_ net171 net1112 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_112_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout975 net977 VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__buf_8
Xfanout986 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 VGND VGND VPWR VPWR net986
+ sky130_fd_sc_hd__buf_6
Xfanout964 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr VGND VGND VPWR VPWR net964
+ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_164_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 net998 VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__buf_2
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4970_ net1100 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_62_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3921_ _0820_ _0826_ _0804_ net1061 VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__a211o_4
X_3852_ _0748_ _0753_ _0762_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__o21ba_1
X_2803_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q _1713_ VGND VGND
+ VPWR VPWR _1714_ sky130_fd_sc_hd__nand2_1
XFILLER_164_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3783_ net1215 net72 net216 net232 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0700_ sky130_fd_sc_hd__mux4_1
XFILLER_157_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2734_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q _1149_ _1655_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q VGND VGND VPWR VPWR
+ _1656_ sky130_fd_sc_hd__a211oi_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2665_ _1562_ _1560_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__xnor2_1
Xoutput501 net501 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[25] sky130_fd_sc_hd__buf_2
X_2596_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q VGND VGND VPWR VPWR
+ _1551_ sky130_fd_sc_hd__mux2_1
X_4404_ net1246 net1152 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput523 net523 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput534 net534 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput545 net545 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput512 net512 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[6] sky130_fd_sc_hd__buf_2
X_4335_ net1240 net1169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput567 net567 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[9] sky130_fd_sc_hd__buf_6
Xoutput556 net556 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[13] sky130_fd_sc_hd__buf_6
Xoutput578 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR
+ Tile_X0Y1_W2BEG[6] sky130_fd_sc_hd__buf_6
XFILLER_59_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput589 net589 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[10] sky130_fd_sc_hd__buf_2
X_4266_ net1234 net1084 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4197_ net27 net1109 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3217_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q net220 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q
+ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__o21a_1
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3148_ net225 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_1
XFILLER_54_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3079_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q VGND VGND VPWR
+ VPWR _0034_ sky130_fd_sc_hd__inv_2
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire617 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q VGND VGND VPWR
+ VPWR net617 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2450_ _1425_ _1424_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q
+ _1427_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q VGND VGND VPWR
+ VPWR _1428_ sky130_fd_sc_hd__a311o_1
XFILLER_5_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2381_ net195 net215 net91 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR
+ _1363_ sky130_fd_sc_hd__mux4_2
X_4120_ net1250 net1124 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4051_ net1245 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput5 Tile_X0Y0_E2END[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3002_ net1014 _1410_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q
+ VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__mux2_4
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4953_ net40 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_135_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3904_ net210 net1067 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__mux2_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4884_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 VGND VGND VPWR VPWR net235
+ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_22_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3835_ _0741_ _0745_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3766_ net1038 net740 net1032 net1021 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR
+ _0684_ sky130_fd_sc_hd__mux4_2
X_2717_ net62 net77 net113 net1053 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_144_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3697_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ net1062 _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__o21ai_4
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput320 net320 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput353 net353 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput342 net342 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
X_2648_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q _1598_ _1600_
+ _0141_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__o211a_1
XFILLER_160_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput375 net375 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[13] sky130_fd_sc_hd__buf_6
Xoutput386 net386 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[9] sky130_fd_sc_hd__buf_6
Xoutput364 net364 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_120_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2579_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 net105 net13 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__mux4_2
XFILLER_160_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4318_ net1223 net1076 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput397 net397 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4249_ net1251 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_153_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_162_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_171_Left_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1950_ _0951_ _0904_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__and2b_1
XFILLER_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_180_Left_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3620_ net174 net182 net120 net128 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR
+ _0549_ sky130_fd_sc_hd__mux4_1
X_3551_ net99 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q VGND
+ VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
X_2502_ _1345_ _1452_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__xnor2_2
X_3482_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0420_ _0421_
+ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__a21o_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5221_ net213 VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__buf_1
X_2433_ _1410_ _1411_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__mux2_1
XFILLER_102_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5152_ net154 VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__buf_1
X_2364_ net202 net128 net74 net218 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q VGND VGND VPWR VPWR
+ _1347_ sky130_fd_sc_hd__mux4_2
X_4103_ net48 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5083_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net425
+ sky130_fd_sc_hd__clkbuf_1
X_2295_ net978 net983 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__mux2_1
XFILLER_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4034_ net1227 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4936_ net51 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_2
XFILLER_20_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4867_ net1206 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_177_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3818_ _0679_ _0680_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4798_ net157 net1164 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_180_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3749_ net83 net91 net215 net229 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0669_ sky130_fd_sc_hd__mux4_1
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone123 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 VGND VGND VPWR VPWR
+ net740 sky130_fd_sc_hd__buf_6
XFILLER_93_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2080_ _0878_ _0981_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__nor2_4
XFILLER_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2982_ _1850_ _1849_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q
+ VGND VGND VPWR VPWR _1851_ sky130_fd_sc_hd__mux2_1
X_1933_ _0933_ _0935_ _0928_ _0120_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__a211o_1
X_4721_ net165 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4652_ net1181 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput30 Tile_X0Y0_FrameData[12] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3603_ net174 net182 net120 net128 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0534_ sky130_fd_sc_hd__mux4_1
Xinput63 Tile_X0Y0_S2END[2] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xinput41 Tile_X0Y0_FrameData[22] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
Xinput52 Tile_X0Y0_FrameData[5] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
X_4583_ net1211 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput85 Tile_X0Y0_SS4END[0] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xinput74 Tile_X0Y0_S2MID[5] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_4
XFILLER_155_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput96 Tile_X0Y0_W1END[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_1
X_3534_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q _0467_ VGND VGND
+ VPWR VPWR _0469_ sky130_fd_sc_hd__nand2_1
XFILLER_170_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3465_ _0405_ _0402_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 sky130_fd_sc_hd__mux2_4
XFILLER_115_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5204_ Tile_X0Y0_SS4END[11] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__buf_6
XFILLER_130_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2416_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q _1393_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q
+ _1395_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_149_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3396_ _0064_ _0341_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o21a_1
XFILLER_96_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2347_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q _1301_ VGND VGND
+ VPWR VPWR _1331_ sky130_fd_sc_hd__nand2_2
X_5135_ net165 VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__buf_1
X_5066_ Tile_X0Y0_W6END[11] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__buf_4
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2278_ _1260_ _1267_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5
+ sky130_fd_sc_hd__nand2_2
X_4017_ net1242 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4919_ Tile_X0Y0_EE4END[7] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_1
XFILLER_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3250_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q _0202_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q
+ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__a21o_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1150 net1151 VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__clkbuf_2
X_2201_ net974 net970 net989 net994 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ _1195_ sky130_fd_sc_hd__mux4_1
X_3181_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q VGND VGND VPWR
+ VPWR _0136_ sky130_fd_sc_hd__inv_1
Xfanout1161 net1162 VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__clkbuf_2
X_2132_ net690 net14 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q
+ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__mux2_2
Xfanout1183 net168 VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__buf_4
Xfanout1172 net1173 VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__buf_2
XFILLER_93_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1194 Tile_X0Y1_FrameData[27] VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__clkbuf_2
X_2063_ _1047_ _1048_ _1042_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_144_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4704_ net1203 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2965_ _0940_ _1329_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__mux2_1
XFILLER_147_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1916_ _0889_ _0911_ _0914_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_60_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2896_ _0818_ _1421_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__mux2_1
XFILLER_162_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4635_ net1197 net1106 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4566_ net1191 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3517_ _0451_ _0452_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q
+ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux2_4
XFILLER_143_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4497_ net1190 net1173 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3448_ net94 net1219 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
XFILLER_134_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3379_ _0042_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q VGND VGND
+ VPWR VPWR _0326_ sky130_fd_sc_hd__and2_1
XFILLER_69_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5118_ Tile_X0Y1_EE4END[5] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5049_ net105 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone99 net994 VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__buf_8
XFILLER_175_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput220 Tile_X0Y1_W2END[7] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput231 Tile_X0Y1_WW4END[0] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_2
XFILLER_48_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2750_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q net1055 VGND
+ VGND VPWR VPWR _1668_ sky130_fd_sc_hd__nor2_1
XFILLER_83_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2681_ _1623_ _1624_ _1625_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR VPWR
+ _1626_ sky130_fd_sc_hd__a221o_1
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4420_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs _0008_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4351_ net1224 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_152_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3302_ net200 net80 net23 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q VGND VGND VPWR VPWR
+ _0252_ sky130_fd_sc_hd__mux4_1
X_4282_ net29 net1083 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3233_ _0186_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q VGND VGND
+ VPWR VPWR _0187_ sky130_fd_sc_hd__or2_4
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3164_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q VGND VGND VPWR
+ VPWR _0119_ sky130_fd_sc_hd__inv_1
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3095_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR
+ VPWR _0050_ sky130_fd_sc_hd__inv_2
X_2115_ _1111_ _1114_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__xnor2_2
XFILLER_81_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2046_ _1045_ _1046_ _1043_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__a21o_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3997_ _0899_ _0900_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__and2_4
XFILLER_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2948_ net999 net1018 net693 net709 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q VGND VGND VPWR VPWR
+ _1822_ sky130_fd_sc_hd__mux4_1
XFILLER_129_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2879_ _0152_ _1764_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__o21a_1
X_4618_ net172 net1112 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4549_ net1209 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout965 _0299_ VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__buf_6
Xfanout976 net977 VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__buf_2
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout987 net988 VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__buf_2
Xfanout998 net999 VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__buf_2
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3920_ _0820_ _0826_ _0804_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B2 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_141_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3851_ _0748_ _0753_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__nor3b_2
X_2802_ _0704_ _1509_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q
+ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__mux2_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3782_ _0698_ _0697_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q
+ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__mux2_4
XFILLER_157_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2733_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q net1054 VGND
+ VGND VPWR VPWR _1655_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2664_ _1613_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 sky130_fd_sc_hd__mux2_4
XFILLER_117_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput502 net502 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[26] sky130_fd_sc_hd__buf_2
XFILLER_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4403_ net1245 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2595_ _0139_ _0274_ _1549_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__a21o_1
Xoutput524 net524 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[4] sky130_fd_sc_hd__buf_8
Xoutput535 net535 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput513 net513 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[7] sky130_fd_sc_hd__buf_2
X_4334_ net1239 net1170 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput568 net568 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput546 net546 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput557 net557 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_115_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput579 net579 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[7] sky130_fd_sc_hd__buf_2
X_4265_ net45 net1084 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4196_ net38 net1109 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3216_ _0166_ _0164_ _0169_ _0034_ _0032_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__a221o_1
XFILLER_94_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3147_ net135 VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_1
XFILLER_54_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3078_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR
+ VPWR _0033_ sky130_fd_sc_hd__inv_2
XFILLER_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2029_ _0740_ net625 VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__nor2_1
XFILLER_24_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2380_ _1360_ net1003 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__mux2_2
XFILLER_110_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4050_ net1244 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 Tile_X0Y0_E2END[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
X_3001_ _1349_ _0672_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q
+ VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__mux2_2
XFILLER_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4952_ net39 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__buf_1
XFILLER_101_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3903_ _0061_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__a21oi_1
X_4883_ net145 net1149 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_177_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3834_ _0741_ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__or2_4
XFILLER_32_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3765_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q _0682_ VGND VGND
+ VPWR VPWR _0683_ sky130_fd_sc_hd__nand2b_1
XFILLER_145_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2716_ net61 net114 net80 net1025 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_1
X_3696_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\] net1062 VGND VGND VPWR VPWR _0619_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_30_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2647_ _0140_ _1599_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__or2_1
Xoutput310 net310 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[5] sky130_fd_sc_hd__buf_2
XFILLER_145_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 net343 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput321 net321 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput332 net332 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
XFILLER_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput387 net387 VGND VGND VPWR VPWR Tile_X0Y0_UserCLKo sky130_fd_sc_hd__buf_1
Xoutput365 net365 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput354 net354 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput376 net376 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[14] sky130_fd_sc_hd__buf_2
X_2578_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q _1531_ _1535_
+ _1525_ _1527_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6
+ sky130_fd_sc_hd__o32a_2
X_4317_ net1222 net1076 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput398 net398 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[6] sky130_fd_sc_hd__buf_2
X_4248_ net1250 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4179_ net1245 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_182_Right_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3550_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q _0484_ VGND VGND
+ VPWR VPWR _0485_ sky130_fd_sc_hd__and2b_1
X_2501_ _1470_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\] net1065 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 sky130_fd_sc_hd__mux2_4
X_3481_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0419_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q
+ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__o21ai_1
X_5220_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net571
+ sky130_fd_sc_hd__buf_1
XFILLER_142_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2432_ net190 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net226
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q
+ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__mux4_2
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2363_ net140 net82 net234 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR
+ _1346_ sky130_fd_sc_hd__mux4_2
X_5151_ net1204 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__clkbuf_2
X_4102_ net1228 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5082_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR net424
+ sky130_fd_sc_hd__buf_4
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4033_ net1226 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2294_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q _1279_ _1277_
+ _1281_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q VGND VGND VPWR
+ VPWR _1282_ sky130_fd_sc_hd__a311o_1
XFILLER_56_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4935_ net50 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__buf_1
XFILLER_177_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4866_ net1205 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_177_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3817_ net665 _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__or2_1
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4797_ net158 net1166 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3748_ net203 net143 net119 net1216 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q VGND VGND VPWR VPWR
+ _0668_ sky130_fd_sc_hd__mux4_1
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3679_ net737 net736 net1030 net1023 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0604_ sky130_fd_sc_hd__mux4_1
XFILLER_101_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2981_ net709 _1410_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q
+ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__mux2_1
X_1932_ _0935_ _0933_ _0928_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4
+ sky130_fd_sc_hd__a21o_1
X_4720_ net166 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4651_ net171 net1105 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput31 Tile_X0Y0_FrameData[13] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput20 Tile_X0Y0_E2MID[7] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_99_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3602_ _0531_ _0530_ _0532_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ _0079_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__a221o_1
Xinput64 Tile_X0Y0_S2END[3] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
XFILLER_174_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput42 Tile_X0Y0_FrameData[23] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput53 Tile_X0Y0_FrameData[6] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
X_4582_ net1210 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput86 Tile_X0Y0_SS4END[1] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
Xinput75 Tile_X0Y0_S2MID[6] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_4
X_3533_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__inv_4
Xinput97 Tile_X0Y0_W2END[0] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3464_ _0403_ _0404_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q
+ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux2_4
XFILLER_115_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5203_ Tile_X0Y0_SS4END[10] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__buf_6
XFILLER_130_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2415_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q _1394_ VGND VGND
+ VPWR VPWR _1395_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_149_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3395_ net1036 net1006 net1031 net1021 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0341_ sky130_fd_sc_hd__mux4_1
XFILLER_130_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5134_ net155 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkbuf_1
XFILLER_96_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2346_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q _1329_ _1328_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR VPWR
+ _1330_ sky130_fd_sc_hd__o211a_1
X_5065_ Tile_X0Y0_W6END[10] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__buf_2
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2277_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q _1262_ _1264_
+ _1266_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q VGND VGND VPWR
+ VPWR _1267_ sky130_fd_sc_hd__a311o_1
X_4016_ net1241 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_108_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4918_ Tile_X0Y0_EE4END[6] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__buf_1
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4849_ net1190 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_165_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2200_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\]
+ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__and2_1
Xfanout1140 net1145 VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__clkbuf_2
X_3180_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q VGND VGND VPWR
+ VPWR _0135_ sky130_fd_sc_hd__inv_1
Xfanout1151 net1152 VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__clkbuf_2
X_2131_ _1129_ _1128_ _1130_ _0090_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__a221o_1
Xfanout1162 Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1173 net1174 VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2062_ _1062_ _1058_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__nor2_1
Xfanout1184 net167 VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__buf_4
Xfanout1195 net162 VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2964_ net996 _0767_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__mux2_1
XFILLER_147_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1915_ _0916_ _0917_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__xnor2_1
X_4703_ net1201 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2895_ net176 net1217 net1067 net716 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR
+ _1776_ sky130_fd_sc_hd__mux4_1
XFILLER_147_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4634_ net1196 net1106 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4565_ net1188 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3516_ net715 net995 net1016 net714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _0452_ sky130_fd_sc_hd__mux4_2
XFILLER_143_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4496_ net1185 net1173 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3447_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q _0388_ VGND VGND
+ VPWR VPWR _0389_ sky130_fd_sc_hd__or2_1
XFILLER_103_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3378_ _0218_ _0217_ _0242_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a211oi_2
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2329_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q _1312_ _1314_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR VPWR
+ _1315_ sky130_fd_sc_hd__o211a_1
XFILLER_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5117_ Tile_X0Y1_EE4END[4] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_1
XFILLER_182_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5048_ net104 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_68_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone45 net1059 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ _0728_ VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__o21ai_4
XFILLER_175_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone78 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 VGND VGND VPWR VPWR
+ net695 sky130_fd_sc_hd__buf_6
XFILLER_175_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput210 Tile_X0Y1_W1END[1] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_4
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput221 Tile_X0Y1_W2MID[0] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_4
Xinput232 Tile_X0Y1_WW4END[1] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ net6 net22 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q VGND
+ VGND VPWR VPWR _1625_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4350_ net1223 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3301_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q _0247_ _0251_
+ _0160_ _0162_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4
+ sky130_fd_sc_hd__o32a_2
XFILLER_152_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4281_ net1251 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3232_ net1009 net1024 net713 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0186_ sky130_fd_sc_hd__mux4_2
X_3163_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q VGND VGND VPWR
+ VPWR _0118_ sky130_fd_sc_hd__inv_1
XFILLER_39_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2114_ _1111_ _1114_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__or2_4
XFILLER_66_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3094_ net187 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2045_ net662 net625 _1000_ _1044_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_65_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3996_ _0766_ _0840_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__xor2_1
XFILLER_22_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2947_ _1820_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q VGND
+ VGND VPWR VPWR _1821_ sky130_fd_sc_hd__nand2b_1
XFILLER_175_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2878_ net981 net995 net1017 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _1764_ sky130_fd_sc_hd__mux4_1
X_4617_ net146 net1112 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4548_ net1208 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4479_ net1201 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout977 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 VGND VGND VPWR VPWR net977
+ sky130_fd_sc_hd__buf_8
Xfanout966 net731 VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__buf_8
XFILLER_38_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout988 net989 VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__buf_2
Xfanout999 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 VGND VGND VPWR VPWR net999
+ sky130_fd_sc_hd__buf_8
XFILLER_161_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3850_ _0761_ _0493_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__xnor2_2
X_2801_ net621 net59 net1220 net1028 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q VGND VGND VPWR VPWR
+ _1712_ sky130_fd_sc_hd__mux4_1
X_3781_ net972 net967 net990 net976 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0698_ sky130_fd_sc_hd__mux4_1
X_2732_ _1654_ _1653_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2663_ _1460_ _1612_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__xor2_1
XFILLER_8_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4402_ net1244 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2594_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR
+ _1549_ sky130_fd_sc_hd__a21bo_1
Xoutput503 net503 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput514 net514 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[8] sky130_fd_sc_hd__buf_2
Xoutput525 net525 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput536 net536 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[0] sky130_fd_sc_hd__buf_2
X_4333_ net1238 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput569 net569 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput547 net547 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput558 net558 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[15] sky130_fd_sc_hd__buf_2
X_4264_ net46 net1084 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3215_ _0164_ _0166_ _0169_ _0034_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2
+ sky130_fd_sc_hd__a22o_1
X_4195_ net1230 net1110 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3146_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q VGND VGND VPWR
+ VPWR _0101_ sky130_fd_sc_hd__inv_1
XFILLER_39_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3077_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q VGND VGND VPWR
+ VPWR _0032_ sky130_fd_sc_hd__inv_1
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2028_ _0998_ _1024_ _1027_ _1026_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__a22o_4
XFILLER_35_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3979_ _0786_ _0879_ _0881_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 Tile_X0Y0_E2END[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
X_3000_ net174 net210 _0529_ net983 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q VGND VGND VPWR VPWR
+ _1865_ sky130_fd_sc_hd__mux4_2
XFILLER_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4951_ net1244 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3902_ _0527_ _0528_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ _0522_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__a211o_1
X_4882_ net155 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3833_ _0621_ _0742_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__xnor2_2
XFILLER_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3764_ net1012 net1047 net1027 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR
+ _0682_ sky130_fd_sc_hd__mux4_1
X_2715_ net1256 net79 net64 net1048 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 sky130_fd_sc_hd__mux4_1
X_3695_ _0618_ _0616_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_30_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput300 net300 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[25] sky130_fd_sc_hd__buf_2
X_2646_ net1 net23 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q VGND
+ VGND VPWR VPWR _1599_ sky130_fd_sc_hd__mux2_1
Xoutput333 net333 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput322 net322 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput344 net344 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput311 net311 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[6] sky130_fd_sc_hd__buf_2
XFILLER_160_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput355 net355 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput377 net377 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[15] sky130_fd_sc_hd__buf_6
Xoutput366 net366 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[5] sky130_fd_sc_hd__buf_2
X_2577_ _0097_ _1534_ _1533_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q
+ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__o211a_1
XFILLER_113_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4316_ net1221 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput399 net399 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput388 net388 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_101_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4247_ net32 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4178_ net1244 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_161_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3129_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR
+ VPWR _0084_ sky130_fd_sc_hd__inv_2
XFILLER_15_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_85_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3480_ net997 net1014 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux2_1
X_2500_ _1451_ _1359_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__xor2_1
XFILLER_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2431_ net189 net225 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q
+ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__mux4_2
X_5150_ net1205 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__buf_1
X_2362_ _1343_ _1344_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__nand2b_4
XFILLER_150_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5081_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR net423
+ sky130_fd_sc_hd__clkbuf_2
X_4101_ net1254 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2293_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q _1280_ VGND VGND
+ VPWR VPWR _1281_ sky130_fd_sc_hd__nor2_1
XFILLER_110_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4032_ net1225 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_regs_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK VGND VGND VPWR VPWR Tile_X0Y1_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_35_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4934_ net47 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__buf_1
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4865_ net1204 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_177_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3816_ net1059 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ _0728_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__o21ai_4
X_4796_ net1198 net1164 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_165_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3747_ _0104_ _0664_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__o21a_1
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3678_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q _0602_ VGND VGND
+ VPWR VPWR _0603_ sky130_fd_sc_hd__or2_4
X_2629_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q _1582_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__a21bo_1
XFILLER_133_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2980_ _1349_ _0598_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q
+ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__mux2_1
X_1931_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _0934_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__o21ba_1
XFILLER_61_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4650_ net1179 net1105 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput21 Tile_X0Y0_E6END[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_147_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput10 Tile_X0Y0_E2END[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_99_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3601_ net210 net1067 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux2_1
XFILLER_174_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput43 Tile_X0Y0_FrameData[24] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xinput32 Tile_X0Y0_FrameData[14] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput54 Tile_X0Y0_FrameData[7] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
X_4581_ net1209 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput65 Tile_X0Y0_S2END[4] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xinput76 Tile_X0Y0_S2MID[7] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
Xinput87 Tile_X0Y0_SS4END[2] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
XFILLER_155_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3532_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q _0464_ _0466_
+ _0460_ _0462_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__o32a_4
Xinput98 Tile_X0Y0_W2END[1] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
XFILLER_170_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3463_ net1256 net65 net101 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0404_ sky130_fd_sc_hd__mux4_1
XFILLER_115_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5202_ Tile_X0Y0_SS4END[9] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__buf_6
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2414_ net131 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q
+ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__mux2_4
X_3394_ _0339_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q VGND VGND
+ VPWR VPWR _0340_ sky130_fd_sc_hd__or2_4
XFILLER_130_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5133_ net145 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__buf_1
X_2345_ net178 net144 net70 net214 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q VGND VGND VPWR VPWR
+ _1329_ sky130_fd_sc_hd__mux4_2
X_5064_ Tile_X0Y0_W6END[9] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_4
XFILLER_123_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2276_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q _1265_ VGND VGND
+ VPWR VPWR _1266_ sky130_fd_sc_hd__nor2_1
X_4015_ net1240 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_108_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4917_ Tile_X0Y0_EE4END[5] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__buf_1
X_4848_ net166 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4779_ net1180 net1070 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_180_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_168_Left_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1141 net1144 VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1130 net1131 VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2130_ net13 net69 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q VGND
+ VGND VPWR VPWR _1130_ sky130_fd_sc_hd__mux2_1
XFILLER_93_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1152 net1153 VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__buf_4
Xfanout1174 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__clkbuf_2
Xfanout1163 net1164 VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__buf_2
XFILLER_120_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2061_ _1043_ _1059_ _1061_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__a21o_1
Xfanout1196 net161 VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__clkbuf_4
Xfanout1185 net166 VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__buf_4
XFILLER_81_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_177_Left_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2963_ net175 net1218 net1068 net986 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q VGND VGND VPWR VPWR
+ _1835_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_103_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1914_ _0916_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__nand2_1
X_4702_ net1200 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2894_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q _1771_ _1773_
+ _1775_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A sky130_fd_sc_hd__o22a_1
XFILLER_8_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4633_ net1195 net1106 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4564_ net1186 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3515_ net691 net707 net991 net975 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _0451_ sky130_fd_sc_hd__mux4_2
XFILLER_170_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4495_ net1184 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3446_ net60 net68 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q VGND
+ VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux2_1
XFILLER_143_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3377_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q net1030 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q
+ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__o21ba_2
XFILLER_111_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2328_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q _1313_ VGND VGND
+ VPWR VPWR _1314_ sky130_fd_sc_hd__nand2_1
X_5116_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 VGND VGND VPWR VPWR net458
+ sky130_fd_sc_hd__buf_6
X_5047_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR net398
+ sky130_fd_sc_hd__buf_4
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2259_ _1249_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__inv_1
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_177_Right_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput200 Tile_X0Y1_N4END[7] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_4
Xinput211 Tile_X0Y1_W1END[2] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_2
XFILLER_102_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput222 Tile_X0Y1_W2MID[1] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_4
Xinput233 Tile_X0Y1_WW4END[2] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
XFILLER_124_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3300_ _0084_ _0250_ _0249_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q
+ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__o211a_1
XFILLER_165_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4280_ net1250 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_125_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3231_ _0183_ _0029_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__a21boi_4
XFILLER_140_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3162_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q VGND VGND VPWR
+ VPWR _0117_ sky130_fd_sc_hd__inv_2
X_2113_ _1113_ _1112_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__xnor2_2
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3093_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q VGND VGND VPWR
+ VPWR _0048_ sky130_fd_sc_hd__inv_1
XFILLER_54_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2044_ net662 _0981_ _1000_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3995_ _0898_ _0897_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__and2b_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2946_ _0767_ _0940_ _1429_ net1003 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q VGND VGND VPWR VPWR
+ _1820_ sky130_fd_sc_hd__mux4_1
X_2877_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q _1762_ VGND VGND
+ VPWR VPWR _1763_ sky130_fd_sc_hd__or2_1
XFILLER_175_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4616_ net147 net1112 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4547_ net1207 net1131 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4478_ net1200 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q _0368_ _0372_
+ _0364_ _0366_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1
+ sky130_fd_sc_hd__o32a_4
XFILLER_131_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout967 net732 VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_164_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout978 net979 VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__buf_2
Xfanout989 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 VGND VGND VPWR VPWR net989
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_57_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2800_ _1708_ _1710_ _1711_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 sky130_fd_sc_hd__o22a_1
X_3780_ net982 net747 net1018 net714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0697_ sky130_fd_sc_hd__mux4_2
XFILLER_157_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2731_ _0199_ net93 net1 net1043 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q VGND VGND VPWR VPWR
+ _1654_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_100_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4401_ net1242 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2662_ _1146_ _1145_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_152_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2593_ _1548_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 sky130_fd_sc_hd__mux2_4
Xoutput504 net504 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput515 net515 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[9] sky130_fd_sc_hd__buf_2
Xoutput526 net526 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_113_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4332_ net1237 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput548 net548 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput537 net537 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput559 net559 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[1] sky130_fd_sc_hd__buf_2
X_4263_ net1229 net1084 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3214_ _0167_ _0168_ _0033_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux2_1
X_4194_ net1227 net1110 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_105_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3145_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR
+ VPWR _0100_ sky130_fd_sc_hd__inv_1
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3076_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q VGND VGND VPWR
+ VPWR _0031_ sky130_fd_sc_hd__inv_2
XFILLER_54_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2027_ _0998_ _1024_ _1027_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3978_ _0786_ _0879_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_114_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2929_ _1801_ _1804_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 sky130_fd_sc_hd__mux2_2
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 Tile_X0Y0_E2END[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_162_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ net36 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_1
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3901_ _0116_ _0808_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q
+ _0807_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__o211a_1
X_4881_ net165 net1149 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_177_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3832_ _0679_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__nand2_1
XFILLER_177_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3763_ _0621_ _0678_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__and2_4
XFILLER_145_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2714_ net1255 net78 net63 net1010 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 sky130_fd_sc_hd__mux4_1
X_3694_ _0617_ _0407_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q
+ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput301 net301 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[26] sky130_fd_sc_hd__buf_2
X_2645_ _0199_ net185 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__mux2_1
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput323 net323 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput334 net334 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
XFILLER_160_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput312 net312 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[7] sky130_fd_sc_hd__buf_2
XFILLER_145_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput367 net367 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput356 net356 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput345 net345 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput378 net378 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[1] sky130_fd_sc_hd__buf_2
X_2576_ net68 net1219 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__mux2_1
X_4315_ net1253 net1076 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput389 net389 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[1] sky130_fd_sc_hd__buf_4
XFILLER_59_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4246_ net33 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4177_ net1242 net1108 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3128_ net19 VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__inv_1
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ net964 _1462_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__and2b_1
XFILLER_82_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_122_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_131_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2430_ _1408_ _0230_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__mux2_4
XFILLER_51_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2361_ _1325_ _1341_ _1342_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__nand3_4
X_5080_ Tile_X0Y0_WW4END[15] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_2
X_4100_ net1243 net1132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2292_ net176 net184 net1217 net130 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR VPWR
+ _1280_ sky130_fd_sc_hd__mux4_1
X_4031_ net1224 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4933_ net1243 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__buf_4
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4864_ net1203 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3815_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\] net1059 VGND VGND VPWR VPWR _0728_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4795_ net1197 net1164 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_177_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3746_ _0665_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q VGND VGND
+ VPWR VPWR _0666_ sky130_fd_sc_hd__or2_4
XFILLER_20_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3677_ net708 net1045 net723 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0602_ sky130_fd_sc_hd__mux4_2
X_2628_ net1043 net740 net1038 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q VGND VGND VPWR VPWR
+ _1582_ sky130_fd_sc_hd__mux4_1
X_2559_ _1118_ _1461_ _1117_ _1503_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__o211a_4
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4229_ net27 net1101 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone126 net977 VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_49_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1930_ net174 net182 net120 net128 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR
+ _0934_ sky130_fd_sc_hd__mux4_1
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput22 Tile_X0Y0_E6END[1] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
Xinput11 Tile_X0Y0_E2END[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_138_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3600_ _0061_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a21oi_1
X_4580_ net1208 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput44 Tile_X0Y0_FrameData[25] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput33 Tile_X0Y0_FrameData[15] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_2
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput55 Tile_X0Y0_FrameData[8] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
XFILLER_155_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3531_ _0082_ _0465_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_99_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput88 Tile_X0Y0_SS4END[3] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 Tile_X0Y0_S4END[0] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput66 Tile_X0Y0_S2END[5] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
XFILLER_155_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3462_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net197 net189 net9 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q VGND VGND VPWR VPWR
+ _0403_ sky130_fd_sc_hd__mux4_2
XFILLER_115_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput99 Tile_X0Y0_W2END[2] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
XFILLER_6_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5201_ Tile_X0Y0_SS4END[8] VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__buf_6
XFILLER_170_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3393_ net708 net1024 net723 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0339_ sky130_fd_sc_hd__mux4_2
XFILLER_130_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2413_ net221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q
+ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__mux2_1
XFILLER_69_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2344_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q _1326_ VGND VGND
+ VPWR VPWR _1328_ sky130_fd_sc_hd__nand2_1
XFILLER_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5063_ Tile_X0Y0_W6END[8] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_4
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2275_ net175 net1218 net183 net129 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q VGND VGND VPWR VPWR
+ _1265_ sky130_fd_sc_hd__mux4_1
X_4014_ net1239 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4916_ Tile_X0Y0_EE4END[4] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__buf_1
X_4847_ net167 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4778_ net1179 net1070 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_180_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3729_ _0533_ _0535_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ _0507_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__a211o_1
XFILLER_161_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1131 net1136 VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1120 net1127 VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__buf_2
Xfanout1142 net1143 VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__buf_2
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1153 Tile_X0Y1_FrameStrobe[12] VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__clkbuf_2
Xfanout1164 net1166 VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__buf_2
Xfanout1175 net1178 VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2060_ _0676_ _0944_ net625 _0601_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__o22a_1
Xfanout1186 net1187 VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__buf_4
Xfanout1197 net160 VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2962_ _1827_ _1829_ _1834_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1
+ sky130_fd_sc_hd__o21ai_1
XFILLER_34_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1913_ _0886_ _0891_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_17_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ net1199 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4632_ net1193 net1106 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2893_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q _1774_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q
+ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__a21bo_1
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4563_ net1214 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3514_ net1062 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ _0449_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__o21ai_4
X_4494_ net1183 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3445_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q _0384_ _0386_
+ _0092_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o211a_1
XFILLER_143_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3376_ _0320_ _0319_ _0321_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ _0074_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a221o_2
XFILLER_69_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2327_ net210 net1067 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__mux2_1
X_5115_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 VGND VGND VPWR VPWR net457
+ sky130_fd_sc_hd__buf_1
XFILLER_57_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5046_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 VGND VGND VPWR VPWR net397
+ sky130_fd_sc_hd__buf_4
X_2258_ _0410_ net69 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_68_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2189_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q _1184_ VGND VGND
+ VPWR VPWR _1185_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput201 Tile_X0Y1_NN4END[0] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_89_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput212 Tile_X0Y1_W1END[3] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
Xinput223 Tile_X0Y1_W2MID[2] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_2
Xinput234 Tile_X0Y1_WW4END[3] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3230_ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__inv_1
X_3161_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q VGND VGND VPWR
+ VPWR _0116_ sky130_fd_sc_hd__inv_2
X_2112_ _0851_ _1105_ _0854_ _1107_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__o31a_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3092_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR
+ VPWR _0047_ sky130_fd_sc_hd__inv_2
XFILLER_81_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2043_ _0878_ _0828_ _0827_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_105_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3994_ _0838_ _0839_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2945_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q _1817_ _1818_
+ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__a21o_1
XFILLER_175_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2876_ net729 net985 net716 net975 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _1762_ sky130_fd_sc_hd__mux4_1
X_4615_ net1211 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4546_ net152 net1131 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_145_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4477_ net1199 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3428_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q _0369_ _0371_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q VGND VGND VPWR VPWR
+ _0372_ sky130_fd_sc_hd__o211a_1
X_3359_ _0304_ _0303_ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a21o_1
Xfanout968 net969 VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_5_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout979 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 VGND VGND VPWR VPWR net979
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5029_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__buf_6
XFILLER_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2730_ _1651_ _1652_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q
+ VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2661_ _1611_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 sky130_fd_sc_hd__mux2_4
XFILLER_8_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4400_ net1241 net1150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_117_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2592_ _1547_ _1521_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__xnor2_2
Xoutput505 net505 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[29] sky130_fd_sc_hd__buf_2
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput527 net527 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[7] sky130_fd_sc_hd__buf_4
Xoutput516 net516 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_125_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4331_ net1236 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput549 net549 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput538 net538 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[11] sky130_fd_sc_hd__buf_2
X_4262_ net1228 net1085 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3213_ net174 net180 net196 net126 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0168_ sky130_fd_sc_hd__mux4_1
X_4193_ net51 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3144_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q VGND VGND VPWR
+ VPWR _0099_ sky130_fd_sc_hd__inv_2
X_3075_ net73 VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_1
XFILLER_27_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2026_ _0574_ _0575_ _0784_ _1025_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__a31o_1
XFILLER_35_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3977_ _0880_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__inv_2
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2928_ _1803_ _1802_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q
+ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__mux2_1
XFILLER_163_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2859_ net691 net985 net716 net743 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _1754_ sky130_fd_sc_hd__mux4_1
XFILLER_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4529_ net1190 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 Tile_X0Y0_E2END[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XFILLER_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3900_ net984 net998 net1020 net1001 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0808_ sky130_fd_sc_hd__mux4_1
X_4880_ net1185 net1149 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_17_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3831_ _0620_ _0729_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__nor2_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3762_ _0620_ _0676_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__nor2_1
XFILLER_32_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2713_ net1005 _0322_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 _0346_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 sky130_fd_sc_hd__mux4_1
X_3693_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 net105 net69 _0274_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q VGND VGND VPWR VPWR
+ _0617_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2644_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q _1596_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__a21bo_1
Xoutput324 net324 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput335 net335 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[0] sky130_fd_sc_hd__buf_2
X_2575_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q _1532_ VGND VGND
+ VPWR VPWR _1533_ sky130_fd_sc_hd__or2_1
Xoutput302 net302 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput313 net313 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[8] sky130_fd_sc_hd__buf_2
XFILLER_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput368 net368 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput357 net357 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput346 net346 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[7] sky130_fd_sc_hd__buf_2
X_4314_ net1252 net1075 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput379 net379 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4245_ net34 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4176_ net1241 net1109 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3127_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q VGND VGND VPWR
+ VPWR _0082_ sky130_fd_sc_hd__inv_2
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ net964 _1613_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__and2b_1
XFILLER_150_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2009_ _1009_ _1008_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_81_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2360_ _1325_ _1341_ _1342_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__a21oi_2
XFILLER_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2291_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1278_ VGND VGND
+ VPWR VPWR _1279_ sky130_fd_sc_hd__nand2_1
XFILLER_110_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4030_ net1223 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4932_ net1254 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__buf_4
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4863_ net1201 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3814_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q _0711_ _0727_
+ _0722_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ sky130_fd_sc_hd__a22o_4
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4794_ net1196 net1164 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_158_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3745_ net971 net985 net716 net976 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0665_ sky130_fd_sc_hd__mux4_2
XFILLER_20_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3676_ net1059 Tile_X0Y1_DSP_bot.A3 _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__o21ai_4
X_2627_ _0143_ _1580_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__and2_1
XFILLER_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2558_ _1506_ _1515_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__xnor2_2
XFILLER_87_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2489_ _1447_ _1463_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__and2_4
X_4228_ net38 net1101 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4159_ net53 net1118 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone105 net1060 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ _0542_ VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__o21ai_4
Xclone127 net745 net725 _0197_ _0198_ VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__a22o_4
Xclone116 net734 VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 Tile_X0Y0_E2END[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput45 Tile_X0Y0_FrameData[28] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xinput34 Tile_X0Y0_FrameData[16] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
Xinput23 Tile_X0Y0_EE4END[0] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
X_3530_ net65 net101 net77 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q VGND VGND VPWR VPWR
+ _0465_ sky130_fd_sc_hd__mux4_1
Xinput89 Tile_X0Y0_SS4END[4] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_4
Xinput78 Tile_X0Y0_S4END[1] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
Xinput67 Tile_X0Y0_S2END[6] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput56 Tile_X0Y0_FrameData[9] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XFILLER_155_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3461_ _0400_ _0401_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q
+ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux2_4
XFILLER_115_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3392_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q _0329_ _0334_
+ _0338_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 sky130_fd_sc_hd__o31ai_2
X_5200_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net542
+ sky130_fd_sc_hd__buf_1
X_2412_ _1391_ _1390_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__mux2_1
XFILLER_170_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2343_ _1326_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__inv_2
X_5131_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 VGND VGND VPWR VPWR net473
+ sky130_fd_sc_hd__buf_6
X_5062_ Tile_X0Y0_W6END[7] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_2
X_4013_ net1238 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2274_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q _1263_ VGND VGND
+ VPWR VPWR _1264_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4915_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 VGND VGND VPWR VPWR net257
+ sky130_fd_sc_hd__clkbuf_2
X_4846_ net168 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1989_ _0966_ _0982_ _0985_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4777_ net1213 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_180_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3728_ net73 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux2_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3659_ net186 net132 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__mux2_1
XFILLER_164_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1132 net1133 VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1121 net1122 VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__buf_2
XFILLER_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1110 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__clkbuf_4
Xfanout1143 net1144 VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1154 net1155 VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__clkbuf_2
Xfanout1165 net1166 VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__clkbuf_2
Xfanout1176 net1177 VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1198 net159 VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__buf_4
Xfanout1187 Tile_X0Y1_FrameData[31] VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2961_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q _1833_ _1831_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q VGND VGND VPWR VPWR
+ _1834_ sky130_fd_sc_hd__a211o_1
XFILLER_34_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1912_ _0909_ _0915_ _0908_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__a21o_1
X_4700_ net1198 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4631_ net1192 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2892_ _0940_ _1364_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__mux2_1
XFILLER_128_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs VGND VGND VPWR
+ VPWR clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4562_ net1202 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3513_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\] net1062 VGND VGND VPWR VPWR _0449_
+ sky130_fd_sc_hd__nand2b_1
X_4493_ net1182 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3444_ _0091_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__or2_1
XFILLER_170_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3375_ _0319_ _0320_ _0321_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__a22o_1
XFILLER_111_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2326_ _0349_ _0045_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__mux2_1
XFILLER_69_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5114_ Tile_X0Y1_E6END[11] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__buf_1
X_5045_ net101 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_1
XFILLER_111_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2257_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q _1245_ _1247_
+ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__o21ai_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2188_ _1182_ _1183_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q
+ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__mux2_1
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone59 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 VGND VGND VPWR VPWR
+ net676 sky130_fd_sc_hd__buf_8
Xclone48 net1061 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ _0708_ VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__o21ai_4
X_4829_ net158 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput202 Tile_X0Y1_NN4END[1] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput224 Tile_X0Y1_W2MID[3] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_2
Xinput213 Tile_X0Y1_W2END[0] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3160_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q VGND VGND VPWR
+ VPWR _0115_ sky130_fd_sc_hd__inv_2
X_2111_ _0843_ _1103_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__nor2_1
XFILLER_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3091_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR
+ VPWR _0046_ sky130_fd_sc_hd__inv_1
XFILLER_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2042_ _0601_ _0944_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__nor2_1
XFILLER_54_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3993_ _0895_ _0896_ _0894_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__a21bo_1
XFILLER_22_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2944_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q _1816_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2875_ net715 _0196_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 _0173_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_175_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4614_ net1210 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_175_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4545_ net153 net1131 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4476_ net1198 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3427_ _0370_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q VGND VGND
+ VPWR VPWR _0371_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3358_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q _0305_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q
+ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a21bo_1
XFILLER_161_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout969 net970 VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__buf_6
X_2309_ net76 net1067 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__mux2_1
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3289_ _0239_ _0233_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_2
X_5028_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_6
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2660_ _1563_ _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_100_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2591_ _1546_ _1544_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__nor2_4
XFILLER_125_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput506 net506 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput517 net517 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[1] sky130_fd_sc_hd__buf_2
X_4330_ net1233 net1169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput528 net528 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput539 net539 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[12] sky130_fd_sc_hd__buf_2
XFILLER_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4261_ net1254 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3212_ net140 net72 net216 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0167_ sky130_fd_sc_hd__mux4_1
X_4192_ net1225 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_79_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3143_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q VGND VGND VPWR
+ VPWR _0098_ sky130_fd_sc_hd__inv_2
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3074_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q VGND VGND VPWR
+ VPWR _0029_ sky130_fd_sc_hd__inv_2
X_2025_ _0827_ _0677_ _0828_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__and3_1
XFILLER_47_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3976_ _0676_ _0709_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__nor2_1
X_2927_ net1000 _1429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__mux2_1
XFILLER_40_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2858_ net980 net995 net1016 net709 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _1753_ sky130_fd_sc_hd__mux4_1
XFILLER_163_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2789_ _1701_ _1702_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_170_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4528_ net1185 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4459_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3830_ net662 _0661_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__nor2_4
XFILLER_32_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3761_ _0601_ _0661_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__nor2_1
X_2712_ net1035 net965 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 _0278_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_145_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3692_ _0615_ _0614_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q
+ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_30_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2643_ net1042 net1007 net1037 net1021 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q VGND VGND VPWR VPWR
+ _1596_ sky130_fd_sc_hd__mux4_1
Xoutput325 net325 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
X_2574_ net58 net60 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q VGND
+ VGND VPWR VPWR _1532_ sky130_fd_sc_hd__mux2_1
Xoutput303 net303 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput314 net314 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[9] sky130_fd_sc_hd__buf_2
XFILLER_160_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput369 net369 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput358 net358 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput347 net347 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput336 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 VGND VGND VPWR VPWR
+ Tile_X0Y0_N1BEG[1] sky130_fd_sc_hd__buf_8
XFILLER_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4313_ net1251 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4244_ net35 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4175_ net1240 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3126_ net109 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__inv_1
XFILLER_67_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3057_ net964 _1478_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__and2b_1
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2008_ net625 net722 VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_81_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3959_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q _0864_ VGND VGND
+ VPWR VPWR _0865_ sky130_fd_sc_hd__and2_1
XFILLER_167_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2290_ net76 net1067 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_63_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4931_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 VGND VGND VPWR VPWR net273
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_177_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4862_ net1200 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3813_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q _0726_ VGND VGND
+ VPWR VPWR _0727_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_72_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4793_ net1195 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3744_ net692 net747 net733 net1013 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0664_ sky130_fd_sc_hd__mux4_1
X_3675_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\] net1059 VGND VGND VPWR VPWR _0600_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2626_ net1012 net1047 net1027 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR VPWR
+ _1580_ sky130_fd_sc_hd__mux4_1
X_2557_ _1506_ _1515_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_81_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2488_ _1416_ _1446_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__nand2_1
X_4227_ net47 net1100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4158_ net54 net1116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4089_ net30 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3109_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q VGND VGND VPWR
+ VPWR _0064_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_90_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone106 net1053 VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__buf_6
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone117 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 VGND VGND VPWR VPWR net734
+ sky130_fd_sc_hd__buf_6
XFILLER_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 Tile_X0Y0_E2MID[0] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XFILLER_52_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput46 Tile_X0Y0_FrameData[29] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput35 Tile_X0Y0_FrameData[17] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput24 Tile_X0Y0_EE4END[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput79 Tile_X0Y0_S4END[2] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
Xinput68 Tile_X0Y0_S2END[7] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
Xinput57 Tile_X0Y0_S1END[0] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_8
XFILLER_155_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3460_ net1034 net1005 net1029 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0401_ sky130_fd_sc_hd__mux4_1
XFILLER_115_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3391_ _0043_ _0335_ _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o21ai_2
X_2411_ net203 net124 net70 net214 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q VGND VGND VPWR VPWR
+ _1391_ sky130_fd_sc_hd__mux4_2
X_5130_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 VGND VGND VPWR VPWR net472
+ sky130_fd_sc_hd__buf_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2342_ _0112_ _0111_ _0021_ _0557_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q VGND VGND VPWR VPWR
+ _1326_ sky130_fd_sc_hd__mux4_2
X_5061_ Tile_X0Y0_W6END[6] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_2
XFILLER_96_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4012_ net44 net1178 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2273_ net209 net1068 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__mux2_1
XFILLER_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4914_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 VGND VGND VPWR VPWR net256
+ sky130_fd_sc_hd__clkbuf_1
X_4845_ net169 net1156 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4776_ net1212 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_165_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3727_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q _0648_ _0644_
+ _0638_ _0640_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4
+ sky130_fd_sc_hd__o32a_4
XFILLER_146_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1988_ _0987_ _0988_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__and2_1
XFILLER_180_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3658_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net222 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__mux2_1
XFILLER_164_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3589_ net198 net86 net101 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q VGND VGND VPWR VPWR
+ _0520_ sky130_fd_sc_hd__mux4_2
X_2609_ _1546_ _1560_ _1561_ _1559_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__o31a_1
XFILLER_161_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5259_ Tile_X0Y1_WW4END[14] VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__clkbuf_2
XFILLER_180_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_119_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1100 net1101 VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1122 net1127 VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__clkbuf_2
Xfanout1111 net1112 VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1133 net1136 VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__clkbuf_2
Xfanout1144 net1145 VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__buf_2
XFILLER_93_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1155 net1156 VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__buf_2
Xfanout1177 net1178 VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_137_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1166 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__buf_2
Xfanout1199 net158 VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__buf_4
Xfanout1188 net1189 VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__buf_4
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2960_ _1832_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__inv_1
X_1911_ _0910_ _0913_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2891_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q _1772_ VGND
+ VGND VPWR VPWR _1773_ sky130_fd_sc_hd__and2b_1
XFILLER_147_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ net1191 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4561_ net1190 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_155_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3512_ _0448_ _0442_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ sky130_fd_sc_hd__mux2_2
X_4492_ net1181 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3443_ net1257 net12 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__mux2_1
XFILLER_170_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ net74 net110 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q VGND
+ VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
XFILLER_69_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5113_ Tile_X0Y1_E6END[10] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__buf_1
X_2325_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q _1308_ _1310_
+ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__o21ai_1
X_5044_ net100 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__buf_1
XFILLER_111_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2256_ _0130_ _1246_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q
+ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__o21a_1
XFILLER_84_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2187_ net59 net67 net93 net1220 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q VGND VGND VPWR VPWR
+ _1183_ sky130_fd_sc_hd__mux4_1
XFILLER_65_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4828_ net159 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_181_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4759_ net1192 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput203 Tile_X0Y1_NN4END[2] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput225 Tile_X0Y1_W2MID[4] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_2
Xinput214 Tile_X0Y1_W2END[1] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_2
XFILLER_102_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2110_ _0857_ _1109_ _1110_ _1100_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__a22oi_4
X_3090_ net76 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__inv_2
XFILLER_66_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2041_ _1026_ _1028_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__xnor2_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3992_ _0892_ _0893_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2943_ net976 net692 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2874_ net70 net81 net229 net990 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_175_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4613_ net1209 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4544_ net154 net1131 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4475_ net1197 net1174 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3426_ net215 net229 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux2_1
X_3357_ net209 net1068 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2308_ _0349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q _1294_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR
+ _1295_ sky130_fd_sc_hd__a211o_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5027_ Tile_X0Y1_NN4END[15] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__buf_1
X_3288_ _0041_ _0238_ _0237_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a21o_1
XFILLER_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2239_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q _1230_ VGND VGND
+ VPWR VPWR _1231_ sky130_fd_sc_hd__or2_1
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2590_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q _1481_ _1543_
+ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__a21oi_1
Xoutput507 net507 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[30] sky130_fd_sc_hd__buf_2
XFILLER_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput518 net518 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_125_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput529 net529 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[1] sky130_fd_sc_hd__buf_2
XFILLER_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4260_ net1243 net1093 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4191_ net53 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3211_ _0165_ _0033_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__o21a_1
X_3142_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR
+ VPWR _0097_ sky130_fd_sc_hd__inv_2
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3073_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q VGND VGND VPWR
+ VPWR _0028_ sky130_fd_sc_hd__inv_2
X_2024_ _0450_ net624 VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__nor2_1
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3975_ _0620_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__nor2_1
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2926_ net1003 _0968_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__mux2_1
X_2857_ net743 _0196_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 _0173_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2788_ net1030 net721 _0652_ _1139_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q VGND VGND VPWR VPWR
+ _1702_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_170_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4527_ net167 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4458_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3409_ _0351_ _0352_ _0353_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ _0075_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__a221o_1
X_4389_ net1254 net1161 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_101_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_110_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3760_ _0659_ _0660_ _0677_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__and3_1
XFILLER_32_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2711_ net1042 _0526_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 _0520_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3691_ net185 net61 net24 net97 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q VGND VGND VPWR VPWR
+ _0615_ sky130_fd_sc_hd__mux4_1
X_2642_ _0141_ _1594_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__and2_1
Xoutput326 net326 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput315 net315 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
X_2573_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q _1528_ _1530_
+ _0098_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__o211a_1
Xoutput304 net304 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput348 net348 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput337 net337 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput359 net359 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[13] sky130_fd_sc_hd__buf_2
XFILLER_160_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4312_ net1250 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_99_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4243_ net36 net1091 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4174_ net1239 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3125_ net17 VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_1
X_3056_ net964 _1476_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__nor2_1
X_2007_ _0601_ _0829_ _0999_ _1001_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__o31ai_4
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3958_ net1043 net1032 net1038 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q VGND VGND VPWR VPWR
+ _0864_ sky130_fd_sc_hd__mux4_1
XFILLER_167_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3889_ net204 net120 net126 net1215 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0798_ sky130_fd_sc_hd__mux4_1
X_2909_ _1787_ VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__inv_1
XFILLER_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4930_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 VGND VGND VPWR VPWR net272
+ sky130_fd_sc_hd__buf_1
X_4861_ net1199 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_177_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3812_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q _0723_ _0725_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q VGND VGND VPWR VPWR
+ _0726_ sky130_fd_sc_hd__o211a_1
XFILLER_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4792_ net1193 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_158_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3743_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q _0382_ VGND VGND
+ VPWR VPWR _0663_ sky130_fd_sc_hd__nand2_1
XFILLER_173_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3674_ _0589_ _0599_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A3 sky130_fd_sc_hd__mux2_2
XFILLER_173_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2625_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q _1564_ _1578_
+ _1577_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q VGND VGND VPWR
+ VPWR _1579_ sky130_fd_sc_hd__o221a_1
XFILLER_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2556_ net1058 _1514_ _1507_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__a21oi_4
X_2487_ _1462_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 sky130_fd_sc_hd__mux2_4
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4226_ net50 net1100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4157_ net1222 net1116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3108_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR
+ VPWR _0063_ sky130_fd_sc_hd__inv_1
XFILLER_95_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4088_ net31 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_102_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3039_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q net703 VGND VGND
+ VPWR VPWR _1901_ sky130_fd_sc_hd__nand2_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone107 net1048 VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__buf_6
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput36 Tile_X0Y0_FrameData[18] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
Xinput25 Tile_X0Y0_EE4END[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
Xinput14 Tile_X0Y0_E2MID[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
Xinput69 Tile_X0Y0_S2MID[0] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_8
Xinput58 Tile_X0Y0_S1END[1] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xinput47 Tile_X0Y0_FrameData[2] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
XFILLER_155_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2410_ net144 net232 net81 _0184_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q VGND VGND VPWR VPWR
+ _1390_ sky130_fd_sc_hd__mux4_1
X_3390_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q _0336_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o21a_1
XFILLER_170_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2341_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\]
+ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__nand2_1
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5060_ Tile_X0Y0_W6END[5] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkbuf_2
X_2272_ _0059_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q
+ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__a211o_1
X_4011_ net1236 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4913_ Tile_X0Y0_E6END[11] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
XFILLER_60_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4844_ net170 net1156 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1987_ _0919_ _0947_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__xor2_1
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4775_ net1211 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_158_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3726_ _0087_ _0647_ _0646_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q
+ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__o211a_1
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3657_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q _0583_ VGND VGND
+ VPWR VPWR _0584_ sky130_fd_sc_hd__and2b_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2608_ _1546_ _1561_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__nor2_1
X_3588_ _0515_ _0078_ _0519_ _0511_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0
+ sky130_fd_sc_hd__a31o_4
X_2539_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[15\] net1064 VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__mux2_4
XFILLER_121_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5258_ Tile_X0Y1_WW4END[13] VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__clkbuf_2
X_5189_ Tile_X0Y0_S4END[12] VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__buf_6
X_4209_ net1242 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1101 net1102 VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__buf_2
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1112 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__clkbuf_2
Xfanout1134 net1136 VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__buf_2
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1123 net1124 VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__buf_2
XFILLER_78_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1145 Tile_X0Y1_FrameStrobe[1] VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__buf_2
Xfanout1156 net1157 VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__clkbuf_4
Xfanout1167 net1170 VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1178 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__buf_2
Xfanout1189 Tile_X0Y1_FrameData[30] VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1910_ _0740_ _0829_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__or3_1
X_2890_ net997 _0767_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__mux2_1
XFILLER_179_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4560_ net1185 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3511_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q _0447_ _0446_
+ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__o21ba_1
X_4491_ net1180 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3442_ net618 net192 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__mux2_4
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _0060_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2324_ _0134_ _1309_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q
+ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__o21a_1
X_5112_ Tile_X0Y1_E6END[9] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__buf_1
XFILLER_111_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5043_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 VGND VGND VPWR VPWR net394
+ sky130_fd_sc_hd__buf_1
XFILLER_84_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2255_ net978 net997 net983 net1014 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q VGND VGND VPWR VPWR
+ _1246_ sky130_fd_sc_hd__mux4_1
X_2186_ net619 net3 net191 net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR VPWR
+ _1182_ sky130_fd_sc_hd__mux4_1
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4827_ net1197 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4758_ net1191 net1069 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_175_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3709_ _0625_ _0623_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__o21ai_4
X_4689_ net1190 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_161_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput204 Tile_X0Y1_NN4END[3] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
Xinput226 Tile_X0Y1_W2MID[5] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_2
Xinput215 Tile_X0Y1_W2END[2] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_2
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2040_ _1022_ _1032_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__xor2_2
XFILLER_47_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3991_ _0832_ _0888_ _0890_ _0887_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2942_ _1815_ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__inv_1
XFILLER_175_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2873_ net69 net84 net230 net986 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4612_ net1208 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4543_ net1201 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_128_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4474_ net1196 net1174 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3425_ net1216 net71 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux2_1
XFILLER_97_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3356_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q _0059_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__a21oi_1
XFILLER_97_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2307_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q _0529_ VGND VGND
+ VPWR VPWR _1294_ sky130_fd_sc_hd__nor2_1
X_3287_ net176 net178 net124 net1215 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _0238_ sky130_fd_sc_hd__mux4_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5026_ Tile_X0Y1_NN4END[14] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__buf_1
X_2238_ net973 net968 net987 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR
+ _1230_ sky130_fd_sc_hd__mux4_1
XFILLER_72_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2169_ net188 net8 net64 net116 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q VGND VGND VPWR VPWR
+ _1166_ sky130_fd_sc_hd__mux4_2
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_156_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_165_Left_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_174_Left_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput508 net508 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[31] sky130_fd_sc_hd__buf_2
XFILLER_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput519 net519 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_140_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4190_ net54 net1107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_111_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3210_ net981 net730 net1017 net1013 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0165_ sky130_fd_sc_hd__mux4_2
X_3141_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR
+ VPWR _0096_ sky130_fd_sc_hd__inv_2
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3072_ net222 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__inv_1
X_2023_ net624 _0575_ _0574_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__and3b_1
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3974_ Tile_X0Y1_DSP_bot.A0 net1059 _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__o21ai_4
XFILLER_50_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2925_ net173 net119 _0410_ net979 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q VGND VGND VPWR VPWR
+ _1801_ sky130_fd_sc_hd__mux4_2
XFILLER_50_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2856_ net747 _0382_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net688
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_163_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2787_ net618 net96 net1257 net1049 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q VGND VGND VPWR VPWR
+ _1701_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_170_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4526_ net1183 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4457_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C9 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3408_ net210 net1067 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__mux2_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4388_ net1243 net1161 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3339_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q _0288_ VGND VGND
+ VPWR VPWR _0289_ sky130_fd_sc_hd__or2_1
XFILLER_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_181_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ Tile_X0Y1_N4END[13] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_1
XFILLER_171_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2710_ _1642_ _1643_ _1646_ _0069_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3690_ net197 net113 net85 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q VGND VGND VPWR VPWR
+ _0614_ sky130_fd_sc_hd__mux4_2
X_2641_ net1011 net1047 net1026 net1052 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR VPWR
+ _1594_ sky130_fd_sc_hd__mux4_1
Xoutput316 net316 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
X_2572_ _0097_ _1529_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__or2_1
Xoutput305 net305 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[2] sky130_fd_sc_hd__buf_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput327 net327 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput349 net349 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput338 net338 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_113_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4311_ net1249 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4242_ net37 net1091 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4173_ net1238 net1109 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3124_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q VGND VGND VPWR
+ VPWR _0079_ sky130_fd_sc_hd__inv_2
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3055_ net964 _1475_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__and2b_1
XFILLER_67_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2006_ _0740_ net626 VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__or2_1
XFILLER_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3957_ net1012 net1047 net1028 net1052 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR VPWR
+ _0863_ sky130_fd_sc_hd__mux4_1
XFILLER_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2908_ net1014 _1410_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q
+ VGND VGND VPWR VPWR _1787_ sky130_fd_sc_hd__mux2_1
X_3888_ _0796_ _0118_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__o21a_1
XFILLER_176_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2839_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q _1744_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q
+ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__a21bo_1
XFILLER_136_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4509_ net1199 net1139 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4860_ net1198 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3811_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q _0724_ VGND VGND
+ VPWR VPWR _0725_ sky130_fd_sc_hd__nand2_1
XFILLER_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4791_ net1192 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3742_ _0023_ _0102_ _0103_ _0229_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q VGND VGND VPWR VPWR
+ _0662_ sky130_fd_sc_hd__mux4_2
XFILLER_173_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3673_ _0598_ _0597_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q
+ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__mux2_1
XFILLER_173_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2624_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q _1127_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q
+ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__o21ai_1
XFILLER_141_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2555_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[16\] net1064 VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_117_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2486_ _1118_ _1461_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__xor2_1
XFILLER_87_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4225_ net1226 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4156_ net56 net1116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3107_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR
+ VPWR _0062_ sky130_fd_sc_hd__inv_2
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4087_ net1249 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_102_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3038_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ _0183_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR
+ VPWR _1900_ sky130_fd_sc_hd__o31a_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4989_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 VGND VGND VPWR VPWR net340
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone119 net1005 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__clkbuf_1
XFILLER_100_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput37 Tile_X0Y0_FrameData[19] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
Xinput26 Tile_X0Y0_EE4END[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
Xinput15 Tile_X0Y0_E2MID[2] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput59 Tile_X0Y0_S1END[2] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_6
Xinput48 Tile_X0Y0_FrameData[30] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
XFILLER_155_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2340_ _1321_ _1323_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_149_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2271_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q _0302_ VGND VGND
+ VPWR VPWR _1261_ sky130_fd_sc_hd__nor2_1
X_4010_ net1234 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4912_ Tile_X0Y0_E6END[10] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4843_ net171 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1986_ _0965_ _0986_ _0964_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__a21o_1
XFILLER_20_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4774_ net1210 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_165_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3725_ net94 net1219 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3656_ net185 net131 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q
+ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__mux2_1
XFILLER_161_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2607_ _1502_ _1517_ _1518_ _1545_ _1516_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__o311a_1
X_3587_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q _0518_ _0517_
+ _0077_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__a211o_1
XFILLER_161_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2538_ _1496_ _1499_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ sky130_fd_sc_hd__mux2_4
XFILLER_114_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5257_ Tile_X0Y1_WW4END[12] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__clkbuf_2
XFILLER_180_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4208_ net1241 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2469_ _1444_ _0981_ _0878_ _1442_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__nor4b_4
XFILLER_57_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5188_ Tile_X0Y0_S4END[11] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__buf_6
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4139_ net1235 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1102 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__clkbuf_2
Xfanout1113 net1114 VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__clkbuf_2
Xfanout1135 net1136 VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1124 net1127 VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__clkbuf_2
Xfanout1146 net1153 VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1168 net1170 VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1157 Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__clkbuf_2
Xfanout1179 net172 VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__buf_4
XFILLER_19_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3510_ net19 net111 net75 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q VGND VGND VPWR VPWR
+ _0447_ sky130_fd_sc_hd__mux4_1
XFILLER_128_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4490_ net172 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_170_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3441_ net980 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 _0382_ net688
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q
+ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__mux4_2
XFILLER_170_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3372_ net712 _0309_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q
+ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__a211o_1
XFILLER_170_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2323_ net978 net1019 net983 net1002 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q VGND VGND VPWR VPWR
+ _1309_ sky130_fd_sc_hd__mux4_1
X_5111_ Tile_X0Y1_E6END[8] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__buf_1
XFILLER_111_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5042_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR net393
+ sky130_fd_sc_hd__clkbuf_1
X_2254_ net974 net969 net988 net993 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q VGND VGND VPWR VPWR
+ _1245_ sky130_fd_sc_hd__mux4_1
X_2185_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q _1180_ VGND VGND
+ VPWR VPWR _1181_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_69_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4826_ net161 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1969_ net227 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q
+ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__o21a_1
X_4757_ net1189 net1072 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_175_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3708_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q _0626_ _0628_
+ _0630_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q VGND VGND VPWR
+ VPWR _0631_ sky130_fd_sc_hd__a221o_1
X_4688_ net1185 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3639_ net185 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q
+ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__mux2_1
XFILLER_161_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput205 Tile_X0Y1_NN4END[4] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_2
XFILLER_0_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput227 Tile_X0Y1_W2MID[6] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_2
Xinput216 Tile_X0Y1_W2END[3] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_87_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3990_ _0892_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_73_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2941_ net986 net990 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__mux2_1
XFILLER_90_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4611_ net1207 net1114 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2872_ net1216 net72 net83 net967 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_175_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4542_ net1200 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4473_ net1195 net1174 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3424_ _0022_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__and2_1
XFILLER_143_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3355_ _0279_ _0292_ _0055_ _0301_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__o211ai_2
XFILLER_97_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2306_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q _1290_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__o21ai_1
X_3286_ _0234_ _0235_ _0236_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR VPWR
+ _0237_ sky130_fd_sc_hd__o221a_1
X_5025_ Tile_X0Y1_NN4END[13] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_1
X_2237_ _0131_ _1228_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__or2_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2168_ _1160_ _1162_ _1165_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 sky130_fd_sc_hd__o22a_4
XFILLER_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2099_ _1097_ _1098_ _0859_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__a21o_4
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4809_ net146 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput509 net509 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[3] sky130_fd_sc_hd__buf_2
XFILLER_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3140_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR
+ VPWR _0095_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3071_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q VGND VGND VPWR
+ VPWR _0026_ sky130_fd_sc_hd__inv_2
XFILLER_82_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2022_ _0729_ net626 VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__or2_4
XFILLER_35_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3973_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\] net1059 VGND VGND VPWR VPWR _0877_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2924_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q _1794_ _1796_
+ _1800_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1
+ sky130_fd_sc_hd__a31oi_1
X_2855_ net692 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 net1003 _1327_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_163_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2786_ _1697_ _1700_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 sky130_fd_sc_hd__mux2_2
X_4525_ net169 net1145 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_170_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4456_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C8 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[8\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4387_ net1230 net1161 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3407_ _0045_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__a21oi_1
X_3338_ net1256 net63 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_1
XFILLER_105_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3269_ net715 net995 net1016 net1013 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ _0221_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_181_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5008_ Tile_X0Y1_N4END[12] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
XFILLER_85_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2640_ _0144_ _1592_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__or2_1
XFILLER_145_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput317 net317 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput306 net306 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[30] sky130_fd_sc_hd__buf_2
X_2571_ net1257 net12 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__mux2_1
Xoutput328 net328 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput339 net339 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_160_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4310_ net1248 net1076 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4241_ net1242 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4172_ net1237 net1109 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3123_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR
+ VPWR _0078_ sky130_fd_sc_hd__inv_1
X_3054_ net963 _1473_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__and2b_1
X_2005_ _0996_ _1004_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__xor2_4
XFILLER_23_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3956_ net192 net138 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 net228
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q
+ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__mux4_2
XFILLER_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2907_ _1349_ _0781_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q
+ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__mux2_1
XFILLER_176_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3887_ net982 net996 net1018 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0796_ sky130_fd_sc_hd__mux4_2
X_2838_ _1150_ _1512_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__mux2_1
X_2769_ _0148_ _1680_ _1685_ _1676_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0
+ sky130_fd_sc_hd__a31o_1
XFILLER_151_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4508_ net1198 net1139 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4439_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer71 _0373_ VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__buf_6
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer93 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 VGND VGND VPWR VPWR
+ net710 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3810_ net76 net112 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q VGND
+ VGND VPWR VPWR _0724_ sky130_fd_sc_hd__mux2_1
XFILLER_82_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4790_ net1191 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3741_ _0659_ _0660_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__nand2_8
XFILLER_20_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3672_ net177 net69 net123 net234 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q VGND VGND VPWR VPWR
+ _0598_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_41_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2623_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q _1572_ _1568_
+ _1576_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q VGND VGND VPWR
+ VPWR _1577_ sky130_fd_sc_hd__o311a_1
XFILLER_173_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2554_ _1513_ _1510_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ sky130_fd_sc_hd__mux2_4
XFILLER_126_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2485_ _1460_ _1144_ _1146_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__a21oi_4
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4224_ net1225 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4155_ net1253 net1116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_50_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3106_ net74 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__inv_2
XFILLER_55_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4086_ net1248 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3037_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q VGND VGND VPWR VPWR
+ _1899_ sky130_fd_sc_hd__o21ai_1
XFILLER_178_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4988_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 VGND VGND VPWR VPWR net339
+ sky130_fd_sc_hd__buf_1
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3939_ _0756_ _0843_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__and2_1
XFILLER_164_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput27 Tile_X0Y0_FrameData[0] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput16 Tile_X0Y0_E2MID[3] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput49 Tile_X0Y0_FrameData[31] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
Xinput38 Tile_X0Y0_FrameData[1] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2270_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q _1257_ _1259_
+ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__o21ai_1
XFILLER_96_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4911_ Tile_X0Y0_E6END[9] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_1
XFILLER_92_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4842_ net172 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1985_ _0984_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__and2_1
X_4773_ net1209 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_165_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3724_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q _0645_ VGND VGND
+ VPWR VPWR _0646_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_119_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3655_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ _0581_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q VGND VGND VPWR
+ VPWR _0582_ sky130_fd_sc_hd__o211a_1
XFILLER_173_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2606_ _1506_ _1558_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__xor2_2
XFILLER_161_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3586_ net98 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q VGND
+ VGND VPWR VPWR _0518_ sky130_fd_sc_hd__mux2_1
X_2537_ _1498_ _1497_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__mux2_1
XFILLER_114_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5256_ Tile_X0Y1_WW4END[11] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__clkbuf_2
X_2468_ _1434_ _1432_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__xor2_4
X_4207_ net41 net1101 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5187_ Tile_X0Y0_S4END[10] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__buf_6
X_2399_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q _1379_ VGND VGND
+ VPWR VPWR _1380_ sky130_fd_sc_hd__nor2_1
X_4138_ net1233 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4069_ net1254 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_126_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1103 net1105 VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__buf_2
XFILLER_160_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1125 net1127 VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__buf_2
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1114 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1147 net1149 VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__buf_2
Xfanout1136 Tile_X0Y1_FrameStrobe[2] VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__buf_4
Xfanout1158 net1161 VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__buf_2
Xfanout1169 net1170 VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__buf_2
XFILLER_120_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3440_ net190 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net226
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux4_2
XFILLER_170_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3371_ _0309_ net739 _0318_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ sky130_fd_sc_hd__a21o_4
XTAP_TAPCELL_ROW_114_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ net973 net968 net987 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR VPWR
+ _1308_ sky130_fd_sc_hd__mux4_1
X_5110_ Tile_X0Y1_E6END[7] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__buf_1
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5041_ net97 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_1
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2253_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ _1243_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__o21ai_1
X_2184_ net1043 net1032 net1008 net1022 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR VPWR
+ _1180_ sky130_fd_sc_hd__mux4_1
XFILLER_111_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4825_ net162 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1968_ _0533_ _0535_ _0125_ _0507_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__a211o_1
X_4756_ net1187 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3707_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q _0629_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q
+ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__o21ba_1
X_4687_ net167 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_173_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3638_ _0561_ _0563_ _0566_ _0073_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ sky130_fd_sc_hd__a22o_4
XFILLER_108_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3569_ net189 net9 net1258 net1256 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q VGND VGND VPWR VPWR
+ _0502_ sky130_fd_sc_hd__mux4_1
XFILLER_108_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput206 Tile_X0Y1_NN4END[5] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_4
Xinput217 Tile_X0Y1_W2END[4] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_2
XFILLER_102_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput228 Tile_X0Y1_W2MID[7] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__buf_2
X_5239_ Tile_X0Y1_W6END[4] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone1 net980 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 _0382_ net672
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q
+ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__mux4_2
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_3__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs VGND VGND VPWR
+ VPWR clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_165_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2940_ _1811_ _1812_ _1813_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q VGND VGND VPWR VPWR
+ _1814_ sky130_fd_sc_hd__a221o_1
X_2871_ net1215 net82 net71 net972 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4610_ net152 net1114 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4541_ net1199 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4472_ net1193 net1174 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3423_ net179 net195 net119 net125 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0367_ sky130_fd_sc_hd__mux4_1
XFILLER_131_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3354_ _0292_ _0279_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_5_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _0135_ _1291_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__nor2_1
X_3285_ net70 net82 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q VGND
+ VGND VPWR VPWR _0236_ sky130_fd_sc_hd__mux2_1
X_5024_ Tile_X0Y1_NN4END[12] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_1
X_2236_ net978 net998 net1019 net1002 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR
+ _1228_ sky130_fd_sc_hd__mux4_1
XFILLER_57_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2167_ _1163_ _1164_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q
+ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__mux2_2
XFILLER_38_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2098_ _0859_ _1098_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__nand2b_1
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4808_ net147 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4739_ net1206 net1079 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_181_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_181_Right_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3070_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q VGND VGND VPWR
+ VPWR _0025_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_78_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2021_ _1003_ _0905_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__xor2_4
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3972_ _0876_ _0861_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A0 sky130_fd_sc_hd__mux2_4
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2923_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q _1797_ _1799_
+ VGND VGND VPWR VPWR _1800_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2854_ net976 _0216_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 _0230_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 sky130_fd_sc_hd__mux4_1
X_2785_ _1698_ _1699_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q
+ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__mux2_1
XFILLER_156_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4524_ net170 net1145 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4455_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C7 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_4386_ net1227 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3406_ _0323_ _0324_ _0348_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a211o_1
X_3337_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q _0284_ _0286_
+ _0058_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__o211a_1
XFILLER_105_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3268_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q _0219_ VGND VGND
+ VPWR VPWR _0220_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_181_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ Tile_X0Y1_N4END[11] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_1
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2219_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q _1207_ _1209_
+ _1211_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q VGND VGND VPWR
+ VPWR _1212_ sky130_fd_sc_hd__a311oi_1
X_3199_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR
+ VPWR _0154_ sky130_fd_sc_hd__inv_1
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput307 net307 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[31] sky130_fd_sc_hd__buf_2
X_2570_ net674 net192 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__mux2_1
Xoutput318 net318 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput329 net329 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
X_4240_ net1241 net1090 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4171_ net1235 net1108 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3122_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q VGND VGND VPWR
+ VPWR _0077_ sky130_fd_sc_hd__inv_2
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3053_ net963 _1616_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__and2b_1
X_2004_ _1004_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__inv_1
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3955_ _0860_ net672 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__mux2_1
XFILLER_50_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2906_ net174 net210 net120 net983 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q VGND VGND VPWR VPWR
+ _1785_ sky130_fd_sc_hd__mux4_1
X_3886_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q _0794_ VGND VGND
+ VPWR VPWR _0795_ sky130_fd_sc_hd__or2_1
XFILLER_176_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2837_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q _1742_ VGND VGND
+ VPWR VPWR _1743_ sky130_fd_sc_hd__and2b_1
X_2768_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q _1683_ _1684_
+ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__a21o_1
X_2699_ net188 net199 net21 net1036 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 sky130_fd_sc_hd__mux4_1
X_4507_ net1197 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4438_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4369_ net39 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer72 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 VGND VGND VPWR VPWR
+ net689 sky130_fd_sc_hd__buf_6
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer94 _0213_ VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3740_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\] net1061 VGND VGND VPWR VPWR _0660_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_13_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3671_ net193 net81 net1216 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q
+ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__mux4_1
XFILLER_173_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2622_ _0146_ _1573_ _1575_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__a21o_1
XFILLER_9_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2553_ _1512_ _1511_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q
+ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__mux2_4
XFILLER_141_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2484_ _1459_ _1157_ _1156_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__a21o_1
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4223_ net1224 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4154_ net1252 net1116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4085_ net1247 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3105_ net18 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__inv_2
XFILLER_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3036_ _1896_ _1897_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q
+ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__mux2_1
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4987_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net338
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3938_ _0756_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__nor2_1
XFILLER_149_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3869_ _0778_ _0779_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q
+ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__mux2_1
XFILLER_164_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 Tile_X0Y0_FrameData[10] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
Xinput17 Tile_X0Y0_E2MID[4] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_10_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput39 Tile_X0Y0_FrameData[20] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_155_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4910_ Tile_X0Y0_E6END[8] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_1
XFILLER_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4841_ net1213 net1157 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1984_ net722 net626 _0983_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__or3_1
XFILLER_60_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4772_ net1208 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_158_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3723_ net58 net66 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q VGND
+ VGND VPWR VPWR _0645_ sky130_fd_sc_hd__mux2_1
XFILLER_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3654_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q _0183_ VGND VGND
+ VPWR VPWR _0581_ sky130_fd_sc_hd__nand2_1
XFILLER_173_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2605_ _1506_ _1558_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__nand2b_1
XFILLER_106_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3585_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q _0516_ VGND VGND
+ VPWR VPWR _0517_ sky130_fd_sc_hd__and2b_1
X_2536_ net188 net8 net85 net100 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q VGND VGND VPWR VPWR
+ _1498_ sky130_fd_sc_hd__mux4_2
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2467_ _1081_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__and2_4
X_5255_ Tile_X0Y1_WW4END[10] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__clkbuf_2
X_4206_ net42 net1100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_87_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5186_ Tile_X0Y0_S4END[9] VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__buf_6
X_2398_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q _1378_ _1376_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q VGND VGND VPWR VPWR
+ _1379_ sky130_fd_sc_hd__o211a_1
X_4137_ net1232 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4068_ net1243 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3019_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q _1882_ _1881_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q VGND VGND VPWR VPWR
+ _1883_ sky130_fd_sc_hd__o211a_1
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1104 net1105 VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__buf_2
Xfanout1126 net1127 VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1115 net1116 VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__clkbuf_2
Xoutput490 net490 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[15] sky130_fd_sc_hd__buf_2
Xfanout1137 net1145 VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__buf_2
Xfanout1159 net1161 VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__buf_2
XFILLER_120_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1148 net1149 VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__buf_1
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3370_ _0311_ _0313_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q
+ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o211a_1
XFILLER_151_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2321_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q VGND VGND VPWR VPWR
+ _1307_ sky130_fd_sc_hd__mux2_1
X_5040_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net391
+ sky130_fd_sc_hd__buf_1
X_2252_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q _0425_ VGND VGND
+ VPWR VPWR _1243_ sky130_fd_sc_hd__nand2_1
XFILLER_2_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2183_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q _1178_ VGND VGND
+ VPWR VPWR _1179_ sky130_fd_sc_hd__nand2b_1
XFILLER_65_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4824_ net1194 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4755_ net1214 net1079 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3706_ net208 net2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q VGND
+ VGND VPWR VPWR _0629_ sky130_fd_sc_hd__mux2_1
X_1967_ _0968_ _0967_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__mux2_4
XFILLER_134_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4686_ net168 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_173_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3637_ _0564_ _0565_ _0072_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__mux2_1
XFILLER_108_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3568_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q _0500_ _0499_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q VGND VGND VPWR VPWR
+ _0501_ sky130_fd_sc_hd__o211a_1
XFILLER_108_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2519_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\]
+ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__and2_1
XFILLER_102_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3499_ net1255 net64 net100 net116 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0437_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_132_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput207 Tile_X0Y1_NN4END[6] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_4
Xinput218 Tile_X0Y1_W2END[5] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput229 Tile_X0Y1_W6END[0] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_4
X_5238_ Tile_X0Y1_W6END[3] VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__clkbuf_2
X_5169_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 VGND VGND VPWR VPWR net520
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2870_ net1016 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 _0382_ net688
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_128_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4540_ net1198 net1130 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_128_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4471_ net163 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3422_ _0022_ _0365_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__a21bo_1
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3353_ _0056_ net965 _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_5_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ net978 net1019 net984 net1014 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q VGND VGND VPWR VPWR
+ _1291_ sky130_fd_sc_hd__mux4_1
X_3284_ net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__a21bo_1
X_5023_ Tile_X0Y1_NN4END[11] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__buf_1
XFILLER_97_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2235_ _1223_ _1225_ _1226_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q
+ _0132_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__o221a_1
X_2166_ net57 net59 net67 net1220 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ _1164_ sky130_fd_sc_hd__mux4_1
XFILLER_38_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2097_ _0841_ _0858_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__nand2_4
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_125_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4807_ net148 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2999_ _1864_ _1863_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 sky130_fd_sc_hd__mux2_1
XFILLER_119_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4738_ net1205 net1079 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_134_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4669_ net1199 net1095 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_134_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_143_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK VGND VGND VPWR VPWR clknet_1_0__leaf_Tile_X0Y1_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_10_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_152_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2020_ _1016_ _1017_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__xor2_4
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_161_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3971_ _0875_ _0862_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_61_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2922_ _0154_ _1798_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q
+ VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__a21o_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2853_ net990 _0196_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 _0173_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 sky130_fd_sc_hd__mux4_1
X_2784_ _0704_ _1522_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q
+ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__mux2_1
XFILLER_116_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4523_ net1180 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_156_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_170_Left_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4454_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C6 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[6\] sky130_fd_sc_hd__dfxtp_1
X_4385_ net1226 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3405_ net738 VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__inv_2
X_3336_ _0057_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__or2_1
XFILLER_112_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5006_ Tile_X0Y1_N4END[10] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__buf_1
X_3267_ net971 net691 net707 net743 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ _0219_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_181_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q _1210_ VGND VGND
+ VPWR VPWR _1211_ sky130_fd_sc_hd__nor2_1
X_3198_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q VGND VGND VPWR
+ VPWR _0153_ sky130_fd_sc_hd__inv_1
XFILLER_38_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2149_ _1147_ _0520_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__mux2_1
XFILLER_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput308 net308 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[3] sky130_fd_sc_hd__buf_2
Xoutput319 net319 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
XFILLER_113_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4170_ net1233 net1108 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3121_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q VGND VGND VPWR
+ VPWR _0076_ sky130_fd_sc_hd__inv_2
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3052_ net963 _1471_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__and2b_1
X_2003_ _1003_ net624 net665 VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_38_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3954_ net183 net129 net92 net219 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q VGND VGND VPWR VPWR
+ _0860_ sky130_fd_sc_hd__mux4_1
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2905_ _1781_ _1784_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A sky130_fd_sc_hd__mux2_1
X_3885_ net971 net967 net990 net976 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0794_ sky130_fd_sc_hd__mux4_1
XFILLER_31_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2836_ net721 _0652_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__mux2_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2767_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q _1682_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q
+ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__o21ai_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2698_ net187 net198 net1255 net1042 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_144_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4506_ net1196 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4437_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4368_ net40 net1161 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3319_ net2 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q VGND
+ VGND VPWR VPWR _0269_ sky130_fd_sc_hd__mux2_1
X_4299_ net1236 net1074 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer40 _1158_ VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer73 net689 VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer95 _0307_ VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3670_ _0593_ _0592_ _0596_ _0101_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1
+ sky130_fd_sc_hd__a22o_4
XFILLER_173_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2621_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q _1574_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q
+ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__a21bo_1
XFILLER_173_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2552_ net17 net109 net73 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q VGND VGND VPWR VPWR
+ _1512_ sky130_fd_sc_hd__mux4_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2483_ _1458_ _1173_ _1172_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__a21o_1
XFILLER_99_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4222_ net1223 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_87_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4153_ net30 net1118 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4084_ net1246 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3104_ net75 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__inv_2
XFILLER_95_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3035_ net221 net658 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__mux4_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4986_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net337
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3937_ _0543_ _0661_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__nor2_1
XFILLER_149_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3868_ net1216 net73 net217 net229 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0779_ sky130_fd_sc_hd__mux4_1
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2819_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q _1726_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__a21bo_1
X_3799_ net708 net724 net750 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0714_ sky130_fd_sc_hd__mux4_2
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 Tile_X0Y0_E2MID[5] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
XFILLER_10_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput29 Tile_X0Y0_FrameData[11] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
XFILLER_10_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_176_Right_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4840_ net147 net1157 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1983_ net722 _0944_ _0983_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__o21ai_1
X_4771_ net1206 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3722_ _0641_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q _0643_
+ _0088_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__o211a_1
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3653_ _0578_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__nand2_1
XFILLER_161_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2604_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\] _1557_ net1058 VGND VGND VPWR VPWR
+ _1558_ sky130_fd_sc_hd__mux2_4
XFILLER_161_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3584_ net1255 net62 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__mux2_1
X_2535_ net199 net87 net99 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q VGND VGND VPWR VPWR
+ _1497_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5254_ Tile_X0Y1_WW4END[9] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__buf_2
X_2466_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\] _1441_ net1057 VGND VGND VPWR VPWR
+ _1442_ sky130_fd_sc_hd__mux2_4
X_5185_ Tile_X0Y0_S4END[8] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__buf_6
X_4205_ net1238 net1100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4136_ net1231 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2397_ _1377_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__inv_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4067_ net1230 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3018_ net997 net1019 net1002 net1014 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q VGND VGND VPWR VPWR
+ _1882_ sky130_fd_sc_hd__mux4_1
XFILLER_36_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4969_ net1109 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput480 net480 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[6] sky130_fd_sc_hd__buf_2
Xfanout1116 net1117 VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__buf_2
XFILLER_154_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1127 Tile_X0Y1_FrameStrobe[3] VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1138 net1140 VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__buf_2
Xoutput491 net491 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[16] sky130_fd_sc_hd__buf_2
Xfanout1105 net1106 VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__buf_2
XFILLER_120_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1149 net1153 VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__clkbuf_2
XFILLER_170_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2320_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q _1305_ VGND VGND
+ VPWR VPWR _1306_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_29_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2251_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 _1241_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR
+ _1242_ sky130_fd_sc_hd__mux4_2
XFILLER_2_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2182_ net1012 net1048 net1027 net1052 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q VGND VGND VPWR VPWR
+ _1178_ sky130_fd_sc_hd__mux4_1
XFILLER_65_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4823_ net163 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1966_ net204 net129 net75 net219 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q VGND VGND VPWR VPWR
+ _0968_ sky130_fd_sc_hd__mux4_1
X_4754_ net1202 net1079 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3705_ _0627_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q VGND VGND
+ VPWR VPWR _0628_ sky130_fd_sc_hd__nand2b_1
XFILLER_119_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4685_ net1182 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3636_ net206 net1257 net6 net1255 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0565_ sky130_fd_sc_hd__mux4_1
X_3567_ net65 net77 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q VGND
+ VGND VPWR VPWR _0500_ sky130_fd_sc_hd__mux2_1
XFILLER_108_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2518_ _1115_ _1480_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__nand2_1
XFILLER_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3498_ _0070_ _0435_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_132_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput208 Tile_X0Y1_NN4END[7] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_4
X_5237_ Tile_X0Y1_W6END[2] VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2449_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q _1426_ VGND VGND
+ VPWR VPWR _1427_ sky130_fd_sc_hd__nor2_1
Xinput219 Tile_X0Y1_W2END[6] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5168_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 VGND VGND VPWR VPWR net519
+ sky130_fd_sc_hd__buf_1
XFILLER_56_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4119_ net1249 net1124 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5099_ net133 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_2
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4470_ net164 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3421_ net972 net985 net991 net976 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0365_ sky130_fd_sc_hd__mux4_2
XFILLER_143_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3352_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q net1004 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q
+ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__o21ba_4
XFILLER_124_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2303_ net973 net968 net987 net992 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR
+ _1290_ sky130_fd_sc_hd__mux4_1
XFILLER_151_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3283_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q net214 VGND VGND
+ VPWR VPWR _0234_ sky130_fd_sc_hd__and2b_1
X_5022_ Tile_X0Y1_NN4END[10] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__buf_1
X_2234_ net175 net1218 net183 net129 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q VGND VGND VPWR VPWR
+ _1226_ sky130_fd_sc_hd__mux4_1
X_2165_ net620 net1258 net191 net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q VGND VGND VPWR VPWR
+ _1163_ sky130_fd_sc_hd__mux4_1
XFILLER_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2096_ _0903_ _1096_ _0901_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__a21o_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4806_ net149 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_166_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2998_ net173 net209 _0410_ net977 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q VGND VGND VPWR VPWR
+ _1864_ sky130_fd_sc_hd__mux4_1
XFILLER_119_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1949_ _0920_ _0945_ _0950_ _0949_ _0948_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__a32oi_1
X_4737_ net153 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4668_ net1198 net1095 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3619_ _0544_ _0108_ _0545_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__a31o_4
XFILLER_88_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4599_ net1192 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3970_ net191 net227 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 net658
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q
+ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__mux4_2
XFILLER_62_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2921_ net176 net1217 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q
+ VGND VGND VPWR VPWR _1798_ sky130_fd_sc_hd__mux2_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2852_ net178 net193 net229 net1016 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A sky130_fd_sc_hd__mux4_1
X_2783_ net1005 _0733_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q
+ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4522_ net1179 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4453_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C5 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3404_ _0324_ _0323_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a21oi_4
X_4384_ net52 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3335_ net199 net7 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q VGND
+ VGND VPWR VPWR _0285_ sky130_fd_sc_hd__mux2_1
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3266_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q net993 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q
+ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5005_ Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__buf_1
X_2217_ net173 net177 net119 net123 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR VPWR
+ _1210_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_181_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q VGND VGND VPWR
+ VPWR _0152_ sky130_fd_sc_hd__inv_2
X_2148_ net190 net86 net10 net102 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q VGND VGND VPWR VPWR
+ _1147_ sky130_fd_sc_hd__mux4_2
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2079_ _1074_ _1077_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput309 net309 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[4] sky130_fd_sc_hd__buf_2
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3120_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q VGND VGND VPWR
+ VPWR _0075_ sky130_fd_sc_hd__inv_2
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3051_ net963 _1470_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__and2b_1
X_2002_ _0997_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__xor2_4
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3953_ _0841_ _0858_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_11_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3884_ _0790_ _0791_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__xor2_1
X_2904_ _1783_ _1782_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q
+ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__mux2_1
XFILLER_31_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2835_ _0149_ _1732_ _1737_ _1741_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0
+ sky130_fd_sc_hd__a31o_1
XFILLER_31_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2766_ net1043 net1038 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__mux2_1
X_2697_ net1035 _0322_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 _0346_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 sky130_fd_sc_hd__mux4_1
X_4505_ net1195 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4436_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\] sky130_fd_sc_hd__dfxtp_1
X_4367_ net41 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3318_ net190 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q VGND VGND
+ VPWR VPWR _0268_ sky130_fd_sc_hd__nand2b_1
XFILLER_116_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4298_ net1234 net1074 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3249_ net1 net5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q VGND
+ VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_92_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer85 _0383_ VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__clkbuf_2
Xrebuffer96 net1049 VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2620_ net1044 net1008 net1038 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q VGND VGND VPWR VPWR
+ _1574_ sky130_fd_sc_hd__mux4_1
XFILLER_9_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2551_ net710 net74 net18 net110 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q VGND VGND VPWR VPWR
+ _1511_ sky130_fd_sc_hd__mux4_2
XFILLER_141_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2482_ _1193_ _1456_ _1274_ _1192_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__a31o_4
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4221_ net55 net1100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4152_ net31 net1118 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4083_ net1245 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3103_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q VGND VGND VPWR
+ VPWR _0058_ sky130_fd_sc_hd__inv_2
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3034_ net191 net131 net137 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__mux4_1
XFILLER_55_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3936_ _0492_ _0709_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__or2_4
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3867_ net175 net181 net193 net127 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0778_ sky130_fd_sc_hd__mux4_1
X_2818_ _1512_ _0540_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q
+ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__mux2_1
X_3798_ _0059_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q
+ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__a21oi_1
XFILLER_164_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2749_ _1664_ _1667_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 sky130_fd_sc_hd__mux2_1
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4419_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0007_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput19 Tile_X0Y0_E2MID[6] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1982_ _0966_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__xnor2_1
X_4770_ net1205 net1071 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3721_ _0087_ _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or2_1
XFILLER_173_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3652_ _0492_ _0576_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__nor2_1
XFILLER_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2603_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[18\] net1064 VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__mux2_2
X_3583_ _0513_ _0512_ _0514_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q VGND VGND VPWR VPWR
+ _0515_ sky130_fd_sc_hd__a221o_1
XFILLER_161_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2534_ _1495_ _0299_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__mux2_4
XFILLER_114_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5253_ Tile_X0Y1_WW4END[8] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__buf_2
X_2465_ Tile_X0Y1_DSP_bot.C0 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[0\] net1063 VGND
+ VGND VPWR VPWR _1441_ sky130_fd_sc_hd__mux2_2
X_4204_ net1237 net1100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5184_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 VGND VGND VPWR VPWR net535
+ sky130_fd_sc_hd__clkbuf_2
X_2396_ net192 net138 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q
+ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__mux2_1
X_4135_ net48 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4066_ net1227 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3017_ _1880_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q VGND VGND
+ VPWR VPWR _1881_ sky130_fd_sc_hd__nand2b_1
XFILLER_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4968_ net1117 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__buf_1
X_4899_ net16 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__buf_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3919_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q _0825_ VGND VGND
+ VPWR VPWR _0826_ sky130_fd_sc_hd__nor2_1
XFILLER_164_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput470 net470 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_160_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1117 net1118 VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1106 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__clkbuf_2
Xoutput492 net492 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[17] sky130_fd_sc_hd__buf_2
XFILLER_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1128 net1136 VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__clkbuf_2
Xoutput481 net481 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1139 net1140 VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__buf_1
XFILLER_170_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2250_ _1235_ _1237_ _1240_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__a22o_1
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2181_ _1176_ _1175_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__mux2_4
XFILLER_77_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4822_ net164 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1965_ net126 net233 net92 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q VGND VGND VPWR VPWR
+ _0967_ sky130_fd_sc_hd__mux4_2
X_4753_ net165 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3704_ net8 net1255 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q VGND
+ VGND VPWR VPWR _0627_ sky130_fd_sc_hd__mux2_1
XFILLER_146_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4684_ net1181 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3635_ net62 net78 net98 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0564_ sky130_fd_sc_hd__mux4_1
XFILLER_108_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3566_ _0498_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q VGND VGND
+ VPWR VPWR _0499_ sky130_fd_sc_hd__nand2b_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3497_ net1036 net1006 net1031 net1054 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0435_ sky130_fd_sc_hd__mux4_1
XFILLER_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2517_ _0843_ _1113_ _1103_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__o21bai_2
XFILLER_142_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5236_ net228 VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__buf_4
X_2448_ net187 net133 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q
+ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__mux2_1
Xinput209 Tile_X0Y1_W1END[0] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_4
XFILLER_68_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5167_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 VGND VGND VPWR VPWR net518
+ sky130_fd_sc_hd__buf_1
X_2379_ net188 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net224
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q
+ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__mux4_2
X_4118_ net1248 net1124 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5098_ net132 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_2
X_4049_ net1242 net1143 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3420_ _0363_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q VGND VGND
+ VPWR VPWR _0364_ sky130_fd_sc_hd__and2_4
X_3351_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net16 net72 net108 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q VGND VGND VPWR VPWR
+ _0299_ sky130_fd_sc_hd__mux4_1
XFILLER_124_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2302_ _1287_ _1289_ _1282_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6
+ sky130_fd_sc_hd__o21ai_4
X_3282_ _0231_ _0232_ _0041_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__mux2_4
X_5021_ Tile_X0Y1_NN4END[9] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__buf_1
X_2233_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q _1224_ _0131_
+ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__a21o_1
XFILLER_38_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2164_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q _1161_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__a21bo_1
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2095_ _1095_ _0954_ _0952_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__a21o_1
XFILLER_80_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4805_ net150 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2997_ _1862_ _1861_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q
+ VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__mux2_1
XFILLER_119_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1948_ _0948_ _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__xor2_1
X_4736_ net154 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_134_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4667_ net160 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3618_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q _0546_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q
+ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__a21bo_1
XFILLER_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4598_ net1191 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3549_ net63 net79 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q VGND
+ VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux2_1
XFILLER_130_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5219_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 VGND VGND VPWR VPWR net570
+ sky130_fd_sc_hd__buf_1
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2920_ _0350_ net990 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q
+ VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__mux2_1
XFILLER_43_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2851_ net177 net196 net230 net997 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A sky130_fd_sc_hd__mux4_1
X_2782_ net621 net1258 net1220 net1025 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q VGND VGND VPWR VPWR
+ _1697_ sky130_fd_sc_hd__mux4_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4521_ net1213 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_156_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4452_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C4 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3403_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2
+ _0347_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q VGND VGND VPWR
+ VPWR _0348_ sky130_fd_sc_hd__o211a_4
XFILLER_171_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4383_ net1224 net1162 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3334_ net744 net187 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_84_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3265_ net711 _0214_ _0215_ _0039_ _0040_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a221o_1
X_5004_ Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_1
X_2216_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q _1208_ VGND VGND
+ VPWR VPWR _1209_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_181_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR
+ VPWR _0151_ sky130_fd_sc_hd__inv_1
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2147_ _1119_ _1142_ _1143_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__a21oi_4
XFILLER_93_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2078_ _1071_ _1067_ _1078_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__nand3_4
XFILLER_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4719_ net1184 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3050_ net963 _1469_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__and2b_1
X_2001_ _0959_ _1000_ _0999_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__a21o_1
XFILLER_90_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3952_ _0855_ _0856_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3883_ _0791_ _0790_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__and2b_1
X_2903_ net1001 _1429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__mux2_1
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2834_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q _1740_ _1739_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q VGND VGND VPWR VPWR
+ _1741_ sky130_fd_sc_hd__o211a_1
XFILLER_176_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2765_ _1681_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__inv_1
XFILLER_129_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4504_ net1194 net1138 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2696_ _1639_ _1638_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 sky130_fd_sc_hd__mux2_1
XFILLER_144_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4435_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.A3 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_4366_ net1239 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3317_ net664 _0218_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ _0242_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a211o_4
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4297_ net1232 net1077 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3248_ _0036_ net617 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3179_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR
+ VPWR _0134_ sky130_fd_sc_hd__inv_1
XFILLER_66_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer86 _0381_ VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_155_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer121 _0349_ VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer110 net966 VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_149_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2550_ _1509_ _1508_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q
+ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__mux2_1
XFILLER_126_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2481_ _1193_ _1456_ _1274_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__and3_1
XFILLER_141_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4220_ net56 net1100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_141_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4151_ net1249 net1118 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_158_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4082_ net1244 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3102_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR
+ VPWR _0057_ sky130_fd_sc_hd__inv_2
XFILLER_95_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3033_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ VGND VGND VPWR VPWR _1895_ sky130_fd_sc_hd__nor2_1
XFILLER_55_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4984_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net335
+ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_34_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3935_ _0840_ _0766_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_167_Left_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3866_ _0776_ _0775_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q
+ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__mux2_4
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2817_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q _1149_ _1724_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q VGND VGND VPWR VPWR
+ _1725_ sky130_fd_sc_hd__a211oi_1
X_3797_ _0354_ _0356_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ _0258_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__a211o_1
X_2748_ _1666_ _1665_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__mux2_1
XFILLER_117_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2679_ _0024_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__a21oi_1
X_4418_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0006_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4349_ net1222 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3720_ net2 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q VGND
+ VGND VPWR VPWR _0642_ sky130_fd_sc_hd__mux2_1
X_1981_ _0492_ net625 VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__nor2_1
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3651_ _0450_ _0543_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__nor2_1
X_2602_ _1556_ _1552_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ sky130_fd_sc_hd__mux2_4
XFILLER_146_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3582_ net198 net24 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q VGND
+ VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux2_1
X_2533_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net107 net71 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q
+ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__mux4_2
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5252_ Tile_X0Y1_WW4END[7] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__clkbuf_2
X_2464_ _1440_ _1438_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C0 sky130_fd_sc_hd__mux2_4
X_4203_ net1235 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5183_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR net534
+ sky130_fd_sc_hd__buf_4
X_2395_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q _1375_ VGND VGND
+ VPWR VPWR _1376_ sky130_fd_sc_hd__nand2_1
X_4134_ net49 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4065_ net1226 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3016_ _0767_ _0940_ _1429_ net1003 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q VGND VGND VPWR VPWR
+ _1880_ sky130_fd_sc_hd__mux4_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4967_ net1126 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4898_ net15 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__buf_1
XFILLER_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3918_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q _0822_ _0824_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q VGND VGND VPWR VPWR
+ _0825_ sky130_fd_sc_hd__o211a_1
XFILLER_138_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3849_ _0760_ _0759_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__nand2_4
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput471 net471 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput460 net460 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[2] sky130_fd_sc_hd__buf_2
Xfanout1107 net1108 VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1118 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__clkbuf_4
Xoutput493 net493 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[18] sky130_fd_sc_hd__buf_2
Xfanout1129 net1136 VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput482 net482 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2180_ net192 net25 net68 net104 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q VGND VGND VPWR VPWR
+ _1176_ sky130_fd_sc_hd__mux4_2
XFILLER_111_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4821_ net1188 net1156 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1964_ _0912_ _0959_ _0960_ _0958_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4752_ net166 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3703_ net64 net100 net80 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q VGND VGND VPWR VPWR
+ _0626_ sky130_fd_sc_hd__mux4_1
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4683_ net1180 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3634_ _0072_ _0562_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__o21a_1
XFILLER_134_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3565_ net101 net117 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux2_1
XFILLER_161_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3496_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q _0433_ VGND VGND
+ VPWR VPWR _0434_ sky130_fd_sc_hd__or2_1
X_2516_ _1118_ _1461_ _1117_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__o21a_1
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5235_ net227 VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__buf_4
X_2447_ _0632_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q VGND VGND
+ VPWR VPWR _1425_ sky130_fd_sc_hd__or2_4
XFILLER_102_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2378_ net187 net223 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q
+ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__mux4_2
X_5166_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 VGND VGND VPWR VPWR net517
+ sky130_fd_sc_hd__clkbuf_1
X_4117_ net34 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5097_ net131 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_2
X_4048_ net1241 net1143 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_104_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput290 net290 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[16] sky130_fd_sc_hd__buf_2
XFILLER_160_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_113_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3350_ _0298_ _0295_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 sky130_fd_sc_hd__mux2_8
X_2301_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q _1288_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q
+ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__o21ai_1
X_5020_ Tile_X0Y1_NN4END[8] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_1
XFILLER_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3281_ net969 net988 net993 net978 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _0232_ sky130_fd_sc_hd__mux4_2
X_2232_ net75 net1068 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__mux2_1
X_2163_ net1043 net1032 net1008 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q VGND VGND VPWR VPWR
+ _1161_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2094_ _0994_ _1094_ _0993_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__a21o_1
XFILLER_80_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4804_ net151 net1164 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_166_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2996_ net714 _1429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__mux2_1
X_4735_ net1201 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1947_ _0895_ _0896_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__xor2_1
XFILLER_174_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4666_ net161 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3617_ net74 net210 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__mux2_1
X_4597_ net1188 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3548_ _0481_ _0480_ _0482_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR VPWR
+ _0483_ sky130_fd_sc_hd__a221o_1
XFILLER_135_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3479_ _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__inv_2
XFILLER_130_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5218_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 VGND VGND VPWR VPWR net569
+ sky130_fd_sc_hd__buf_1
XFILLER_96_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5149_ net1206 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__buf_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_121_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2850_ net180 net139 net195 net983 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_130_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2781_ _1691_ _1696_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1
+ sky130_fd_sc_hd__or2_1
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4520_ net1212 net1137 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_156_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4451_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C3 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_3402_ _0346_ _0074_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2_4
XFILLER_124_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4382_ net1223 net1162 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3333_ _0282_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__a21bo_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3264_ _0213_ _0214_ _0215_ _0039_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a22o_4
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5003_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 VGND VGND VPWR VPWR net354
+ sky130_fd_sc_hd__buf_4
XFILLER_78_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2215_ net89 net231 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__mux2_1
XFILLER_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3195_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q VGND VGND VPWR
+ VPWR _0150_ sky130_fd_sc_hd__inv_1
X_2146_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__inv_2
XFILLER_38_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2077_ _1074_ _1076_ _1072_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__o21a_1
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2979_ net174 net210 net120 net692 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q VGND VGND VPWR VPWR
+ _1848_ sky130_fd_sc_hd__mux4_1
XFILLER_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4718_ net1183 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4649_ net1213 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2000_ _0959_ _1000_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__nand2_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3951_ _0855_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__nor2_1
XFILLER_90_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2902_ net1003 _0921_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__mux2_1
XFILLER_16_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3882_ _0730_ _0731_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2833_ net1006 net1033 net1021 net1054 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR
+ _1740_ sky130_fd_sc_hd__mux4_1
XFILLER_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2764_ net1027 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__mux2_1
XFILLER_129_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4503_ net1192 net1139 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2695_ net1039 net965 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q
+ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__mux2_1
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4434_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.A2 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_4365_ net1238 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3316_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q _0261_ _0265_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q VGND VGND VPWR VPWR
+ _0266_ sky130_fd_sc_hd__o211a_1
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4296_ net1231 net1074 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3247_ _0185_ _0174_ _0197_ _0198_ net617 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__a221o_1
Xrebuffer10 _0394_ VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__buf_6
X_3178_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR
+ VPWR _0133_ sky130_fd_sc_hd__inv_1
XFILLER_73_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2129_ net105 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q
+ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__o21a_1
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer87 net731 VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_179_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer122 _0307_ VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer111 net966 VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2480_ _1453_ _1454_ _1324_ _1275_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__a211o_4
XFILLER_56_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4150_ net1248 net1118 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3101_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q VGND VGND VPWR
+ VPWR _0056_ sky130_fd_sc_hd__inv_2
X_4081_ net1242 net1134 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput190 Tile_X0Y1_N2MID[5] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_4
X_3032_ _1889_ _1887_ _1894_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1
+ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_128_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4983_ Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3934_ _0838_ _0839_ _0837_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__a21bo_4
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3865_ net971 net691 net707 net975 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0776_ sky130_fd_sc_hd__mux4_2
XFILLER_176_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2816_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q net1054 VGND
+ VGND VPWR VPWR _1724_ sky130_fd_sc_hd__nor2_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3796_ _0710_ _0346_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__mux2_1
XFILLER_164_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2747_ net1022 net657 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__mux2_1
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2678_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q net673 VGND VGND
+ VPWR VPWR _1623_ sky130_fd_sc_hd__or2_1
XFILLER_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4417_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0005_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4348_ net1221 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4279_ net1249 net1084 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ Tile_X0Y1_DSP_bot.B0 net1061 _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__o21ai_4
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3650_ _0543_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__nor2_1
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2601_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q _1553_ _1555_
+ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__o21ba_1
X_3581_ _0024_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__a21oi_1
X_2532_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q _1490_ _1494_
+ _1486_ _1484_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6
+ sky130_fd_sc_hd__o32a_4
XFILLER_161_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5251_ Tile_X0Y1_WW4END[6] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__clkbuf_2
X_4202_ net1233 net1099 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_114_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2463_ _1439_ _0216_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__mux2_4
X_5182_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR net533
+ sky130_fd_sc_hd__buf_4
X_2394_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 net228 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q
+ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__mux2_1
X_4133_ net1254 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4064_ net1225 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3015_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q _1877_ _1878_
+ VGND VGND VPWR VPWR _1879_ sky130_fd_sc_hd__a21o_1
XFILLER_36_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4966_ net1135 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_1
XFILLER_149_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4897_ net14 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3917_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q _0823_ VGND VGND
+ VPWR VPWR _0824_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_137_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3848_ _0744_ _0746_ _0758_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__a21o_1
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3779_ _0696_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4
+ sky130_fd_sc_hd__inv_4
XFILLER_138_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput450 net450 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput461 net461 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_160_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1108 net1109 VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__clkbuf_2
Xoutput494 net494 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[19] sky130_fd_sc_hd__buf_2
XFILLER_59_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1119 net1120 VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__clkbuf_2
Xoutput483 net483 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput472 net472 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[13] sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_148_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4820_ net1186 net1156 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1963_ _0962_ _0963_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_16_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ net167 net1080 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3702_ _0624_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__a21bo_1
X_4682_ net1179 net1097 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3633_ net1035 net736 net695 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0562_ sky130_fd_sc_hd__mux4_1
XFILLER_161_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3564_ _0494_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__a21bo_1
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3495_ net1011 net1046 net1050 net1042 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0433_ sky130_fd_sc_hd__mux4_1
XFILLER_142_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2515_ _1478_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 sky130_fd_sc_hd__mux2_4
XFILLER_88_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2446_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5
+ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__nand2_1
X_5234_ net226 VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__clkbuf_2
X_5165_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 VGND VGND VPWR VPWR net516
+ sky130_fd_sc_hd__buf_1
X_4116_ net1246 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2377_ _1357_ _1356_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__xnor2_2
XFILLER_110_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5096_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 VGND VGND VPWR VPWR net447
+ sky130_fd_sc_hd__buf_6
X_4047_ net1240 net1143 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4949_ net1246 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__buf_1
XFILLER_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput280 net280 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_181_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput291 net291 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[17] sky130_fd_sc_hd__buf_2
XFILLER_133_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2300_ net973 net969 net987 net993 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR VPWR
+ _1288_ sky130_fd_sc_hd__mux4_1
X_3280_ net983 net997 net1019 net1014 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _0231_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_131_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2231_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q _1222_ VGND VGND
+ VPWR VPWR _1223_ sky130_fd_sc_hd__and2b_1
X_2162_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q _1159_ VGND VGND
+ VPWR VPWR _1160_ sky130_fd_sc_hd__and2b_1
XFILLER_65_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2093_ _1020_ _1039_ _1091_ _1019_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__a31o_1
XFILLER_80_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4803_ net1207 net1164 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2995_ net1003 _0802_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__mux2_1
X_4734_ net1200 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1946_ _0919_ _0947_ _0918_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__o21ai_1
XFILLER_119_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4665_ net1195 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3616_ _0323_ _0324_ _0348_ _0107_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__a211o_1
X_4596_ net1186 net1113 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3547_ net7 net1256 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q VGND
+ VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux2_1
XFILLER_88_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3478_ net978 net983 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
XFILLER_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5217_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net568
+ sky130_fd_sc_hd__buf_1
X_2429_ net182 net128 net90 net218 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q VGND VGND VPWR VPWR
+ _1408_ sky130_fd_sc_hd__mux4_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5148_ net151 VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__buf_1
XFILLER_151_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5079_ Tile_X0Y0_WW4END[14] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2780_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q _1692_ _1695_
+ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__o21a_1
XFILLER_171_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4450_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C2 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4381_ net1222 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3401_ net208 net115 net80 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q VGND VGND VPWR VPWR
+ _0346_ sky130_fd_sc_hd__mux4_2
X_3332_ net737 net1005 net1030 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0282_ sky130_fd_sc_hd__mux4_2
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3263_ net192 net138 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q
+ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_1
X_3194_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q VGND VGND VPWR
+ VPWR _0149_ sky130_fd_sc_hd__inv_1
X_5002_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 VGND VGND VPWR VPWR net353
+ sky130_fd_sc_hd__buf_2
XFILLER_85_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2214_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q _1206_ VGND VGND
+ VPWR VPWR _1207_ sky130_fd_sc_hd__nand2b_1
X_2145_ _1143_ _1142_ _1119_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__nand3_4
XFILLER_93_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2076_ _1072_ _1076_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2978_ _1844_ _1847_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 sky130_fd_sc_hd__mux2_1
X_1929_ _0929_ _0122_ _0930_ _0932_ _0123_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__a311o_1
X_4717_ net1182 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4648_ net1212 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4579_ net1206 net1122 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3950_ _0580_ _0763_ _0764_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__o21ba_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2901_ net173 net119 net209 net979 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q VGND VGND VPWR VPWR
+ _1781_ sky130_fd_sc_hd__mux4_1
XFILLER_16_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3881_ _0680_ _0786_ _0788_ _0789_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_31_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2832_ _1738_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q VGND VGND
+ VPWR VPWR _1739_ sky130_fd_sc_hd__nand2b_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2763_ _1677_ _1678_ _1679_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q VGND VGND VPWR VPWR
+ _1680_ sky130_fd_sc_hd__a221o_1
XFILLER_144_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4502_ net1191 net1139 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2694_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 _0278_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q
+ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__mux2_1
XFILLER_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4433_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.A1 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_4364_ net1237 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3315_ _0053_ _0262_ _0263_ _0264_ _0054_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a221o_1
XFILLER_112_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4295_ net1229 net1074 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3246_ net745 net725 _0197_ _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a22o_4
X_3177_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q VGND VGND VPWR
+ VPWR _0132_ sky130_fd_sc_hd__inv_1
XFILLER_66_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2128_ _1127_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q VGND VGND
+ VPWR VPWR _1128_ sky130_fd_sc_hd__nand2_2
Xrebuffer55 _0373_ VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_37_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ _1043_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__nand2_2
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer88 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 VGND VGND VPWR VPWR
+ net705 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer77 net658 VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_80_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer112 net728 VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_22_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3100_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR
+ VPWR _0055_ sky130_fd_sc_hd__inv_2
X_4080_ net1241 net1135 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput180 Tile_X0Y1_N2END[3] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_2
X_3031_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q _1893_ _1891_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q VGND VGND VPWR VPWR
+ _1894_ sky130_fd_sc_hd__a211o_1
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput191 Tile_X0Y1_N2MID[6] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_8
XFILLER_48_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4982_ Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3933_ _0835_ _0836_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3864_ net715 net995 net1016 net714 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0775_ sky130_fd_sc_hd__mux4_1
X_2815_ _1723_ _1722_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 sky130_fd_sc_hd__mux2_1
X_3795_ net191 net11 net88 net103 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q VGND VGND VPWR VPWR
+ _0710_ sky130_fd_sc_hd__mux4_2
XFILLER_157_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2746_ net965 _0441_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__mux2_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2677_ _1622_ _1619_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 sky130_fd_sc_hd__mux2_4
XFILLER_132_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput610 net610 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_172_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4416_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0004_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4347_ net1253 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4278_ net1248 net1084 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3229_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q _0180_ _0182_
+ _0178_ _0176_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__o32a_4
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_99_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2600_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q _0696_ _1554_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR
+ _1555_ sky130_fd_sc_hd__o211a_1
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer2 net684 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__buf_6
X_3580_ _0383_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q VGND VGND
+ VPWR VPWR _0512_ sky130_fd_sc_hd__or2_4
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2531_ _0093_ _1493_ _1492_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q
+ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__o211a_1
XFILLER_154_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5250_ Tile_X0Y1_WW4END[5] VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__clkbuf_2
XFILLER_181_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4201_ net1232 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2462_ net191 net227 net137 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__mux4_2
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5181_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR net532
+ sky130_fd_sc_hd__buf_2
XFILLER_68_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2393_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q _1371_ _1373_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q VGND VGND VPWR VPWR
+ _1374_ sky130_fd_sc_hd__a211o_1
XFILLER_122_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4132_ net1243 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4063_ net1224 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3014_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q _1876_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q
+ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4965_ net1143 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__buf_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3916_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net226 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q
+ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__mux2_1
XFILLER_149_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4896_ net13 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
XFILLER_164_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3847_ _0744_ _0746_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__nand3_4
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3778_ _0685_ _0683_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q
+ _0690_ _0695_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__a32o_2
XFILLER_138_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2729_ net965 _0706_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__mux2_1
XFILLER_3_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput440 net440 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput451 net451 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput462 net462 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_160_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1109 net1110 VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__clkbuf_2
Xoutput484 net484 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput473 net473 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[14] sky130_fd_sc_hd__buf_6
Xoutput495 net495 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ _0962_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ net168 net1081 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3701_ net1035 net1005 net1030 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0624_ sky130_fd_sc_hd__mux4_2
X_4681_ net1213 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3632_ _0560_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q VGND VGND
+ VPWR VPWR _0561_ sky130_fd_sc_hd__or2_4
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3563_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q _0495_ VGND VGND
+ VPWR VPWR _0496_ sky130_fd_sc_hd__and2b_1
XFILLER_127_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3494_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\] _0431_ net1058 VGND VGND VPWR VPWR
+ _0432_ sky130_fd_sc_hd__mux2_1
X_2514_ _1459_ _1157_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__xor2_1
XFILLER_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2445_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1422_ _1420_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q VGND VGND VPWR VPWR
+ _1423_ sky130_fd_sc_hd__o211a_1
X_5233_ net225 VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__clkbuf_2
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5164_ net1187 VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkbuf_2
X_4115_ net36 net1125 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2376_ _1357_ _1356_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__and2b_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5095_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 VGND VGND VPWR VPWR net446
+ sky130_fd_sc_hd__buf_6
X_4046_ net1239 net1143 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xclone7 Tile_X0Y1_DSP_bot.A0 net1059 _0877_ VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__o21ai_1
XFILLER_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4948_ net1247 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_2
XFILLER_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4879_ net1184 net1149 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_152_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput270 net270 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[12] sky130_fd_sc_hd__buf_2
XFILLER_133_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput292 net292 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[18] sky130_fd_sc_hd__buf_2
XFILLER_160_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput281 net281 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2230_ _0410_ _0302_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__mux2_1
X_2161_ net1012 net1047 net1027 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ _1159_ sky130_fd_sc_hd__mux4_1
XFILLER_38_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2092_ _1020_ _1091_ _1039_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__and3_1
XFILLER_38_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2994_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q _1860_ _1859_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 sky130_fd_sc_hd__o21a_1
X_4802_ net152 net1164 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_166_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1945_ _0920_ _0945_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__xnor2_1
X_4733_ net1199 net1079 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4664_ net1193 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3615_ _0527_ _0528_ _0522_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__a211o_1
X_4595_ net1214 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3546_ _0049_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a21oi_1
XFILLER_115_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3477_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q _0416_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__o21ba_1
X_5216_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net558
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_130_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2428_ _1404_ _1405_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__xor2_1
XFILLER_96_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2359_ _1090_ _1092_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__xnor2_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5147_ net150 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__buf_1
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5078_ Tile_X0Y0_WW4END[13] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_2
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4029_ net55 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_44_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4380_ net1221 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3400_ _0342_ _0340_ _0345_ _0065_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1
+ sky130_fd_sc_hd__a22o_4
XFILLER_7_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3331_ _0280_ _0058_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__and2_4
XFILLER_124_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3262_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q _0038_ _0039_
+ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a21oi_1
X_3193_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q VGND VGND VPWR
+ VPWR _0148_ sky130_fd_sc_hd__inv_1
XFILLER_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5001_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 VGND VGND VPWR VPWR net352
+ sky130_fd_sc_hd__buf_4
X_2213_ _0410_ _0302_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__mux2_2
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2144_ _1110_ _1100_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__xnor2_4
XFILLER_38_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2075_ _1044_ _1075_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__and2_1
XFILLER_19_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2977_ _1846_ _1845_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q
+ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__mux2_1
X_1928_ net210 _0121_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q
+ _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_62_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4716_ net1181 net1086 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_107_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4647_ net1211 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4578_ net1205 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3529_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q _0463_ VGND VGND
+ VPWR VPWR _0464_ sky130_fd_sc_hd__nor2_1
XFILLER_115_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2900_ _1776_ _1780_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3880_ _0678_ _0787_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2831_ _0733_ net622 _0704_ net965 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q VGND VGND VPWR VPWR
+ _1738_ sky130_fd_sc_hd__mux4_1
XFILLER_31_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2762_ net1012 net1047 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__mux2_1
XFILLER_129_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4501_ net1188 net1139 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2693_ _1637_ _1636_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 sky130_fd_sc_hd__mux2_4
X_4432_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs net735 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4363_ net1235 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3314_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q net1031 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__o21a_1
X_4294_ net1228 net1073 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3245_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q net988 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__o21ba_1
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3176_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q VGND VGND VPWR
+ VPWR _0131_ sky130_fd_sc_hd__inv_2
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2127_ _1127_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5
+ sky130_fd_sc_hd__inv_1
XFILLER_81_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer67 net741 VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__buf_6
Xrebuffer56 net702 VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__buf_6
X_2058_ _0981_ _0676_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__nor2_4
XFILLER_179_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer89 net705 VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer113 net999 VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__buf_2
XFILLER_182_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer124 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 VGND VGND VPWR VPWR
+ net741 sky130_fd_sc_hd__clkbuf_2
XFILLER_135_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_118_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput170 Tile_X0Y1_FrameData[7] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_2
Xinput181 Tile_X0Y1_N2END[4] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
X_3030_ _1892_ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__inv_1
XFILLER_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput192 Tile_X0Y1_N2MID[7] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_127_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4981_ Tile_X0Y1_FrameStrobe[17] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3932_ _0577_ _0831_ _0833_ _0830_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3863_ _0770_ _0771_ _0774_ _0114_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2814_ net744 net93 net57 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q VGND VGND VPWR VPWR
+ _1723_ sky130_fd_sc_hd__mux4_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3794_ net1061 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ _0708_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__o21ai_4
X_2745_ net744 net57 net1 net1043 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _1664_ sky130_fd_sc_hd__mux4_1
XFILLER_117_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2676_ _1620_ _1621_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q
+ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__mux2_4
Xoutput600 net600 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput611 net611 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_132_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4415_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0003_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4346_ net1252 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4277_ net1247 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3228_ _0031_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__nor2_1
XFILLER_27_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3159_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q VGND VGND VPWR
+ VPWR _0114_ sky130_fd_sc_hd__inv_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer3 net619 VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_139_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2530_ net68 net1219 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__mux2_1
XFILLER_158_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2461_ _1437_ _1436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__mux2_1
XFILLER_114_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4200_ net1231 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5180_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR net531
+ sky130_fd_sc_hd__buf_4
X_2392_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q _1372_ VGND VGND
+ VPWR VPWR _1373_ sky130_fd_sc_hd__and2b_1
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4131_ net1230 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4062_ net1223 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3013_ net978 net983 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__mux2_1
X_4964_ net1176 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3915_ _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__inv_1
X_4895_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 VGND VGND VPWR VPWR net246
+ sky130_fd_sc_hd__buf_1
XFILLER_149_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3846_ _0757_ _0754_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__xnor2_4
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3777_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q _0694_ VGND VGND
+ VPWR VPWR _0695_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2728_ net1022 net657 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__mux2_1
XFILLER_160_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2659_ _1609_ _1506_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__xnor2_2
Xoutput430 net430 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput441 net441 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput452 net452 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[4] sky130_fd_sc_hd__buf_2
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput496 net496 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput474 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 VGND VGND VPWR VPWR
+ Tile_X0Y1_EE4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput463 net463 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput485 net485 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[10] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4329_ net1232 net1169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3700_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q _0622_ VGND VGND
+ VPWR VPWR _0623_ sky130_fd_sc_hd__and2b_1
X_1961_ _0909_ _0915_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_16_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4680_ net1212 net1094 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3631_ net724 net750 net1049 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0560_ sky130_fd_sc_hd__mux4_2
X_3562_ net1009 net1045 net750 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ _0495_ sky130_fd_sc_hd__mux4_2
XFILLER_127_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2513_ _1477_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 sky130_fd_sc_hd__mux2_4
XFILLER_154_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3493_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[14\] net1064 VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2444_ _1421_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__inv_2
X_5232_ net224 VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__buf_1
X_2375_ _1089_ _1055_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__xnor2_2
X_5163_ net1189 VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkbuf_2
X_4114_ net37 net1127 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5094_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 VGND VGND VPWR VPWR net445
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4045_ net43 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone8 net1061 Tile_X0Y1_DSP_bot.B0 _0980_ VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_67_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4947_ net33 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_2
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4878_ net1183 net1149 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3829_ net665 _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__or2_1
XFILLER_180_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput260 net260 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput271 net271 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[13] sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_7_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput293 net293 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[19] sky130_fd_sc_hd__buf_2
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput282 net282 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net16 net72 net108 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q VGND VGND VPWR VPWR
+ _1158_ sky130_fd_sc_hd__mux4_2
XFILLER_93_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2091_ _1021_ _1038_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__xor2_2
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2993_ net176 net1067 _0350_ net990 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q VGND VGND VPWR VPWR
+ _1860_ sky130_fd_sc_hd__mux4_1
X_4801_ net1204 net1164 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_159_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1944_ _0920_ _0945_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__nand2_2
X_4732_ net1198 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4663_ net163 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3614_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ net1060 _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__o21ai_4
XFILLER_174_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4594_ net1202 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3545_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q _0199_ VGND VGND
+ VPWR VPWR _0480_ sky130_fd_sc_hd__or2_1
XFILLER_115_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3476_ net173 net177 net119 net141 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR VPWR
+ _0416_ sky130_fd_sc_hd__mux4_1
XFILLER_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2427_ _1405_ _1404_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__nand2b_4
X_5215_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net557
+ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_4_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2358_ net1057 _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__nand2_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5146_ net149 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__buf_1
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5077_ Tile_X0Y0_WW4END[12] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_2
XFILLER_96_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2289_ _0349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q _1276_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR VPWR
+ _1277_ sky130_fd_sc_hd__a211o_1
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4028_ net1221 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3330_ net708 net750 net723 net1041 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0280_ sky130_fd_sc_hd__mux4_2
XFILLER_124_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5000_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 VGND VGND VPWR VPWR net351
+ sky130_fd_sc_hd__buf_4
X_3261_ _0204_ _0206_ _0212_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q
+ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a211o_1
X_3192_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q VGND VGND VPWR
+ VPWR _0147_ sky130_fd_sc_hd__inv_1
X_2212_ _1200_ _1201_ _1205_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5
+ sky130_fd_sc_hd__o21a_1
X_2143_ net1058 _1141_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__nand2_4
XFILLER_78_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2074_ _1059_ _1073_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__xor2_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2976_ net693 _1429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__mux2_1
X_1927_ net74 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q VGND VGND
+ VPWR VPWR _0931_ sky130_fd_sc_hd__or2_1
X_4715_ net1180 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_32_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4646_ net1210 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4577_ net1204 net1122 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3528_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net9 net189 net1256 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q VGND VGND VPWR VPWR
+ _0463_ sky130_fd_sc_hd__mux4_1
XFILLER_115_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3459_ net1010 net724 net1024 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0400_ sky130_fd_sc_hd__mux4_2
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5129_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 VGND VGND VPWR VPWR net471
+ sky130_fd_sc_hd__buf_1
XFILLER_84_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2830_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q _1735_ _1736_
+ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__a21o_1
XFILLER_91_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2761_ net1257 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__o21ba_1
X_2692_ net1050 _0526_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q
+ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__mux2_4
XFILLER_129_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4500_ net1186 net1139 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_61_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4431_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0019_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4362_ net1233 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3313_ net1021 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q VGND
+ VGND VPWR VPWR _0263_ sky130_fd_sc_hd__nand2b_1
XFILLER_112_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4293_ net1254 net1085 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3244_ _0193_ _0194_ _0195_ _0028_ _0029_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a221o_1
XFILLER_58_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1090 net1091 VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__clkbuf_2
X_3175_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR
+ VPWR _0130_ sky130_fd_sc_hd__inv_1
X_2126_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q _1126_ _1123_
+ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__o21ai_4
Xrebuffer46 _0217_ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__clkbuf_2
Xrebuffer57 net673 VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__dlygate4sd1_1
X_2057_ _1000_ _1044_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__a21o_1
XFILLER_25_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2959_ net986 net976 net990 net692 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q VGND VGND VPWR VPWR
+ _1832_ sky130_fd_sc_hd__mux4_1
XFILLER_41_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer125 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 VGND VGND VPWR VPWR net742
+ sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer114 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 VGND VGND VPWR VPWR net731
+ sky130_fd_sc_hd__buf_6
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4629_ net1188 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_173_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput160 Tile_X0Y1_FrameData[24] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
Xinput171 Tile_X0Y1_FrameData[8] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_2
XFILLER_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput193 Tile_X0Y1_N4END[0] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput182 Tile_X0Y1_N2END[5] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_2
XFILLER_48_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4980_ Tile_X0Y1_FrameStrobe[16] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3931_ _0835_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__nand2b_1
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3862_ _0772_ _0773_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q
+ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__mux2_1
X_2813_ _1720_ _1721_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q
+ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3793_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\] net1061 VGND VGND VPWR VPWR _0708_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2744_ _1663_ _1662_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 sky130_fd_sc_hd__mux2_1
XFILLER_117_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2675_ net59 net67 net93 net1220 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR
+ _1621_ sky130_fd_sc_hd__mux4_1
XFILLER_8_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput601 net601 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[10] sky130_fd_sc_hd__buf_2
XFILLER_172_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput612 net612 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[6] sky130_fd_sc_hd__buf_2
X_4414_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0002_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4345_ net1251 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4276_ net1246 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3227_ net73 net81 net217 net229 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0181_ sky130_fd_sc_hd__mux4_1
XFILLER_94_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3158_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q VGND VGND VPWR
+ VPWR _0113_ sky130_fd_sc_hd__inv_1
XFILLER_39_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2109_ _1109_ _1101_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__xnor2_4
XFILLER_94_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3089_ net20 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer4 net619 VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2460_ net184 net143 net76 net220 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q VGND VGND VPWR VPWR
+ _1437_ sky130_fd_sc_hd__mux4_1
XFILLER_174_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4130_ net1227 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2391_ net191 net137 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q
+ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__mux2_1
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4061_ net1222 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3012_ _1875_ VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__inv_1
XFILLER_36_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4963_ net1228 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3914_ net190 net136 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q
+ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__mux2_1
X_4894_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 VGND VGND VPWR VPWR net245
+ sky130_fd_sc_hd__buf_1
XFILLER_137_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3845_ _0743_ _0755_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3776_ _0086_ _0693_ _0692_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q
+ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__o211a_1
X_2727_ _1649_ _1650_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 sky130_fd_sc_hd__mux2_1
XFILLER_172_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput420 net420 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_160_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2658_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\] _1608_ net1058 VGND VGND VPWR VPWR
+ _1609_ sky130_fd_sc_hd__mux2_4
Xoutput431 net431 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_105_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput442 net442 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput453 net453 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[5] sky130_fd_sc_hd__buf_2
XFILLER_160_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2589_ _1506_ _1543_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__nand2b_1
Xoutput486 net486 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput475 net475 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput464 net464 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4328_ net1231 net1169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput497 net497 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[21] sky130_fd_sc_hd__buf_2
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4259_ net1230 net1092 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_146_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_155_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_164_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1960_ _0957_ _0961_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3630_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q net221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q
+ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__o21a_1
X_3561_ net1036 net1006 net1031 net1021 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ _0494_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_136_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_180_Right_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2512_ _1476_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__inv_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3492_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q _0254_ _0393_
+ _0430_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_173_Left_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5231_ net223 VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__clkbuf_2
X_2443_ net180 net126 net72 net232 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q VGND VGND VPWR VPWR
+ _1421_ sky130_fd_sc_hd__mux4_1
XFILLER_68_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2374_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\] _1355_ net1057 VGND VGND VPWR VPWR
+ _1356_ sky130_fd_sc_hd__mux2_4
X_5162_ net164 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__buf_1
X_4113_ net1242 net1126 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5093_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 VGND VGND VPWR VPWR net444
+ sky130_fd_sc_hd__buf_1
XFILLER_110_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4044_ net44 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone9 Tile_X0Y1_DSP_bot.B1 net1061 _0943_ VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__o21ai_4
XPHY_EDGE_ROW_182_Left_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4946_ net32 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__buf_2
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4877_ net1182 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_137_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3828_ net1059 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ _0739_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__o21ai_4
XFILLER_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3759_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__inv_2
XFILLER_145_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput261 net261 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput250 net250 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[3] sky130_fd_sc_hd__buf_2
XFILLER_133_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput294 net294 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput283 net283 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput272 net272 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_59_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2090_ _1021_ _1038_ _1055_ _1089_ _1054_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__a221o_1
XFILLER_38_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ net1203 net1166 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_72_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2992_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q _1856_ _1857_
+ _1858_ _0156_ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__a221o_1
X_1943_ net626 _0492_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__nor2_4
X_4731_ net1197 net1078 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4662_ net164 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3613_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\] net1060 VGND VGND VPWR VPWR _0542_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_174_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4593_ net1190 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3544_ _0478_ _0050_ _0477_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q
+ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__o211a_1
XFILLER_115_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3475_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0412_ _0411_
+ _0414_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q VGND VGND VPWR
+ VPWR _0415_ sky130_fd_sc_hd__o311ai_4
XFILLER_142_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2426_ _1080_ _1084_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__xnor2_1
X_5214_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR net556
+ sky130_fd_sc_hd__buf_4
XFILLER_130_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5145_ net1211 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__buf_4
X_2357_ Tile_X0Y1_DSP_bot.C7 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[7\] net1063 VGND
+ VGND VPWR VPWR _1340_ sky130_fd_sc_hd__mux2_4
XFILLER_151_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5076_ Tile_X0Y0_WW4END[11] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_2
X_2288_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q _0529_ VGND VGND
+ VPWR VPWR _1276_ sky130_fd_sc_hd__nor2_2
XFILLER_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4027_ net1253 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4929_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 VGND VGND VPWR VPWR net271
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_165_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3260_ _0206_ _0204_ _0212_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7
+ sky130_fd_sc_hd__a21o_4
X_3191_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q VGND VGND VPWR
+ VPWR _0146_ sky130_fd_sc_hd__inv_2
Xfanout1250 net31 VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__buf_4
X_2211_ _1202_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q _1204_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q VGND VGND VPWR VPWR
+ _1205_ sky130_fd_sc_hd__a211o_1
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2142_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[13\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q
+ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__mux2_4
XFILLER_93_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2073_ _1059_ _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__and2_1
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4714_ net1179 net1087 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2975_ net1003 _0571_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__mux2_1
X_1926_ _0527_ _0528_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ _0522_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_32_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4645_ net1209 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4576_ net1203 net1121 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3527_ _0461_ _0082_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__o21ai_2
XFILLER_115_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3458_ _0394_ _0395_ _0397_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q VGND VGND VPWR VPWR
+ _0399_ sky130_fd_sc_hd__o221a_4
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3389_ net1009 net1045 net1049 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0336_ sky130_fd_sc_hd__mux4_2
X_2409_ _1388_ _1387_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__nor2_4
XFILLER_84_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5128_ Tile_X0Y1_EE4END[15] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__buf_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5059_ Tile_X0Y0_W6END[4] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkbuf_2
XFILLER_55_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2760_ net1219 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q VGND
+ VGND VPWR VPWR _1677_ sky130_fd_sc_hd__nand2b_1
XFILLER_129_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2691_ _1635_ _0520_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q
+ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__mux2_1
XFILLER_144_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4430_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0018_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_4361_ net45 net1160 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3312_ net1036 net1006 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__mux2_1
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4292_ net1243 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3243_ _0193_ _0194_ _0195_ _0028_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__a22o_2
XFILLER_66_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1091 net1092 VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__buf_2
X_3174_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR
+ VPWR _0129_ sky130_fd_sc_hd__inv_1
Xfanout1080 net1081 VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__clkbuf_2
X_2125_ _1124_ _1125_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q
+ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__mux2_4
XFILLER_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer58 net673 VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer47 net663 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__dlygate4sd1_1
X_2056_ _0785_ _0829_ _1024_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_37_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer104 _0537_ VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_20_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2958_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q _1830_ VGND
+ VGND VPWR VPWR _1831_ sky130_fd_sc_hd__nor2_1
XFILLER_175_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1909_ _0889_ _0911_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__xnor2_1
Xrebuffer115 net731 VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4628_ net1186 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2889_ net175 net1218 net1068 net987 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q VGND VGND VPWR VPWR
+ _1771_ sky130_fd_sc_hd__mux4_1
XFILLER_135_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4559_ net1184 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput161 Tile_X0Y1_FrameData[25] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_2
Xinput150 Tile_X0Y1_FrameData[14] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_2
Xinput172 Tile_X0Y1_FrameData[9] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_2
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput194 Tile_X0Y1_N4END[1] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
Xinput183 Tile_X0Y1_N2END[6] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_4
X_3930_ _0750_ _0752_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__xor2_1
XFILLER_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3861_ net1216 net71 net215 net234 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0773_ sky130_fd_sc_hd__mux4_1
X_3792_ _0705_ _0707_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ sky130_fd_sc_hd__mux2_4
X_2812_ net965 _0634_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__mux2_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2743_ net618 net1257 net60 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q VGND VGND VPWR VPWR
+ _1663_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_139_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2674_ net619 net1258 net191 net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q VGND VGND VPWR VPWR
+ _1620_ sky130_fd_sc_hd__mux4_2
Xoutput602 net602 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_172_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput613 net613 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[7] sky130_fd_sc_hd__buf_2
X_4413_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0001_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4344_ net1250 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4275_ net1245 net1082 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3226_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q _0179_ VGND VGND
+ VPWR VPWR _0180_ sky130_fd_sc_hd__nor2_1
XFILLER_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3157_ net201 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_146_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ _1108_ _0851_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__xnor2_4
XFILLER_54_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3088_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR
+ VPWR _0043_ sky130_fd_sc_hd__inv_2
XFILLER_153_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2039_ _1037_ _1036_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_59_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer5 _1158_ VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2390_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q VGND VGND VPWR VPWR
+ _1371_ sky130_fd_sc_hd__mux2_1
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4060_ net1221 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_95_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3011_ net988 net993 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__mux2_1
X_4962_ net1229 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4893_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 VGND VGND VPWR VPWR net244
+ sky130_fd_sc_hd__buf_4
X_3913_ _0117_ _0805_ _0817_ _0816_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q
+ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__a221o_1
XFILLER_149_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3844_ _0620_ _0740_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__nor2_1
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3775_ net66 net94 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q VGND
+ VGND VPWR VPWR _0693_ sky130_fd_sc_hd__mux2_1
X_2726_ net1031 net721 _0652_ _1166_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q VGND VGND VPWR VPWR
+ _1650_ sky130_fd_sc_hd__mux4_1
XFILLER_160_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2657_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\] net1064 VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__mux2_4
Xoutput410 net410 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[11] sky130_fd_sc_hd__buf_6
XFILLER_160_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput421 net421 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput432 net432 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_105_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput443 net443 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2588_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q _1543_ _1481_
+ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__and3_1
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput487 net487 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput454 net454 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput476 net476 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput465 net465 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[7] sky130_fd_sc_hd__buf_2
X_4327_ net1229 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput498 net498 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[22] sky130_fd_sc_hd__buf_2
X_4258_ net1227 net1092 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3209_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q _0163_ VGND VGND
+ VPWR VPWR _0164_ sky130_fd_sc_hd__or2_4
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4189_ net55 net1109 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_107_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_177_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3560_ _0450_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2511_ _1174_ _1458_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__xor2_2
XFILLER_142_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3491_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q _0429_ VGND VGND
+ VPWR VPWR _0430_ sky130_fd_sc_hd__nor2_1
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5230_ net222 VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__buf_1
XFILLER_142_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2442_ _0138_ _1417_ _1419_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2373_ Tile_X0Y1_DSP_bot.C6 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[6\] net1063 VGND
+ VGND VPWR VPWR _1355_ sky130_fd_sc_hd__mux2_1
X_5161_ net163 VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_2
X_4112_ net40 net1126 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5092_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 VGND VGND VPWR VPWR net443
+ sky130_fd_sc_hd__clkbuf_2
X_4043_ net1235 net1142 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4945_ net31 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_2
XFILLER_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4876_ net1181 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3827_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\] net1059 VGND VGND VPWR VPWR _0739_
+ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3758_ Tile_X0Y1_DSP_bot.A2 net1059 _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_154_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2709_ _1644_ _1645_ _0068_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__mux2_1
XFILLER_152_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3689_ _0063_ _0609_ _0613_ _0605_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2
+ sky130_fd_sc_hd__a31o_1
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput262 net262 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput251 net251 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput240 net240 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput295 net295 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput284 net284 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[10] sky130_fd_sc_hd__buf_2
XFILLER_160_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput273 net273 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[15] sky130_fd_sc_hd__buf_6
XFILLER_133_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2991_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q net733 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q
+ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__o21ba_1
XFILLER_159_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4730_ net1196 net1081 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1942_ Tile_X0Y1_DSP_bot.B1 net1061 _0943_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__o21ai_4
XPHY_EDGE_ROW_14_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4661_ net1188 net1095 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3612_ _0538_ _0541_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_12_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4592_ net1185 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3543_ net737 net736 net1029 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0478_ sky130_fd_sc_hd__mux4_2
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3474_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q _0413_ VGND VGND
+ VPWR VPWR _0414_ sky130_fd_sc_hd__nand2_1
X_2425_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\] _1403_ net1057 VGND VGND VPWR VPWR
+ _1404_ sky130_fd_sc_hd__mux2_4
X_5213_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net555
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5144_ net1212 VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__buf_4
XFILLER_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2356_ _0137_ _1334_ _1339_ _1330_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C7 sky130_fd_sc_hd__a31o_4
X_5075_ Tile_X0Y0_WW4END[10] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_2
XFILLER_96_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2287_ _1194_ _1271_ _1272_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__o21a_1
XFILLER_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4026_ net1252 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4928_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 VGND VGND VPWR VPWR net270
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4859_ net1197 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2210_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q _1203_ VGND VGND
+ VPWR VPWR _1204_ sky130_fd_sc_hd__and2b_1
Xfanout1240 net41 VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__buf_4
X_3190_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR
+ VPWR _0145_ sky130_fd_sc_hd__inv_2
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1251 net30 VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__buf_4
X_2141_ _1137_ _1131_ _1140_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2072_ _0785_ _0944_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__nor2_1
XFILLER_75_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2974_ net173 net119 net209 net976 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q VGND VGND VPWR VPWR
+ _1844_ sky130_fd_sc_hd__mux4_1
X_1925_ _0323_ _0324_ _0121_ _0348_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__a211o_1
X_4713_ net1213 net1088 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_32_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4644_ net1208 net1104 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4575_ net156 net1122 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_162_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3526_ net737 net1005 net1029 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0461_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_31_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3457_ _0395_ net627 _0397_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q
+ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o22ai_4
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3388_ net1034 net1004 net695 net676 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0335_ sky130_fd_sc_hd__mux4_1
XFILLER_69_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2408_ _1087_ _1386_ _1385_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__a21oi_1
X_2339_ _1093_ _1322_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__nor2_4
X_5127_ Tile_X0Y1_EE4END[14] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__buf_1
XFILLER_29_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5058_ Tile_X0Y0_W6END[3] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4009_ net1232 net1178 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_40_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2690_ _0048_ _1626_ _1630_ _1634_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__a31o_1
XFILLER_129_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4360_ net46 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3311_ net1011 net1046 net1026 net1050 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR
+ _0261_ sky130_fd_sc_hd__mux4_1
X_4291_ net47 net1083 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3242_ net186 net132 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q
+ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3173_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q VGND VGND VPWR
+ VPWR _0128_ sky130_fd_sc_hd__inv_2
X_2124_ net57 net59 net67 net95 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR
+ _1125_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_175_Right_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1081 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__clkbuf_4
Xfanout1092 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1070 net1072 VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__clkbuf_4
XFILLER_81_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2055_ _1051_ _1050_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__xor2_1
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2957_ net1218 net1068 net972 net967 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q VGND VGND VPWR VPWR
+ _1830_ sky130_fd_sc_hd__mux4_1
XFILLER_41_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1908_ _0601_ _0575_ _0574_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__and3b_1
X_2888_ net971 _0382_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 net688
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_30_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4627_ net1214 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4558_ net1183 net1128 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_173_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3509_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q _0443_ _0445_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q VGND VGND VPWR VPWR
+ _0446_ sky130_fd_sc_hd__o211a_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4489_ net1213 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_106_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput162 Tile_X0Y1_FrameData[26] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_2
Xinput151 Tile_X0Y1_FrameData[15] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_2
Xinput140 Tile_X0Y1_E6END[1] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
Xinput195 Tile_X0Y1_N4END[2] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
Xinput184 Tile_X0Y1_N2END[7] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_4
Xinput173 Tile_X0Y1_N1END[0] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_4
XFILLER_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3860_ net173 net179 net195 net125 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0772_ sky130_fd_sc_hd__mux4_1
XFILLER_176_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3791_ _0706_ _0398_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q
+ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__mux2_4
X_2811_ net676 net623 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2742_ net1032 net721 _0652_ _1176_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q VGND VGND VPWR VPWR
+ _1662_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_139_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2673_ _1617_ _1618_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q
+ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__mux2_4
XFILLER_172_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4412_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0000_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput614 net614 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput603 net603 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[12] sky130_fd_sc_hd__buf_2
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4343_ net32 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4274_ net1244 net1083 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3225_ net175 net181 net127 net1216 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0179_ sky130_fd_sc_hd__mux4_1
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3156_ net213 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_1
X_3087_ net188 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
X_2107_ _1105_ _1106_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__or2_1
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _1038_ _1021_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__or2_4
XPHY_EDGE_ROW_6_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3989_ _0793_ _0834_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__xor2_1
XFILLER_10_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer6 _1158_ VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3010_ _1871_ _1872_ _1873_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q VGND VGND VPWR VPWR
+ _1874_ sky130_fd_sc_hd__a221o_1
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4961_ net1231 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__buf_1
XFILLER_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4892_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 VGND VGND VPWR VPWR net243
+ sky130_fd_sc_hd__buf_1
X_3912_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__inv_2
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3843_ _0661_ _0740_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK VGND VGND VPWR VPWR clknet_0_Tile_X0Y1_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
X_3774_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q _0691_ VGND VGND
+ VPWR VPWR _0692_ sky130_fd_sc_hd__or2_1
X_2725_ net618 net1219 net1257 net1050 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q VGND VGND VPWR VPWR
+ _1649_ sky130_fd_sc_hd__mux4_1
XFILLER_172_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2656_ _0147_ _1593_ _1607_ _1579_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput411 net411 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput400 net400 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput422 net422 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput433 net433 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput444 net444 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_160_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2587_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\] _1542_ net1058 VGND VGND VPWR VPWR
+ _1543_ sky130_fd_sc_hd__mux2_4
XFILLER_113_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput477 net477 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput455 net455 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput466 net466 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4326_ net1228 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput499 net499 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput488 net488 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[13] sky130_fd_sc_hd__buf_2
X_4257_ net51 net1092 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4188_ net56 net1109 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3208_ net971 net966 net991 net977 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0163_ sky130_fd_sc_hd__mux4_2
X_3139_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q VGND VGND VPWR
+ VPWR _0094_ sky130_fd_sc_hd__inv_2
XFILLER_103_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_177_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3490_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q _0426_ _0428_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q VGND VGND VPWR VPWR
+ _0429_ sky130_fd_sc_hd__o211a_1
X_2510_ _1475_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\] net1066 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 sky130_fd_sc_hd__mux2_4
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2441_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q _1418_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q
+ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__o21a_1
XFILLER_142_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5160_ net1194 VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__buf_2
X_2372_ _1354_ _1348_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C6 sky130_fd_sc_hd__mux2_4
X_4111_ net1240 net1126 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5091_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 VGND VGND VPWR VPWR net442
+ sky130_fd_sc_hd__clkbuf_2
X_4042_ net1233 net1143 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4944_ net30 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_96_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4875_ net1180 net1147 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_15_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3826_ _0735_ _0738_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ sky130_fd_sc_hd__mux2_2
X_3757_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\] net1059 VGND VGND VPWR VPWR _0675_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_165_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2708_ net186 net198 net4 net6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _1645_ sky130_fd_sc_hd__mux4_1
XFILLER_160_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3688_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q _0612_ _0611_
+ _0062_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__a211o_1
X_2639_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q VGND VGND VPWR VPWR
+ _1592_ sky130_fd_sc_hd__mux2_1
Xoutput252 net252 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput241 net241 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput285 net285 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[11] sky130_fd_sc_hd__buf_2
XFILLER_160_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput263 net263 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput274 net274 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_99_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput296 net296 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[21] sky130_fd_sc_hd__buf_2
X_4309_ net34 net1076 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2990_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q _0662_ VGND VGND
+ VPWR VPWR _1857_ sky130_fd_sc_hd__nand2_1
XFILLER_159_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1941_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\] net1061 VGND VGND VPWR VPWR _0943_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_159_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4660_ net1186 net1095 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_174_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3611_ _0540_ _0539_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q
+ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4591_ net1184 net1120 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3542_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q _0476_ VGND VGND
+ VPWR VPWR _0477_ sky130_fd_sc_hd__or2_4
XFILLER_142_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3473_ net209 net1068 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
X_5212_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net554
+ sky130_fd_sc_hd__buf_6
XFILLER_142_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2424_ Tile_X0Y1_DSP_bot.C3 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[3\] net1063 VGND
+ VGND VPWR VPWR _1403_ sky130_fd_sc_hd__mux2_4
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5143_ net1213 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__buf_2
X_2355_ _1335_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q _1338_
+ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__a21o_1
XFILLER_96_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5074_ Tile_X0Y0_WW4END[9] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkbuf_2
X_2286_ net616 VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__inv_2
XFILLER_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4025_ net1251 net1178 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4927_ Tile_X0Y0_EE4END[15] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
XFILLER_100_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4858_ net1196 net1146 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3809_ _0425_ _0044_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q
+ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__mux2_1
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4789_ net1188 net1165 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1241 net40 VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__buf_4
Xfanout1230 net47 VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__buf_4
XFILLER_78_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2140_ _1139_ _1138_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__mux2_4
Xfanout1252 net29 VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__buf_4
XFILLER_78_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2071_ _1058_ _1062_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__xor2_1
XFILLER_81_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2973_ _1839_ _1843_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 sky130_fd_sc_hd__mux2_1
X_1924_ _0923_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _0925_
+ _0927_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q VGND VGND VPWR
+ VPWR _0928_ sky130_fd_sc_hd__o221a_1
X_4712_ net1212 net1089 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4643_ net1207 net1103 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4574_ net157 net1122 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_151_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3525_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q _0459_ VGND VGND
+ VPWR VPWR _0460_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3456_ net199 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q _0396_
+ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__o21ai_2
XFILLER_162_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3387_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0331_ _0333_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR VPWR
+ _0334_ sky130_fd_sc_hd__o211a_1
XFILLER_69_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2407_ _1087_ _1385_ _1386_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_179_Left_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2338_ _1039_ _1091_ _1020_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5126_ Tile_X0Y1_EE4END[13] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__buf_1
X_5057_ Tile_X0Y0_W6END[2] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkbuf_2
X_2269_ _0129_ _1258_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__o21a_1
XFILLER_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4008_ net46 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3310_ net1256 _0052_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4290_ net50 net1083 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3241_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q _0027_ _0028_
+ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__a21oi_1
X_3172_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q VGND VGND VPWR
+ VPWR _0127_ sky130_fd_sc_hd__inv_1
XFILLER_66_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2123_ net619 net1258 net191 net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q VGND VGND VPWR VPWR
+ _1124_ sky130_fd_sc_hd__mux4_2
Xfanout1082 net1085 VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__buf_2
Xfanout1060 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q VGND VGND
+ VPWR VPWR net1060 sky130_fd_sc_hd__buf_2
Xfanout1071 net1072 VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__buf_2
Xfanout1093 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__clkbuf_2
X_2054_ _1053_ _1040_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__xnor2_4
Xrebuffer49 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 VGND VGND VPWR VPWR
+ net666 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_37_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2956_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q _1828_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q
+ VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__o21ai_1
XFILLER_175_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1907_ _0450_ _0601_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__nor2_1
Xrebuffer128 _0185_ VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlygate4sd1_1
X_2887_ _1769_ _1770_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 sky130_fd_sc_hd__mux2_1
XFILLER_30_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4626_ net1202 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4557_ net1182 net1129 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_173_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3508_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q _0444_ VGND VGND
+ VPWR VPWR _0445_ sky130_fd_sc_hd__nand2_1
X_4488_ net1212 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_103_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3439_ _0381_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ sky130_fd_sc_hd__inv_4
X_5109_ Tile_X0Y1_E6END[6] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__buf_1
XFILLER_122_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput163 Tile_X0Y1_FrameData[28] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_2
Xinput152 Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_2
Xinput130 Tile_X0Y1_E2END[7] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
Xinput141 Tile_X0Y1_EE4END[0] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput196 Tile_X0Y1_N4END[3] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_2
Xinput185 Tile_X0Y1_N2MID[0] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_8
Xinput174 Tile_X0Y1_N1END[1] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2810_ _1719_ _1718_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 sky130_fd_sc_hd__mux2_1
X_3790_ net187 net63 net7 net117 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q VGND VGND VPWR VPWR
+ _0706_ sky130_fd_sc_hd__mux4_2
XFILLER_72_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2741_ _1660_ _1661_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2672_ net1043 net1032 net1008 net1022 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q VGND VGND VPWR VPWR
+ _1618_ sky130_fd_sc_hd__mux4_2
X_4411_ net1253 net1152 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput615 net615 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput604 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR
+ Tile_X0Y1_WW4BEG[13] sky130_fd_sc_hd__buf_6
X_4342_ net33 net1170 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4273_ net39 net1083 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3224_ _0177_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__o21ai_2
.ends

