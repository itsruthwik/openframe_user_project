module RegFile (UserCLK,
    UserCLKo,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire AD0;
 wire AD1;
 wire AD2;
 wire AD3;
 wire A_ADR0;
 wire BD0;
 wire BD1;
 wire BD2;
 wire BD3;
 wire B_ADR0;
 wire net434;
 wire net141;
 wire net403;
 wire net433;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net435;
 wire net149;
 wire net437;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net395;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net446;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire \Inst_RegFile_32x4.AD_comb[0] ;
 wire \Inst_RegFile_32x4.AD_comb[1] ;
 wire \Inst_RegFile_32x4.AD_comb[2] ;
 wire \Inst_RegFile_32x4.AD_comb[3] ;
 wire \Inst_RegFile_32x4.AD_reg[0] ;
 wire \Inst_RegFile_32x4.AD_reg[1] ;
 wire \Inst_RegFile_32x4.AD_reg[2] ;
 wire \Inst_RegFile_32x4.AD_reg[3] ;
 wire \Inst_RegFile_32x4.BD_comb[0] ;
 wire \Inst_RegFile_32x4.BD_comb[1] ;
 wire \Inst_RegFile_32x4.BD_comb[2] ;
 wire \Inst_RegFile_32x4.BD_comb[3] ;
 wire \Inst_RegFile_32x4.BD_reg[0] ;
 wire \Inst_RegFile_32x4.BD_reg[1] ;
 wire \Inst_RegFile_32x4.BD_reg[2] ;
 wire \Inst_RegFile_32x4.BD_reg[3] ;
 wire \Inst_RegFile_32x4.mem[0][0] ;
 wire \Inst_RegFile_32x4.mem[0][1] ;
 wire \Inst_RegFile_32x4.mem[0][2] ;
 wire \Inst_RegFile_32x4.mem[0][3] ;
 wire \Inst_RegFile_32x4.mem[10][0] ;
 wire \Inst_RegFile_32x4.mem[10][1] ;
 wire \Inst_RegFile_32x4.mem[10][2] ;
 wire \Inst_RegFile_32x4.mem[10][3] ;
 wire \Inst_RegFile_32x4.mem[11][0] ;
 wire \Inst_RegFile_32x4.mem[11][1] ;
 wire \Inst_RegFile_32x4.mem[11][2] ;
 wire \Inst_RegFile_32x4.mem[11][3] ;
 wire \Inst_RegFile_32x4.mem[12][0] ;
 wire \Inst_RegFile_32x4.mem[12][1] ;
 wire \Inst_RegFile_32x4.mem[12][2] ;
 wire \Inst_RegFile_32x4.mem[12][3] ;
 wire \Inst_RegFile_32x4.mem[13][0] ;
 wire \Inst_RegFile_32x4.mem[13][1] ;
 wire \Inst_RegFile_32x4.mem[13][2] ;
 wire \Inst_RegFile_32x4.mem[13][3] ;
 wire \Inst_RegFile_32x4.mem[14][0] ;
 wire \Inst_RegFile_32x4.mem[14][1] ;
 wire \Inst_RegFile_32x4.mem[14][2] ;
 wire \Inst_RegFile_32x4.mem[14][3] ;
 wire \Inst_RegFile_32x4.mem[15][0] ;
 wire \Inst_RegFile_32x4.mem[15][1] ;
 wire \Inst_RegFile_32x4.mem[15][2] ;
 wire \Inst_RegFile_32x4.mem[15][3] ;
 wire \Inst_RegFile_32x4.mem[16][0] ;
 wire \Inst_RegFile_32x4.mem[16][1] ;
 wire \Inst_RegFile_32x4.mem[16][2] ;
 wire \Inst_RegFile_32x4.mem[16][3] ;
 wire \Inst_RegFile_32x4.mem[17][0] ;
 wire \Inst_RegFile_32x4.mem[17][1] ;
 wire \Inst_RegFile_32x4.mem[17][2] ;
 wire \Inst_RegFile_32x4.mem[17][3] ;
 wire \Inst_RegFile_32x4.mem[18][0] ;
 wire \Inst_RegFile_32x4.mem[18][1] ;
 wire \Inst_RegFile_32x4.mem[18][2] ;
 wire \Inst_RegFile_32x4.mem[18][3] ;
 wire \Inst_RegFile_32x4.mem[19][0] ;
 wire \Inst_RegFile_32x4.mem[19][1] ;
 wire \Inst_RegFile_32x4.mem[19][2] ;
 wire \Inst_RegFile_32x4.mem[19][3] ;
 wire \Inst_RegFile_32x4.mem[1][0] ;
 wire \Inst_RegFile_32x4.mem[1][1] ;
 wire \Inst_RegFile_32x4.mem[1][2] ;
 wire \Inst_RegFile_32x4.mem[1][3] ;
 wire \Inst_RegFile_32x4.mem[20][0] ;
 wire \Inst_RegFile_32x4.mem[20][1] ;
 wire \Inst_RegFile_32x4.mem[20][2] ;
 wire \Inst_RegFile_32x4.mem[20][3] ;
 wire \Inst_RegFile_32x4.mem[21][0] ;
 wire \Inst_RegFile_32x4.mem[21][1] ;
 wire \Inst_RegFile_32x4.mem[21][2] ;
 wire \Inst_RegFile_32x4.mem[21][3] ;
 wire \Inst_RegFile_32x4.mem[22][0] ;
 wire \Inst_RegFile_32x4.mem[22][1] ;
 wire \Inst_RegFile_32x4.mem[22][2] ;
 wire \Inst_RegFile_32x4.mem[22][3] ;
 wire \Inst_RegFile_32x4.mem[23][0] ;
 wire \Inst_RegFile_32x4.mem[23][1] ;
 wire \Inst_RegFile_32x4.mem[23][2] ;
 wire \Inst_RegFile_32x4.mem[23][3] ;
 wire \Inst_RegFile_32x4.mem[24][0] ;
 wire \Inst_RegFile_32x4.mem[24][1] ;
 wire \Inst_RegFile_32x4.mem[24][2] ;
 wire \Inst_RegFile_32x4.mem[24][3] ;
 wire \Inst_RegFile_32x4.mem[25][0] ;
 wire \Inst_RegFile_32x4.mem[25][1] ;
 wire \Inst_RegFile_32x4.mem[25][2] ;
 wire \Inst_RegFile_32x4.mem[25][3] ;
 wire \Inst_RegFile_32x4.mem[26][0] ;
 wire \Inst_RegFile_32x4.mem[26][1] ;
 wire \Inst_RegFile_32x4.mem[26][2] ;
 wire \Inst_RegFile_32x4.mem[26][3] ;
 wire \Inst_RegFile_32x4.mem[27][0] ;
 wire \Inst_RegFile_32x4.mem[27][1] ;
 wire \Inst_RegFile_32x4.mem[27][2] ;
 wire \Inst_RegFile_32x4.mem[27][3] ;
 wire \Inst_RegFile_32x4.mem[28][0] ;
 wire \Inst_RegFile_32x4.mem[28][1] ;
 wire \Inst_RegFile_32x4.mem[28][2] ;
 wire \Inst_RegFile_32x4.mem[28][3] ;
 wire \Inst_RegFile_32x4.mem[29][0] ;
 wire \Inst_RegFile_32x4.mem[29][1] ;
 wire \Inst_RegFile_32x4.mem[29][2] ;
 wire \Inst_RegFile_32x4.mem[29][3] ;
 wire \Inst_RegFile_32x4.mem[2][0] ;
 wire \Inst_RegFile_32x4.mem[2][1] ;
 wire \Inst_RegFile_32x4.mem[2][2] ;
 wire \Inst_RegFile_32x4.mem[2][3] ;
 wire \Inst_RegFile_32x4.mem[30][0] ;
 wire \Inst_RegFile_32x4.mem[30][1] ;
 wire \Inst_RegFile_32x4.mem[30][2] ;
 wire \Inst_RegFile_32x4.mem[30][3] ;
 wire \Inst_RegFile_32x4.mem[31][0] ;
 wire \Inst_RegFile_32x4.mem[31][1] ;
 wire \Inst_RegFile_32x4.mem[31][2] ;
 wire \Inst_RegFile_32x4.mem[31][3] ;
 wire \Inst_RegFile_32x4.mem[3][0] ;
 wire \Inst_RegFile_32x4.mem[3][1] ;
 wire \Inst_RegFile_32x4.mem[3][2] ;
 wire \Inst_RegFile_32x4.mem[3][3] ;
 wire \Inst_RegFile_32x4.mem[4][0] ;
 wire \Inst_RegFile_32x4.mem[4][1] ;
 wire \Inst_RegFile_32x4.mem[4][2] ;
 wire \Inst_RegFile_32x4.mem[4][3] ;
 wire \Inst_RegFile_32x4.mem[5][0] ;
 wire \Inst_RegFile_32x4.mem[5][1] ;
 wire \Inst_RegFile_32x4.mem[5][2] ;
 wire \Inst_RegFile_32x4.mem[5][3] ;
 wire \Inst_RegFile_32x4.mem[6][0] ;
 wire \Inst_RegFile_32x4.mem[6][1] ;
 wire \Inst_RegFile_32x4.mem[6][2] ;
 wire \Inst_RegFile_32x4.mem[6][3] ;
 wire \Inst_RegFile_32x4.mem[7][0] ;
 wire \Inst_RegFile_32x4.mem[7][1] ;
 wire \Inst_RegFile_32x4.mem[7][2] ;
 wire \Inst_RegFile_32x4.mem[7][3] ;
 wire \Inst_RegFile_32x4.mem[8][0] ;
 wire \Inst_RegFile_32x4.mem[8][1] ;
 wire \Inst_RegFile_32x4.mem[8][2] ;
 wire \Inst_RegFile_32x4.mem[8][3] ;
 wire \Inst_RegFile_32x4.mem[9][0] ;
 wire \Inst_RegFile_32x4.mem[9][1] ;
 wire \Inst_RegFile_32x4.mem[9][2] ;
 wire \Inst_RegFile_32x4.mem[9][3] ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_RegFile_switch_matrix.E1BEG0 ;
 wire \Inst_RegFile_switch_matrix.E1BEG1 ;
 wire \Inst_RegFile_switch_matrix.E1BEG2 ;
 wire \Inst_RegFile_switch_matrix.E1BEG3 ;
 wire \Inst_RegFile_switch_matrix.E2BEG0 ;
 wire \Inst_RegFile_switch_matrix.E2BEG1 ;
 wire \Inst_RegFile_switch_matrix.E2BEG2 ;
 wire \Inst_RegFile_switch_matrix.E2BEG3 ;
 wire \Inst_RegFile_switch_matrix.E2BEG4 ;
 wire \Inst_RegFile_switch_matrix.E2BEG5 ;
 wire \Inst_RegFile_switch_matrix.E2BEG6 ;
 wire \Inst_RegFile_switch_matrix.E2BEG7 ;
 wire \Inst_RegFile_switch_matrix.E6BEG0 ;
 wire \Inst_RegFile_switch_matrix.E6BEG1 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG0 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG1 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG2 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG3 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG7 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG7 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG7 ;
 wire \Inst_RegFile_switch_matrix.N1BEG0 ;
 wire \Inst_RegFile_switch_matrix.N1BEG1 ;
 wire \Inst_RegFile_switch_matrix.N1BEG2 ;
 wire \Inst_RegFile_switch_matrix.N1BEG3 ;
 wire \Inst_RegFile_switch_matrix.N4BEG0 ;
 wire \Inst_RegFile_switch_matrix.N4BEG1 ;
 wire \Inst_RegFile_switch_matrix.N4BEG2 ;
 wire \Inst_RegFile_switch_matrix.N4BEG3 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG0 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG1 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG2 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG3 ;
 wire \Inst_RegFile_switch_matrix.S1BEG0 ;
 wire \Inst_RegFile_switch_matrix.S1BEG1 ;
 wire \Inst_RegFile_switch_matrix.S1BEG2 ;
 wire \Inst_RegFile_switch_matrix.S1BEG3 ;
 wire \Inst_RegFile_switch_matrix.S4BEG0 ;
 wire \Inst_RegFile_switch_matrix.S4BEG1 ;
 wire \Inst_RegFile_switch_matrix.S4BEG2 ;
 wire \Inst_RegFile_switch_matrix.S4BEG3 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG0 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG1 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG2 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG3 ;
 wire \Inst_RegFile_switch_matrix.W1BEG0 ;
 wire \Inst_RegFile_switch_matrix.W1BEG1 ;
 wire \Inst_RegFile_switch_matrix.W1BEG2 ;
 wire \Inst_RegFile_switch_matrix.W1BEG3 ;
 wire \Inst_RegFile_switch_matrix.W6BEG0 ;
 wire \Inst_RegFile_switch_matrix.W6BEG1 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG0 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG1 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG2 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG3 ;
 wire net240;
 wire net241;
 wire net242;
 wire net432;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net444;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net456;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net454;
 wire net447;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net428;
 wire net402;
 wire net427;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net452;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net453;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net431;
 wire net397;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net436;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net439;
 wire net445;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net455;
 wire net394;
 wire net382;
 wire net398;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net393;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_4_0_0_UserCLK_regs;
 wire clknet_4_1_0_UserCLK_regs;
 wire clknet_4_2_0_UserCLK_regs;
 wire clknet_4_3_0_UserCLK_regs;
 wire clknet_4_4_0_UserCLK_regs;
 wire clknet_4_5_0_UserCLK_regs;
 wire clknet_4_6_0_UserCLK_regs;
 wire clknet_4_7_0_UserCLK_regs;
 wire clknet_4_8_0_UserCLK_regs;
 wire clknet_4_9_0_UserCLK_regs;
 wire clknet_4_10_0_UserCLK_regs;
 wire clknet_4_11_0_UserCLK_regs;
 wire clknet_4_12_0_UserCLK_regs;
 wire clknet_4_13_0_UserCLK_regs;
 wire clknet_4_14_0_UserCLK_regs;
 wire clknet_4_15_0_UserCLK_regs;
 wire net396;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;

 sky130_fd_sc_hd__inv_1 _1074_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0968_));
 sky130_fd_sc_hd__inv_1 _1075_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ),
    .Y(_0969_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(net72),
    .Y(_0970_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .Y(_0971_));
 sky130_fd_sc_hd__inv_1 _1078_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .Y(_0972_));
 sky130_fd_sc_hd__inv_2 _1079_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ),
    .Y(_0973_));
 sky130_fd_sc_hd__inv_1 _1080_ (.A(net128),
    .Y(_0974_));
 sky130_fd_sc_hd__inv_2 _1081_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ),
    .Y(_0975_));
 sky130_fd_sc_hd__inv_2 _1082_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_0976_));
 sky130_fd_sc_hd__inv_1 _1083_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ),
    .Y(_0977_));
 sky130_fd_sc_hd__inv_2 _1084_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ),
    .Y(_0978_));
 sky130_fd_sc_hd__inv_1 _1085_ (.A(net17),
    .Y(_0979_));
 sky130_fd_sc_hd__inv_1 _1086_ (.A(net102),
    .Y(_0980_));
 sky130_fd_sc_hd__inv_1 _1087_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .Y(_0981_));
 sky130_fd_sc_hd__inv_1 _1088_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ),
    .Y(_0982_));
 sky130_fd_sc_hd__inv_2 _1089_ (.A(net130),
    .Y(_0983_));
 sky130_fd_sc_hd__inv_1 _1090_ (.A(net139),
    .Y(_0984_));
 sky130_fd_sc_hd__inv_2 _1091_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ),
    .Y(_0985_));
 sky130_fd_sc_hd__inv_2 _1092_ (.A(net13),
    .Y(_0986_));
 sky130_fd_sc_hd__inv_1 _1093_ (.A(net126),
    .Y(_0987_));
 sky130_fd_sc_hd__inv_1 _1094_ (.A(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ),
    .Y(_0988_));
 sky130_fd_sc_hd__inv_2 _1095_ (.A(net15),
    .Y(_0989_));
 sky130_fd_sc_hd__inv_1 _1096_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .Y(_0990_));
 sky130_fd_sc_hd__inv_1 _1097_ (.A(net691),
    .Y(_0991_));
 sky130_fd_sc_hd__inv_2 _1098_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ),
    .Y(_0992_));
 sky130_fd_sc_hd__inv_1 _1099_ (.A(\Inst_RegFile_32x4.mem[10][1] ),
    .Y(_0993_));
 sky130_fd_sc_hd__inv_2 _1100_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ),
    .Y(_0994_));
 sky130_fd_sc_hd__inv_2 _1101_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ),
    .Y(_0995_));
 sky130_fd_sc_hd__inv_2 _1102_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ),
    .Y(_0996_));
 sky130_fd_sc_hd__inv_2 _1103_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .Y(_0997_));
 sky130_fd_sc_hd__inv_2 _1104_ (.A(net74),
    .Y(_0998_));
 sky130_fd_sc_hd__inv_1 _1105_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .Y(_0999_));
 sky130_fd_sc_hd__inv_2 _1106_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ),
    .Y(_1000_));
 sky130_fd_sc_hd__inv_1 _1107_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .Y(_1001_));
 sky130_fd_sc_hd__inv_1 _1108_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ),
    .Y(_1002_));
 sky130_fd_sc_hd__inv_1 _1109_ (.A(net98),
    .Y(_1003_));
 sky130_fd_sc_hd__inv_1 _1110_ (.A(\Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ),
    .Y(_1004_));
 sky130_fd_sc_hd__inv_2 _1111_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ),
    .Y(_1005_));
 sky130_fd_sc_hd__inv_2 _1112_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_1006_));
 sky130_fd_sc_hd__inv_1 _1113_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(_1007_));
 sky130_fd_sc_hd__inv_1 _1114_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ),
    .Y(_1008_));
 sky130_fd_sc_hd__inv_2 _1115_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_1009_));
 sky130_fd_sc_hd__inv_2 _1116_ (.A(net1),
    .Y(_1010_));
 sky130_fd_sc_hd__inv_1 _1117_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .Y(_1011_));
 sky130_fd_sc_hd__inv_1 _1118_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ),
    .Y(_1012_));
 sky130_fd_sc_hd__inv_2 _1119_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ),
    .Y(_1013_));
 sky130_fd_sc_hd__inv_1 _1120_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ),
    .Y(_1014_));
 sky130_fd_sc_hd__inv_1 _1121_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_1015_));
 sky130_fd_sc_hd__inv_1 _1122_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ),
    .Y(_1016_));
 sky130_fd_sc_hd__inv_2 _1123_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .Y(_1017_));
 sky130_fd_sc_hd__inv_1 _1124_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ),
    .Y(_1018_));
 sky130_fd_sc_hd__inv_1 _1125_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .Y(_1019_));
 sky130_fd_sc_hd__inv_1 _1126_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ),
    .Y(_1020_));
 sky130_fd_sc_hd__inv_1 _1127_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ),
    .Y(_1021_));
 sky130_fd_sc_hd__inv_2 _1128_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .Y(_1022_));
 sky130_fd_sc_hd__inv_1 _1129_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ),
    .Y(_1023_));
 sky130_fd_sc_hd__inv_1 _1130_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ),
    .Y(_1024_));
 sky130_fd_sc_hd__inv_1 _1131_ (.A(\Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ),
    .Y(_1025_));
 sky130_fd_sc_hd__inv_1 _1132_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .Y(_1026_));
 sky130_fd_sc_hd__inv_2 _1133_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ),
    .Y(_1027_));
 sky130_fd_sc_hd__inv_2 _1134_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .Y(_1028_));
 sky130_fd_sc_hd__inv_2 _1135_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .Y(_1029_));
 sky130_fd_sc_hd__inv_2 _1136_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_1030_));
 sky130_fd_sc_hd__inv_2 _1137_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ),
    .Y(_1031_));
 sky130_fd_sc_hd__mux4_2 _1138_ (.A0(net650),
    .A1(net684),
    .A2(net398),
    .A3(net404),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1032_));
 sky130_fd_sc_hd__or2_4 _1139_ (.A(_1032_),
    .B(_0995_),
    .X(_1033_));
 sky130_fd_sc_hd__mux4_1 _1140_ (.A0(net116),
    .A1(net674),
    .A2(net660),
    .A3(net413),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1034_));
 sky130_fd_sc_hd__o21a_1 _1141_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_1034_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_1035_));
 sky130_fd_sc_hd__mux4_1 _1142_ (.A0(net25),
    .A1(net86),
    .A2(net88),
    .A3(net96),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1036_));
 sky130_fd_sc_hd__mux4_1 _1143_ (.A0(net60),
    .A1(net68),
    .A2(net784),
    .A3(net11),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _1144_ (.A0(_1036_),
    .A1(_1037_),
    .S(_0995_),
    .X(_1038_));
 sky130_fd_sc_hd__a22o_1 _1145_ (.A1(_1033_),
    .A2(_1035_),
    .B1(_1038_),
    .B2(_0996_),
    .X(\Inst_RegFile_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__a221o_2 _1146_ (.A1(_1033_),
    .A2(_1035_),
    .B1(_1038_),
    .B2(_0996_),
    .C1(_0994_),
    .X(_1039_));
 sky130_fd_sc_hd__o21a_1 _1147_ (.A1(net100),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _1148_ (.A0(_0970_),
    .A1(_0989_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_1041_));
 sky130_fd_sc_hd__nor2_1 _1149_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__a211o_1 _1150_ (.A1(_1039_),
    .A2(_1040_),
    .B1(_1042_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_1043_));
 sky130_fd_sc_hd__mux4_2 _1151_ (.A0(net73),
    .A1(net16),
    .A2(net101),
    .A3(net129),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_1044_));
 sky130_fd_sc_hd__clkinv_2 _1152_ (.A(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a21oi_1 _1153_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_1045_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ),
    .Y(_1046_));
 sky130_fd_sc_hd__mux4_2 _1154_ (.A0(net691),
    .A1(net671),
    .A2(net657),
    .A3(net652),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1047_));
 sky130_fd_sc_hd__or2_4 _1155_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .B(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__mux4_1 _1156_ (.A0(net681),
    .A1(net634),
    .A2(net406),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .X(_1049_));
 sky130_fd_sc_hd__o21a_1 _1157_ (.A1(_0990_),
    .A2(_1049_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_1050_));
 sky130_fd_sc_hd__mux4_1 _1158_ (.A0(net60),
    .A1(net66),
    .A2(net78),
    .A3(net9),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1051_));
 sky130_fd_sc_hd__mux4_1 _1159_ (.A0(net782),
    .A1(net94),
    .A2(net113),
    .A3(net122),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _1160_ (.A0(_1051_),
    .A1(_1052_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .X(_1053_));
 sky130_fd_sc_hd__a22o_4 _1161_ (.A1(_1050_),
    .A2(_1048_),
    .B1(_1053_),
    .B2(_0992_),
    .X(\Inst_RegFile_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__a221o_1 _1162_ (.A1(_1048_),
    .A2(_1050_),
    .B1(_1053_),
    .B2(_0992_),
    .C1(_0997_),
    .X(_1054_));
 sky130_fd_sc_hd__or2_1 _1163_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .B(net108),
    .X(_1055_));
 sky130_fd_sc_hd__mux2_1 _1164_ (.A0(net84),
    .A1(net7),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1056_));
 sky130_fd_sc_hd__inv_1 _1165_ (.A(_1056_),
    .Y(_1057_));
 sky130_fd_sc_hd__o21ai_1 _1166_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_1057_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .Y(_1058_));
 sky130_fd_sc_hd__a31o_1 _1167_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_1054_),
    .A3(_1055_),
    .B1(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__mux4_2 _1168_ (.A0(net65),
    .A1(net8),
    .A2(net93),
    .A3(net137),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_1060_));
 sky130_fd_sc_hd__o21a_1 _1169_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_1060_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ),
    .X(_1061_));
 sky130_fd_sc_hd__a22oi_2 _1170_ (.A1(_1043_),
    .A2(_1046_),
    .B1(_1059_),
    .B2(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__mux2_1 _1171_ (.A0(\Inst_RegFile_32x4.mem[8][0] ),
    .A1(\Inst_RegFile_32x4.mem[9][0] ),
    .S(net616),
    .X(_1063_));
 sky130_fd_sc_hd__mux4_1 _1172_ (.A0(net693),
    .A1(net672),
    .A2(net658),
    .A3(net419),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1064_));
 sky130_fd_sc_hd__or2_1 _1173_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .B(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__mux4_2 _1174_ (.A0(net649),
    .A1(net683),
    .A2(net428),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1066_));
 sky130_fd_sc_hd__o21a_1 _1175_ (.A1(_1066_),
    .A2(_0999_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_1067_));
 sky130_fd_sc_hd__mux4_1 _1176_ (.A0(net60),
    .A1(net68),
    .A2(net784),
    .A3(net11),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1068_));
 sky130_fd_sc_hd__mux4_1 _1177_ (.A0(net88),
    .A1(net96),
    .A2(net112),
    .A3(net114),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_1 _1178_ (.A0(_1068_),
    .A1(_1069_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_1070_));
 sky130_fd_sc_hd__a22oi_4 _1179_ (.A1(_1067_),
    .A2(_1065_),
    .B1(_1070_),
    .B2(_1000_),
    .Y(_1071_));
 sky130_fd_sc_hd__inv_6 _1180_ (.A(net436),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _1181_ (.A0(_0998_),
    .A1(_0983_),
    .A2(_0980_),
    .A3(_1071_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1072_));
 sky130_fd_sc_hd__inv_2 _1182_ (.A(net433),
    .Y(_1073_));
 sky130_fd_sc_hd__mux4_2 _1183_ (.A0(net75),
    .A1(net18),
    .A2(net103),
    .A3(net131),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ),
    .X(_0128_));
 sky130_fd_sc_hd__nand2_1 _1184_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ),
    .B(_0128_),
    .Y(_0129_));
 sky130_fd_sc_hd__o21ai_1 _1185_ (.A1(_1072_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ),
    .B1(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__mux4_2 _1186_ (.A0(net691),
    .A1(net671),
    .A2(net657),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0131_));
 sky130_fd_sc_hd__or2_4 _1187_ (.A(_0131_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0132_));
 sky130_fd_sc_hd__mux4_2 _1188_ (.A0(net681),
    .A1(net634),
    .A2(net406),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0133_));
 sky130_fd_sc_hd__o21a_1 _1189_ (.A1(_0133_),
    .A2(_1001_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0134_));
 sky130_fd_sc_hd__mux4_1 _1190_ (.A0(net66),
    .A1(net9),
    .A2(net784),
    .A3(net26),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0135_));
 sky130_fd_sc_hd__mux4_1 _1191_ (.A0(net21),
    .A1(net94),
    .A2(net106),
    .A3(net122),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _1192_ (.A0(_0135_),
    .A1(_0136_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_4 _1193_ (.A1(_0132_),
    .A2(_0134_),
    .B1(_0137_),
    .B2(_1002_),
    .X(\Inst_RegFile_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__inv_1 _1194_ (.A(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .Y(_0138_));
 sky130_fd_sc_hd__mux4_2 _1195_ (.A0(net79),
    .A1(net122),
    .A2(net111),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_0139_));
 sky130_fd_sc_hd__mux4_2 _1196_ (.A0(net67),
    .A1(net10),
    .A2(net111),
    .A3(net123),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_4 _1197_ (.A0(_0140_),
    .A1(_0139_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_4 _1198_ (.A0(_0130_),
    .A1(_0141_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _1199_ (.A0(\Inst_RegFile_32x4.mem[10][0] ),
    .A1(\Inst_RegFile_32x4.mem[11][0] ),
    .S(net616),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _1200_ (.A0(_0143_),
    .A1(_1063_),
    .S(net444),
    .X(_0144_));
 sky130_fd_sc_hd__nand2b_1 _1201_ (.A_N(net416),
    .B(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__mux4_2 _1202_ (.A0(net691),
    .A1(net414),
    .A2(net415),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0146_));
 sky130_fd_sc_hd__mux4_2 _1203_ (.A0(net681),
    .A1(net634),
    .A2(net406),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_4 _1204_ (.A0(_0146_),
    .A1(_0147_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .X(_0148_));
 sky130_fd_sc_hd__mux4_1 _1205_ (.A0(net60),
    .A1(net66),
    .A2(net85),
    .A3(net9),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0149_));
 sky130_fd_sc_hd__mux4_1 _1206_ (.A0(net21),
    .A1(net94),
    .A2(net106),
    .A3(net122),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _1207_ (.A0(_0149_),
    .A1(_0150_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_4 _1208_ (.A0(_0151_),
    .A1(_0148_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Inst_RegFile_switch_matrix.JW2BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1209_ (.A0(net26),
    .A1(net137),
    .A2(net106),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_0152_));
 sky130_fd_sc_hd__mux4_2 _1210_ (.A0(net84),
    .A1(net6),
    .A2(net91),
    .A3(net119),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_4 _1211_ (.A0(_0153_),
    .A1(_0152_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_0154_));
 sky130_fd_sc_hd__mux4_1 _1212_ (.A0(net138),
    .A1(net673),
    .A2(net659),
    .A3(net413),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0155_));
 sky130_fd_sc_hd__nand2b_1 _1213_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .B(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__mux4_2 _1214_ (.A0(net649),
    .A1(net683),
    .A2(net637),
    .A3(net447),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0157_));
 sky130_fd_sc_hd__a21boi_2 _1215_ (.A1(_0157_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ),
    .Y(_0158_));
 sky130_fd_sc_hd__mux4_1 _1216_ (.A0(net60),
    .A1(net68),
    .A2(net784),
    .A3(net11),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0159_));
 sky130_fd_sc_hd__mux4_1 _1217_ (.A0(net86),
    .A1(net96),
    .A2(net88),
    .A3(net693),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _1218_ (.A0(_0159_),
    .A1(_0160_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_0161_));
 sky130_fd_sc_hd__a2bb2o_4 _1219_ (.A1_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ),
    .A2_N(_0161_),
    .B1(_0158_),
    .B2(_0156_),
    .X(_0162_));
 sky130_fd_sc_hd__inv_2 _1220_ (.A(_0162_),
    .Y(\Inst_RegFile_switch_matrix.JW2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _1221_ (.A0(_0986_),
    .A1(_0987_),
    .A2(_1003_),
    .A3(_0162_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _1222_ (.A0(net71),
    .A1(net14),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _1223_ (.A0(net99),
    .A1(net127),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_0165_));
 sky130_fd_sc_hd__o21a_1 _1224_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ),
    .A2(_0164_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_0166_));
 sky130_fd_sc_hd__o21ai_1 _1225_ (.A1(_1004_),
    .A2(_0165_),
    .B1(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__o21a_1 _1226_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_0163_),
    .B1(_1005_),
    .X(_0168_));
 sky130_fd_sc_hd__a2bb2o_4 _1227_ (.A1_N(_1005_),
    .A2_N(_0154_),
    .B1(_0167_),
    .B2(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _1228_ (.A0(\Inst_RegFile_32x4.mem[12][0] ),
    .A1(\Inst_RegFile_32x4.mem[13][0] ),
    .S(net394),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _1229_ (.A0(\Inst_RegFile_32x4.mem[14][0] ),
    .A1(\Inst_RegFile_32x4.mem[15][0] ),
    .S(net395),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _1230_ (.A0(_0171_),
    .A1(_0170_),
    .S(net445),
    .X(_0172_));
 sky130_fd_sc_hd__a21oi_1 _1231_ (.A1(net416),
    .A2(_0172_),
    .B1(net393),
    .Y(_0173_));
 sky130_fd_sc_hd__mux2_1 _1232_ (.A0(\Inst_RegFile_32x4.mem[0][0] ),
    .A1(\Inst_RegFile_32x4.mem[1][0] ),
    .S(net615),
    .X(_0174_));
 sky130_fd_sc_hd__and2b_1 _1233_ (.A_N(_0174_),
    .B(net446),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _1234_ (.A0(\Inst_RegFile_32x4.mem[2][0] ),
    .A1(\Inst_RegFile_32x4.mem[3][0] ),
    .S(net615),
    .X(_0176_));
 sky130_fd_sc_hd__nor2_1 _1235_ (.A(net445),
    .B(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__mux2_1 _1236_ (.A0(\Inst_RegFile_32x4.mem[4][0] ),
    .A1(\Inst_RegFile_32x4.mem[5][0] ),
    .S(net394),
    .X(_0178_));
 sky130_fd_sc_hd__nand2b_1 _1237_ (.A_N(_0178_),
    .B(net445),
    .Y(_0179_));
 sky130_fd_sc_hd__mux2_1 _1238_ (.A0(\Inst_RegFile_32x4.mem[6][0] ),
    .A1(\Inst_RegFile_32x4.mem[7][0] ),
    .S(net394),
    .X(_0180_));
 sky130_fd_sc_hd__o211ai_1 _1239_ (.A1(net445),
    .A2(_0180_),
    .B1(_0179_),
    .C1(net416),
    .Y(_0181_));
 sky130_fd_sc_hd__o311a_1 _1240_ (.A1(net416),
    .A2(_0175_),
    .A3(_0177_),
    .B1(_0181_),
    .C1(net393),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _1241_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .B(_0162_),
    .Y(_0183_));
 sky130_fd_sc_hd__o21a_1 _1242_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ),
    .X(_0184_));
 sky130_fd_sc_hd__mux4_1 _1243_ (.A0(net693),
    .A1(net674),
    .A2(net660),
    .A3(net656),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0185_));
 sky130_fd_sc_hd__mux4_2 _1244_ (.A0(net405),
    .A1(BD0),
    .A2(BD2),
    .A3(net412),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_4 _1245_ (.A0(_0185_),
    .A1(_0186_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0187_));
 sky130_fd_sc_hd__mux4_1 _1246_ (.A0(net11),
    .A1(net88),
    .A2(net96),
    .A3(net114),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0188_));
 sky130_fd_sc_hd__mux4_1 _1247_ (.A0(net60),
    .A1(net84),
    .A2(net68),
    .A3(net784),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _1248_ (.A0(_0189_),
    .A1(_0188_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_4 _1249_ (.A0(_0190_),
    .A1(_0187_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ),
    .X(\Inst_RegFile_switch_matrix.JN2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _1250_ (.A0(net62),
    .A1(net90),
    .A2(net24),
    .A3(net118),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_4 _1251_ (.A0(_0191_),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0192_));
 sky130_fd_sc_hd__a22o_1 _1252_ (.A1(_0183_),
    .A2(_0184_),
    .B1(_1006_),
    .B2(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__mux4_1 _1253_ (.A0(net117),
    .A1(net674),
    .A2(net660),
    .A3(net656),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0194_));
 sky130_fd_sc_hd__or2_4 _1254_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__mux4_2 _1255_ (.A0(net405),
    .A1(net684),
    .A2(net668),
    .A3(net404),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0196_));
 sky130_fd_sc_hd__o21a_1 _1256_ (.A1(_0972_),
    .A2(_0196_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ),
    .X(_0197_));
 sky130_fd_sc_hd__mux4_1 _1257_ (.A0(net61),
    .A1(net69),
    .A2(net783),
    .A3(net12),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0198_));
 sky130_fd_sc_hd__mux4_1 _1258_ (.A0(net24),
    .A1(net87),
    .A2(net89),
    .A3(net97),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _1259_ (.A0(_0198_),
    .A1(_0199_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_4 _1260_ (.A1(_0195_),
    .A2(_0197_),
    .B1(_0200_),
    .B2(_0973_),
    .X(\Inst_RegFile_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__a221o_1 _1261_ (.A1(_0195_),
    .A2(_0197_),
    .B1(_0200_),
    .B2(_0973_),
    .C1(_0971_),
    .X(_0201_));
 sky130_fd_sc_hd__o21a_1 _1262_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .A2(net128),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _1263_ (.A0(net72),
    .A1(net100),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_0203_));
 sky130_fd_sc_hd__a22o_1 _1264_ (.A1(_0201_),
    .A2(_0202_),
    .B1(_0203_),
    .B2(_0975_),
    .X(_0204_));
 sky130_fd_sc_hd__mux4_1 _1265_ (.A0(net75),
    .A1(net18),
    .A2(net103),
    .A3(net131),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _1266_ (.A0(_0204_),
    .A1(_0205_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _1267_ (.A0(net63),
    .A1(net91),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _1268_ (.A0(_0206_),
    .A1(_0207_),
    .S(_1006_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_4 _1269_ (.A0(_0208_),
    .A1(_0193_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0209_));
 sky130_fd_sc_hd__a21o_1 _1270_ (.A1(_0145_),
    .A2(_0173_),
    .B1(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _1271_ (.A0(\Inst_RegFile_32x4.mem[26][0] ),
    .A1(\Inst_RegFile_32x4.mem[27][0] ),
    .S(net619),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _1272_ (.A0(\Inst_RegFile_32x4.mem[24][0] ),
    .A1(\Inst_RegFile_32x4.mem[25][0] ),
    .S(net619),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _1273_ (.A0(_0211_),
    .A1(_0212_),
    .S(net678),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _1274_ (.A0(\Inst_RegFile_32x4.mem[30][0] ),
    .A1(\Inst_RegFile_32x4.mem[31][0] ),
    .S(net615),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _1275_ (.A0(\Inst_RegFile_32x4.mem[28][0] ),
    .A1(\Inst_RegFile_32x4.mem[29][0] ),
    .S(net615),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _1276_ (.A0(_0214_),
    .A1(_0215_),
    .S(net446),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _1277_ (.A0(_0213_),
    .A1(_0216_),
    .S(net663),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _1278_ (.A0(\Inst_RegFile_32x4.mem[16][0] ),
    .A1(\Inst_RegFile_32x4.mem[17][0] ),
    .S(net618),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _1279_ (.A0(\Inst_RegFile_32x4.mem[18][0] ),
    .A1(\Inst_RegFile_32x4.mem[19][0] ),
    .S(net618),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _1280_ (.A0(_0219_),
    .A1(_0218_),
    .S(net679),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _1281_ (.A0(\Inst_RegFile_32x4.mem[22][0] ),
    .A1(\Inst_RegFile_32x4.mem[23][0] ),
    .S(net617),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _1282_ (.A0(\Inst_RegFile_32x4.mem[20][0] ),
    .A1(\Inst_RegFile_32x4.mem[21][0] ),
    .S(net617),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _1283_ (.A0(_0221_),
    .A1(_0222_),
    .S(net678),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _1284_ (.A0(_0220_),
    .A1(_0223_),
    .S(net664),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _1285_ (.A0(_0217_),
    .A1(_0224_),
    .S(_0169_),
    .X(_0225_));
 sky130_fd_sc_hd__a2bb2o_4 _1286_ (.A1_N(_0182_),
    .A2_N(_0210_),
    .B1(_0209_),
    .B2(_0225_),
    .X(\Inst_RegFile_32x4.AD_comb[0] ));
 sky130_fd_sc_hd__mux2_4 _1287_ (.A0(\Inst_RegFile_32x4.AD_comb[0] ),
    .A1(\Inst_RegFile_32x4.AD_reg[0] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD0));
 sky130_fd_sc_hd__mux2_1 _1288_ (.A0(\Inst_RegFile_32x4.mem[10][1] ),
    .A1(\Inst_RegFile_32x4.mem[11][1] ),
    .S(net614),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _1289_ (.A0(\Inst_RegFile_32x4.mem[8][1] ),
    .A1(\Inst_RegFile_32x4.mem[9][1] ),
    .S(net614),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _1290_ (.A0(_0226_),
    .A1(_0227_),
    .S(net444),
    .X(_0228_));
 sky130_fd_sc_hd__and2b_1 _1291_ (.A_N(net416),
    .B(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _1292_ (.A0(\Inst_RegFile_32x4.mem[14][1] ),
    .A1(\Inst_RegFile_32x4.mem[15][1] ),
    .S(A_ADR0),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _1293_ (.A0(\Inst_RegFile_32x4.mem[12][1] ),
    .A1(\Inst_RegFile_32x4.mem[13][1] ),
    .S(net612),
    .X(_0231_));
 sky130_fd_sc_hd__nand2b_1 _1294_ (.A_N(_0231_),
    .B(net445),
    .Y(_0232_));
 sky130_fd_sc_hd__o211a_1 _1295_ (.A1(net446),
    .A2(_0230_),
    .B1(_0232_),
    .C1(net662),
    .X(_0233_));
 sky130_fd_sc_hd__nor3_2 _1296_ (.A(_0233_),
    .B(_0229_),
    .C(net651),
    .Y(_0234_));
 sky130_fd_sc_hd__mux2_1 _1297_ (.A0(\Inst_RegFile_32x4.mem[0][1] ),
    .A1(\Inst_RegFile_32x4.mem[1][1] ),
    .S(net616),
    .X(_0235_));
 sky130_fd_sc_hd__inv_2 _1298_ (.A(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__mux2_1 _1299_ (.A0(\Inst_RegFile_32x4.mem[2][1] ),
    .A1(\Inst_RegFile_32x4.mem[3][1] ),
    .S(net614),
    .X(_0237_));
 sky130_fd_sc_hd__nor2_1 _1300_ (.A(net444),
    .B(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__a211o_1 _1301_ (.A1(net444),
    .A2(_0236_),
    .B1(_0238_),
    .C1(net662),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_4 _1302_ (.A0(\Inst_RegFile_32x4.mem[4][1] ),
    .A1(\Inst_RegFile_32x4.mem[5][1] ),
    .S(net394),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_2 _1303_ (.A0(\Inst_RegFile_32x4.mem[6][1] ),
    .A1(\Inst_RegFile_32x4.mem[7][1] ),
    .S(net394),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_4 _1304_ (.A0(_0241_),
    .A1(_0240_),
    .S(net675),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _1305_ (.A(net662),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__a31o_1 _1306_ (.A1(net393),
    .A2(_0239_),
    .A3(_0243_),
    .B1(_0209_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _1307_ (.A0(\Inst_RegFile_32x4.mem[26][1] ),
    .A1(\Inst_RegFile_32x4.mem[27][1] ),
    .S(net619),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _1308_ (.A0(\Inst_RegFile_32x4.mem[24][1] ),
    .A1(\Inst_RegFile_32x4.mem[25][1] ),
    .S(net619),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _1309_ (.A0(_0245_),
    .A1(_0246_),
    .S(net678),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _1310_ (.A0(\Inst_RegFile_32x4.mem[30][1] ),
    .A1(\Inst_RegFile_32x4.mem[31][1] ),
    .S(net615),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _1311_ (.A0(\Inst_RegFile_32x4.mem[28][1] ),
    .A1(\Inst_RegFile_32x4.mem[29][1] ),
    .S(net615),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _1312_ (.A0(_0248_),
    .A1(_0249_),
    .S(net446),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _1313_ (.A0(_0247_),
    .A1(_0250_),
    .S(net664),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _1314_ (.A0(\Inst_RegFile_32x4.mem[16][1] ),
    .A1(\Inst_RegFile_32x4.mem[17][1] ),
    .S(net618),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _1315_ (.A0(\Inst_RegFile_32x4.mem[18][1] ),
    .A1(\Inst_RegFile_32x4.mem[19][1] ),
    .S(net618),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _1316_ (.A0(_0253_),
    .A1(_0252_),
    .S(net678),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _1317_ (.A0(\Inst_RegFile_32x4.mem[22][1] ),
    .A1(\Inst_RegFile_32x4.mem[23][1] ),
    .S(net617),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _1318_ (.A0(\Inst_RegFile_32x4.mem[20][1] ),
    .A1(\Inst_RegFile_32x4.mem[21][1] ),
    .S(net617),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _1319_ (.A0(_0255_),
    .A1(_0256_),
    .S(net678),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _1320_ (.A0(_0254_),
    .A1(_0257_),
    .S(net664),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _1321_ (.A0(_0251_),
    .A1(_0258_),
    .S(net393),
    .X(_0259_));
 sky130_fd_sc_hd__a2bb2o_4 _1322_ (.A1_N(_0244_),
    .A2_N(_0234_),
    .B1(_0259_),
    .B2(_0209_),
    .X(\Inst_RegFile_32x4.AD_comb[1] ));
 sky130_fd_sc_hd__mux2_4 _1323_ (.A0(\Inst_RegFile_32x4.AD_comb[1] ),
    .A1(\Inst_RegFile_32x4.AD_reg[1] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD1));
 sky130_fd_sc_hd__mux2_1 _1324_ (.A0(\Inst_RegFile_32x4.mem[10][2] ),
    .A1(\Inst_RegFile_32x4.mem[11][2] ),
    .S(net616),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _1325_ (.A0(\Inst_RegFile_32x4.mem[8][2] ),
    .A1(\Inst_RegFile_32x4.mem[9][2] ),
    .S(net614),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_4 _1326_ (.A0(_0260_),
    .A1(_0261_),
    .S(net444),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _1327_ (.A0(\Inst_RegFile_32x4.mem[12][2] ),
    .A1(\Inst_RegFile_32x4.mem[13][2] ),
    .S(net614),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _1328_ (.A0(\Inst_RegFile_32x4.mem[14][2] ),
    .A1(\Inst_RegFile_32x4.mem[15][2] ),
    .S(net614),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_4 _1329_ (.A0(_0264_),
    .A1(_0263_),
    .S(net676),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_4 _1330_ (.A0(_0262_),
    .A1(_0265_),
    .S(net663),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _1331_ (.A0(\Inst_RegFile_32x4.mem[2][2] ),
    .A1(\Inst_RegFile_32x4.mem[3][2] ),
    .S(net614),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _1332_ (.A0(\Inst_RegFile_32x4.mem[0][2] ),
    .A1(\Inst_RegFile_32x4.mem[1][2] ),
    .S(net614),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_2 _1333_ (.A0(_0267_),
    .A1(_0268_),
    .S(net676),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _1334_ (.A0(\Inst_RegFile_32x4.mem[6][2] ),
    .A1(\Inst_RegFile_32x4.mem[7][2] ),
    .S(net612),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _1335_ (.A0(\Inst_RegFile_32x4.mem[4][2] ),
    .A1(\Inst_RegFile_32x4.mem[5][2] ),
    .S(net612),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_2 _1336_ (.A0(_0270_),
    .A1(_0271_),
    .S(net675),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_4 _1337_ (.A0(_0269_),
    .A1(_0272_),
    .S(net662),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_4 _1338_ (.A0(_0266_),
    .A1(_0273_),
    .S(net651),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _1339_ (.A0(\Inst_RegFile_32x4.mem[26][2] ),
    .A1(\Inst_RegFile_32x4.mem[27][2] ),
    .S(net619),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _1340_ (.A0(\Inst_RegFile_32x4.mem[24][2] ),
    .A1(\Inst_RegFile_32x4.mem[25][2] ),
    .S(net619),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _1341_ (.A0(_0275_),
    .A1(_0276_),
    .S(net678),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _1342_ (.A0(\Inst_RegFile_32x4.mem[30][2] ),
    .A1(\Inst_RegFile_32x4.mem[31][2] ),
    .S(net615),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _1343_ (.A0(\Inst_RegFile_32x4.mem[28][2] ),
    .A1(\Inst_RegFile_32x4.mem[29][2] ),
    .S(net615),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _1344_ (.A0(_0278_),
    .A1(_0279_),
    .S(net676),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _1345_ (.A0(_0277_),
    .A1(_0280_),
    .S(net663),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _1346_ (.A0(\Inst_RegFile_32x4.mem[16][2] ),
    .A1(\Inst_RegFile_32x4.mem[17][2] ),
    .S(net618),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _1347_ (.A0(\Inst_RegFile_32x4.mem[18][2] ),
    .A1(\Inst_RegFile_32x4.mem[19][2] ),
    .S(net618),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _1348_ (.A0(_0283_),
    .A1(_0282_),
    .S(net678),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _1349_ (.A0(\Inst_RegFile_32x4.mem[22][2] ),
    .A1(\Inst_RegFile_32x4.mem[23][2] ),
    .S(net617),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _1350_ (.A0(\Inst_RegFile_32x4.mem[20][2] ),
    .A1(\Inst_RegFile_32x4.mem[21][2] ),
    .S(net617),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _1351_ (.A0(_0285_),
    .A1(_0286_),
    .S(net679),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _1352_ (.A0(_0284_),
    .A1(_0287_),
    .S(net664),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_4 _1353_ (.A0(_0281_),
    .A1(_0288_),
    .S(net393),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_4 _1354_ (.A0(_0274_),
    .A1(_0289_),
    .S(_0209_),
    .X(\Inst_RegFile_32x4.AD_comb[2] ));
 sky130_fd_sc_hd__mux2_4 _1355_ (.A0(\Inst_RegFile_32x4.AD_comb[2] ),
    .A1(\Inst_RegFile_32x4.AD_reg[2] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD2));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(\Inst_RegFile_32x4.mem[26][3] ),
    .A1(\Inst_RegFile_32x4.mem[27][3] ),
    .S(net619),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _1357_ (.A0(\Inst_RegFile_32x4.mem[24][3] ),
    .A1(\Inst_RegFile_32x4.mem[25][3] ),
    .S(net619),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _1358_ (.A0(_0290_),
    .A1(_0291_),
    .S(net678),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _1359_ (.A0(\Inst_RegFile_32x4.mem[30][3] ),
    .A1(\Inst_RegFile_32x4.mem[31][3] ),
    .S(net619),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _1360_ (.A0(\Inst_RegFile_32x4.mem[28][3] ),
    .A1(\Inst_RegFile_32x4.mem[29][3] ),
    .S(net615),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _1361_ (.A0(_0293_),
    .A1(_0294_),
    .S(net678),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _1362_ (.A0(_0292_),
    .A1(_0295_),
    .S(net664),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _1363_ (.A0(\Inst_RegFile_32x4.mem[16][3] ),
    .A1(\Inst_RegFile_32x4.mem[17][3] ),
    .S(net617),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _1364_ (.A0(\Inst_RegFile_32x4.mem[18][3] ),
    .A1(\Inst_RegFile_32x4.mem[19][3] ),
    .S(net617),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _1365_ (.A0(_0298_),
    .A1(_0297_),
    .S(net678),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _1366_ (.A0(\Inst_RegFile_32x4.mem[22][3] ),
    .A1(\Inst_RegFile_32x4.mem[23][3] ),
    .S(net617),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _1367_ (.A0(\Inst_RegFile_32x4.mem[20][3] ),
    .A1(\Inst_RegFile_32x4.mem[21][3] ),
    .S(net617),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _1368_ (.A0(_0300_),
    .A1(_0301_),
    .S(net679),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _1369_ (.A0(_0299_),
    .A1(_0302_),
    .S(net664),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _1370_ (.A0(_0296_),
    .A1(_0303_),
    .S(net651),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _1371_ (.A0(\Inst_RegFile_32x4.mem[10][3] ),
    .A1(\Inst_RegFile_32x4.mem[11][3] ),
    .S(net616),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _1372_ (.A0(\Inst_RegFile_32x4.mem[8][3] ),
    .A1(\Inst_RegFile_32x4.mem[9][3] ),
    .S(net614),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _1373_ (.A0(_0305_),
    .A1(_0306_),
    .S(net676),
    .X(_0307_));
 sky130_fd_sc_hd__and2b_1 _1374_ (.A_N(net663),
    .B(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_2 _1375_ (.A0(\Inst_RegFile_32x4.mem[14][3] ),
    .A1(\Inst_RegFile_32x4.mem[15][3] ),
    .S(net395),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_4 _1376_ (.A0(\Inst_RegFile_32x4.mem[12][3] ),
    .A1(\Inst_RegFile_32x4.mem[13][3] ),
    .S(net395),
    .X(_0310_));
 sky130_fd_sc_hd__nand2b_4 _1377_ (.A_N(_0310_),
    .B(net675),
    .Y(_0311_));
 sky130_fd_sc_hd__o211a_1 _1378_ (.A1(net677),
    .A2(_0309_),
    .B1(net663),
    .C1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__or3_4 _1379_ (.A(_0312_),
    .B(_0308_),
    .C(net651),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _1380_ (.A0(\Inst_RegFile_32x4.mem[2][3] ),
    .A1(\Inst_RegFile_32x4.mem[3][3] ),
    .S(net614),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _1381_ (.A0(\Inst_RegFile_32x4.mem[0][3] ),
    .A1(\Inst_RegFile_32x4.mem[1][3] ),
    .S(net615),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _1382_ (.A0(_0314_),
    .A1(_0315_),
    .S(net676),
    .X(_0316_));
 sky130_fd_sc_hd__nand2b_1 _1383_ (.A_N(net663),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__mux2_1 _1384_ (.A0(\Inst_RegFile_32x4.mem[4][3] ),
    .A1(\Inst_RegFile_32x4.mem[5][3] ),
    .S(net612),
    .X(_0318_));
 sky130_fd_sc_hd__nand2b_1 _1385_ (.A_N(_0318_),
    .B(net675),
    .Y(_0319_));
 sky130_fd_sc_hd__mux2_1 _1386_ (.A0(\Inst_RegFile_32x4.mem[6][3] ),
    .A1(\Inst_RegFile_32x4.mem[7][3] ),
    .S(net612),
    .X(_0320_));
 sky130_fd_sc_hd__o211ai_1 _1387_ (.A1(net675),
    .A2(_0320_),
    .B1(_0319_),
    .C1(net662),
    .Y(_0321_));
 sky130_fd_sc_hd__a31oi_1 _1388_ (.A1(_0321_),
    .A2(_0317_),
    .A3(net651),
    .B1(_0209_),
    .Y(_0322_));
 sky130_fd_sc_hd__a22o_1 _1389_ (.A1(_0209_),
    .A2(_0304_),
    .B1(_0322_),
    .B2(_0313_),
    .X(\Inst_RegFile_32x4.AD_comb[3] ));
 sky130_fd_sc_hd__mux2_4 _1390_ (.A0(\Inst_RegFile_32x4.AD_comb[3] ),
    .A1(\Inst_RegFile_32x4.AD_reg[3] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD3));
 sky130_fd_sc_hd__a221o_1 _1391_ (.A1(_0201_),
    .A2(_0202_),
    .B1(_0203_),
    .B2(_0975_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_0323_));
 sky130_fd_sc_hd__mux4_1 _1392_ (.A0(net73),
    .A1(net16),
    .A2(net101),
    .A3(net129),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ),
    .X(_0324_));
 sky130_fd_sc_hd__inv_1 _1393_ (.A(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__a21oi_1 _1394_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(_0325_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ),
    .Y(_0326_));
 sky130_fd_sc_hd__mux4_2 _1395_ (.A0(net648),
    .A1(net636),
    .A2(net668),
    .A3(net447),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0327_));
 sky130_fd_sc_hd__or2_4 _1396_ (.A(_0327_),
    .B(_0977_),
    .X(_0328_));
 sky130_fd_sc_hd__mux4_1 _1397_ (.A0(net115),
    .A1(net672),
    .A2(net658),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0329_));
 sky130_fd_sc_hd__o21a_1 _1398_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0329_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0330_));
 sky130_fd_sc_hd__mux4_2 _1399_ (.A0(net59),
    .A1(net67),
    .A2(net2),
    .A3(net10),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0331_));
 sky130_fd_sc_hd__mux4_2 _1400_ (.A0(net26),
    .A1(net87),
    .A2(net89),
    .A3(net95),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_4 _1401_ (.A0(_0331_),
    .A1(_0332_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0333_));
 sky130_fd_sc_hd__a22oi_4 _1402_ (.A1(_0330_),
    .A2(_0328_),
    .B1(_0333_),
    .B2(_0978_),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_4 _1403_ (.A(_0334_),
    .Y(\Inst_RegFile_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__a221o_1 _1404_ (.A1(_0328_),
    .A2(_0330_),
    .B1(_0978_),
    .B2(_0333_),
    .C1(_0976_),
    .X(_0335_));
 sky130_fd_sc_hd__or2_1 _1405_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .B(net120),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _1406_ (.A0(net80),
    .A1(net112),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0337_));
 sky130_fd_sc_hd__inv_2 _1407_ (.A(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__o21ai_1 _1408_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_0338_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .Y(_0339_));
 sky130_fd_sc_hd__a31o_1 _1409_ (.A1(_0335_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ),
    .A3(_0336_),
    .B1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__mux4_2 _1410_ (.A0(net65),
    .A1(net8),
    .A2(net110),
    .A3(net121),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_0341_));
 sky130_fd_sc_hd__o21a_1 _1411_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(_0341_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_4 _1412_ (.A1(_0323_),
    .A2(_0326_),
    .B1(_0340_),
    .B2(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _1413_ (.A0(\Inst_RegFile_32x4.mem[26][0] ),
    .A1(\Inst_RegFile_32x4.mem[27][0] ),
    .S(net628),
    .X(_0344_));
 sky130_fd_sc_hd__mux4_1 _1414_ (.A0(net692),
    .A1(net674),
    .A2(net660),
    .A3(net656),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0345_));
 sky130_fd_sc_hd__or2_1 _1415_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .B(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__mux4_2 _1416_ (.A0(net650),
    .A1(net684),
    .A2(net431),
    .A3(net642),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0347_));
 sky130_fd_sc_hd__o21a_1 _1417_ (.A1(_0347_),
    .A2(_0981_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ),
    .X(_0348_));
 sky130_fd_sc_hd__mux4_1 _1418_ (.A0(net61),
    .A1(net69),
    .A2(net783),
    .A3(net12),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0349_));
 sky130_fd_sc_hd__mux4_1 _1419_ (.A0(net89),
    .A1(net97),
    .A2(net111),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _1420_ (.A0(_0349_),
    .A1(_0350_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0351_));
 sky130_fd_sc_hd__a22o_4 _1421_ (.A1(_0346_),
    .A2(_0348_),
    .B1(_0351_),
    .B2(_0982_),
    .X(\Inst_RegFile_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1422_ (.A0(net17),
    .A1(net102),
    .A2(net130),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ),
    .X(_0352_));
 sky130_fd_sc_hd__and2b_1 _1423_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .B(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__a21o_1 _1424_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(_0205_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_0354_));
 sky130_fd_sc_hd__mux4_1 _1425_ (.A0(net692),
    .A1(net672),
    .A2(net658),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0355_));
 sky130_fd_sc_hd__mux4_2 _1426_ (.A0(net648),
    .A1(net428),
    .A2(net431),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_4 _1427_ (.A0(_0355_),
    .A1(_0356_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0357_));
 sky130_fd_sc_hd__mux4_1 _1428_ (.A0(net59),
    .A1(net67),
    .A2(net2),
    .A3(net10),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0358_));
 sky130_fd_sc_hd__mux4_1 _1429_ (.A0(net87),
    .A1(net95),
    .A2(net113),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _1430_ (.A0(_0358_),
    .A1(_0359_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_4 _1431_ (.A0(_0360_),
    .A1(_0357_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ),
    .X(\Inst_RegFile_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__o21ai_1 _1432_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_0984_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_0361_));
 sky130_fd_sc_hd__a21o_1 _1433_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .B1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _1434_ (.A0(net22),
    .A1(net107),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_0363_));
 sky130_fd_sc_hd__o211a_1 _1435_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0363_),
    .B1(_0362_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .X(_0364_));
 sky130_fd_sc_hd__mux4_1 _1436_ (.A0(net83),
    .A1(net10),
    .A2(net95),
    .A3(net123),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ),
    .X(_0365_));
 sky130_fd_sc_hd__inv_2 _1437_ (.A(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__o21ai_1 _1438_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(_0366_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ),
    .Y(_0367_));
 sky130_fd_sc_hd__o22a_1 _1439_ (.A1(_0354_),
    .A2(_0353_),
    .B1(_0364_),
    .B2(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(\Inst_RegFile_32x4.mem[24][0] ),
    .A1(\Inst_RegFile_32x4.mem[25][0] ),
    .S(net628),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _1441_ (.A0(_0369_),
    .A1(_0344_),
    .S(net688),
    .X(_0370_));
 sky130_fd_sc_hd__mux4_1 _1442_ (.A0(net139),
    .A1(net672),
    .A2(net658),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0371_));
 sky130_fd_sc_hd__mux4_2 _1443_ (.A0(net648),
    .A1(net636),
    .A2(net667),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_4 _1444_ (.A0(_0371_),
    .A1(_0372_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0373_));
 sky130_fd_sc_hd__mux4_1 _1445_ (.A0(net59),
    .A1(net67),
    .A2(net2),
    .A3(net10),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0374_));
 sky130_fd_sc_hd__mux4_1 _1446_ (.A0(net87),
    .A1(net95),
    .A2(net89),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _1447_ (.A0(_0374_),
    .A1(_0375_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_4 _1448_ (.A0(_0376_),
    .A1(_0373_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Inst_RegFile_switch_matrix.JW2BEG4 ));
 sky130_fd_sc_hd__mux4_2 _1449_ (.A0(net82),
    .A1(net782),
    .A2(net118),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ),
    .X(_0377_));
 sky130_fd_sc_hd__mux4_2 _1450_ (.A0(net63),
    .A1(net91),
    .A2(net26),
    .A3(net119),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_2 _1451_ (.A0(_0377_),
    .A1(_0378_),
    .S(_0985_),
    .X(_0379_));
 sky130_fd_sc_hd__mux4_2 _1452_ (.A0(net137),
    .A1(net672),
    .A2(net658),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0380_));
 sky130_fd_sc_hd__and2b_1 _1453_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .B(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__mux4_2 _1454_ (.A0(net648),
    .A1(net683),
    .A2(net667),
    .A3(net447),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0382_));
 sky130_fd_sc_hd__a21bo_1 _1455_ (.A1(_0382_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ),
    .X(_0383_));
 sky130_fd_sc_hd__mux4_1 _1456_ (.A0(net61),
    .A1(net69),
    .A2(net783),
    .A3(net12),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0384_));
 sky130_fd_sc_hd__mux4_1 _1457_ (.A0(net87),
    .A1(net97),
    .A2(net89),
    .A3(net692),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _1458_ (.A0(_0384_),
    .A1(_0385_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .X(_0386_));
 sky130_fd_sc_hd__o22a_4 _1459_ (.A1(_0383_),
    .A2(_0381_),
    .B1(_0386_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_RegFile_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1460_ (.A0(net70),
    .A1(net13),
    .A2(net126),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(net71),
    .A1(net14),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _1462_ (.A(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ),
    .B(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _1463_ (.A0(net99),
    .A1(net127),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_0390_));
 sky130_fd_sc_hd__o211a_1 _1464_ (.A1(_0988_),
    .A2(_0390_),
    .B1(_0389_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_0391_));
 sky130_fd_sc_hd__a21o_1 _1465_ (.A1(_0985_),
    .A2(_0387_),
    .B1(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_4 _1466_ (.A0(_0392_),
    .A1(_0379_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ),
    .X(_0393_));
 sky130_fd_sc_hd__inv_8 _1467_ (.A(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__mux2_1 _1468_ (.A0(\Inst_RegFile_32x4.mem[28][0] ),
    .A1(\Inst_RegFile_32x4.mem[29][0] ),
    .S(net624),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _1469_ (.A0(\Inst_RegFile_32x4.mem[30][0] ),
    .A1(\Inst_RegFile_32x4.mem[31][0] ),
    .S(net624),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _1470_ (.A0(_0395_),
    .A1(_0396_),
    .S(net687),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _1471_ (.A0(_0370_),
    .A1(_0397_),
    .S(net644),
    .X(_0398_));
 sky130_fd_sc_hd__mux4_1 _1472_ (.A0(net692),
    .A1(net673),
    .A2(net659),
    .A3(net655),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0399_));
 sky130_fd_sc_hd__mux4_1 _1473_ (.A0(net648),
    .A1(net683),
    .A2(net667),
    .A3(net642),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_2 _1474_ (.A0(_0399_),
    .A1(_0400_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0401_));
 sky130_fd_sc_hd__mux4_1 _1475_ (.A0(net61),
    .A1(net69),
    .A2(net83),
    .A3(net783),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0402_));
 sky130_fd_sc_hd__mux4_1 _1476_ (.A0(net12),
    .A1(net89),
    .A2(net97),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(_0402_),
    .A1(_0403_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_4 _1478_ (.A0(_0404_),
    .A1(_0401_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ),
    .X(\Inst_RegFile_switch_matrix.JN2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _1479_ (.A0(_0153_),
    .A1(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_0405_));
 sky130_fd_sc_hd__mux4_2 _1480_ (.A0(net15),
    .A1(net128),
    .A2(net100),
    .A3(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0406_));
 sky130_fd_sc_hd__mux4_2 _1481_ (.A0(net75),
    .A1(net18),
    .A2(net103),
    .A3(net131),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0407_));
 sky130_fd_sc_hd__mux4_2 _1482_ (.A0(net64),
    .A1(net92),
    .A2(_0406_),
    .A3(_0407_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_4 _1483_ (.A0(_0408_),
    .A1(_0405_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(\Inst_RegFile_32x4.mem[16][0] ),
    .A1(\Inst_RegFile_32x4.mem[17][0] ),
    .S(net627),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _1485_ (.A0(\Inst_RegFile_32x4.mem[18][0] ),
    .A1(\Inst_RegFile_32x4.mem[19][0] ),
    .S(net627),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(_0410_),
    .A1(_0411_),
    .S(net688),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _1487_ (.A0(\Inst_RegFile_32x4.mem[20][0] ),
    .A1(\Inst_RegFile_32x4.mem[21][0] ),
    .S(net626),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _1488_ (.A0(\Inst_RegFile_32x4.mem[22][0] ),
    .A1(\Inst_RegFile_32x4.mem[23][0] ),
    .S(net626),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(_0413_),
    .A1(_0414_),
    .S(_0343_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _1490_ (.A0(_0412_),
    .A1(_0415_),
    .S(net645),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _1491_ (.A0(_0398_),
    .A1(_0416_),
    .S(_0394_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _1492_ (.A0(\Inst_RegFile_32x4.mem[8][0] ),
    .A1(\Inst_RegFile_32x4.mem[9][0] ),
    .S(net623),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _1493_ (.A0(\Inst_RegFile_32x4.mem[10][0] ),
    .A1(\Inst_RegFile_32x4.mem[11][0] ),
    .S(net623),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _1494_ (.A0(_0418_),
    .A1(_0419_),
    .S(net685),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(\Inst_RegFile_32x4.mem[12][0] ),
    .A1(\Inst_RegFile_32x4.mem[13][0] ),
    .S(net432),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _1496_ (.A0(\Inst_RegFile_32x4.mem[14][0] ),
    .A1(\Inst_RegFile_32x4.mem[15][0] ),
    .S(net432),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _1497_ (.A0(_0421_),
    .A1(_0422_),
    .S(net685),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _1498_ (.A0(_0420_),
    .A1(_0423_),
    .S(net417),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _1499_ (.A0(\Inst_RegFile_32x4.mem[2][0] ),
    .A1(\Inst_RegFile_32x4.mem[3][0] ),
    .S(net625),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _1500_ (.A0(\Inst_RegFile_32x4.mem[0][0] ),
    .A1(\Inst_RegFile_32x4.mem[1][0] ),
    .S(net624),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _1501_ (.A0(_0426_),
    .A1(_0425_),
    .S(net687),
    .X(_0427_));
 sky130_fd_sc_hd__and2b_1 _1502_ (.A_N(net417),
    .B(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _1503_ (.A0(\Inst_RegFile_32x4.mem[6][0] ),
    .A1(\Inst_RegFile_32x4.mem[7][0] ),
    .S(net432),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _1504_ (.A0(\Inst_RegFile_32x4.mem[4][0] ),
    .A1(\Inst_RegFile_32x4.mem[5][0] ),
    .S(net432),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _1505_ (.A0(_0430_),
    .A1(_0429_),
    .S(net686),
    .X(_0431_));
 sky130_fd_sc_hd__a21o_1 _1506_ (.A1(net417),
    .A2(_0431_),
    .B1(_0393_),
    .X(_0432_));
 sky130_fd_sc_hd__o22a_1 _1507_ (.A1(net397),
    .A2(_0424_),
    .B1(_0432_),
    .B2(_0428_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_4 _1508_ (.A0(_0433_),
    .A1(_0417_),
    .S(_0409_),
    .X(\Inst_RegFile_32x4.BD_comb[0] ));
 sky130_fd_sc_hd__mux2_4 _1509_ (.A0(\Inst_RegFile_32x4.BD_comb[0] ),
    .A1(\Inst_RegFile_32x4.BD_reg[0] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD0));
 sky130_fd_sc_hd__mux2_1 _1510_ (.A0(\Inst_RegFile_32x4.mem[26][1] ),
    .A1(\Inst_RegFile_32x4.mem[27][1] ),
    .S(net628),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _1511_ (.A0(\Inst_RegFile_32x4.mem[24][1] ),
    .A1(\Inst_RegFile_32x4.mem[25][1] ),
    .S(net628),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(_0435_),
    .A1(_0434_),
    .S(net688),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _1513_ (.A0(\Inst_RegFile_32x4.mem[28][1] ),
    .A1(\Inst_RegFile_32x4.mem[29][1] ),
    .S(net624),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _1514_ (.A0(\Inst_RegFile_32x4.mem[30][1] ),
    .A1(\Inst_RegFile_32x4.mem[31][1] ),
    .S(net624),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _1515_ (.A0(_0437_),
    .A1(_0438_),
    .S(net687),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _1516_ (.A0(_0436_),
    .A1(_0439_),
    .S(net645),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _1517_ (.A0(\Inst_RegFile_32x4.mem[16][1] ),
    .A1(\Inst_RegFile_32x4.mem[17][1] ),
    .S(net627),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _1518_ (.A0(\Inst_RegFile_32x4.mem[18][1] ),
    .A1(\Inst_RegFile_32x4.mem[19][1] ),
    .S(net627),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _1519_ (.A0(_0441_),
    .A1(_0442_),
    .S(net688),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _1520_ (.A0(\Inst_RegFile_32x4.mem[20][1] ),
    .A1(\Inst_RegFile_32x4.mem[21][1] ),
    .S(net627),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _1521_ (.A0(\Inst_RegFile_32x4.mem[22][1] ),
    .A1(\Inst_RegFile_32x4.mem[23][1] ),
    .S(net626),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_4 _1522_ (.A0(_0444_),
    .A1(_0445_),
    .S(_0343_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_4 _1523_ (.A0(_0443_),
    .A1(_0446_),
    .S(net645),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_4 _1524_ (.A0(_0440_),
    .A1(_0447_),
    .S(_0394_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(\Inst_RegFile_32x4.mem[8][1] ),
    .A1(\Inst_RegFile_32x4.mem[9][1] ),
    .S(net622),
    .X(_0449_));
 sky130_fd_sc_hd__nor2_1 _1526_ (.A(net685),
    .B(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__nand2_1 _1527_ (.A(\Inst_RegFile_32x4.mem[11][1] ),
    .B(net622),
    .Y(_0451_));
 sky130_fd_sc_hd__o211a_1 _1528_ (.A1(_0993_),
    .A2(net622),
    .B1(net685),
    .C1(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _1529_ (.A0(\Inst_RegFile_32x4.mem[14][1] ),
    .A1(\Inst_RegFile_32x4.mem[15][1] ),
    .S(net621),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _1530_ (.A0(\Inst_RegFile_32x4.mem[12][1] ),
    .A1(\Inst_RegFile_32x4.mem[13][1] ),
    .S(net621),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _1531_ (.A0(_0454_),
    .A1(_0453_),
    .S(net686),
    .X(_0455_));
 sky130_fd_sc_hd__nand2_1 _1532_ (.A(net417),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__o31a_1 _1533_ (.A1(net417),
    .A2(_0450_),
    .A3(_0452_),
    .B1(_0393_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _1534_ (.A0(\Inst_RegFile_32x4.mem[2][1] ),
    .A1(\Inst_RegFile_32x4.mem[3][1] ),
    .S(net622),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _1535_ (.A0(\Inst_RegFile_32x4.mem[0][1] ),
    .A1(\Inst_RegFile_32x4.mem[1][1] ),
    .S(net622),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _1536_ (.A0(_0459_),
    .A1(_0458_),
    .S(net685),
    .X(_0460_));
 sky130_fd_sc_hd__and2b_1 _1537_ (.A_N(net644),
    .B(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _1538_ (.A0(\Inst_RegFile_32x4.mem[4][1] ),
    .A1(\Inst_RegFile_32x4.mem[5][1] ),
    .S(net432),
    .X(_0462_));
 sky130_fd_sc_hd__or2_1 _1539_ (.A(net686),
    .B(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _1540_ (.A0(\Inst_RegFile_32x4.mem[6][1] ),
    .A1(\Inst_RegFile_32x4.mem[7][1] ),
    .S(net620),
    .X(_0464_));
 sky130_fd_sc_hd__inv_1 _1541_ (.A(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2_1 _1542_ (.A(net686),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__a31o_1 _1543_ (.A1(net643),
    .A2(_0463_),
    .A3(_0466_),
    .B1(_0393_),
    .X(_0467_));
 sky130_fd_sc_hd__o2bb2a_1 _1544_ (.A1_N(_0456_),
    .A2_N(_0457_),
    .B1(_0461_),
    .B2(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_4 _1545_ (.A0(_0468_),
    .A1(_0448_),
    .S(_0409_),
    .X(\Inst_RegFile_32x4.BD_comb[1] ));
 sky130_fd_sc_hd__mux2_4 _1546_ (.A0(\Inst_RegFile_32x4.BD_comb[1] ),
    .A1(\Inst_RegFile_32x4.BD_reg[1] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD1));
 sky130_fd_sc_hd__mux2_1 _1547_ (.A0(\Inst_RegFile_32x4.mem[26][3] ),
    .A1(\Inst_RegFile_32x4.mem[27][3] ),
    .S(net628),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _1548_ (.A0(\Inst_RegFile_32x4.mem[24][3] ),
    .A1(\Inst_RegFile_32x4.mem[25][3] ),
    .S(net628),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _1549_ (.A0(_0470_),
    .A1(_0469_),
    .S(net688),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _1550_ (.A0(\Inst_RegFile_32x4.mem[28][3] ),
    .A1(\Inst_RegFile_32x4.mem[29][3] ),
    .S(net624),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _1551_ (.A0(\Inst_RegFile_32x4.mem[30][3] ),
    .A1(\Inst_RegFile_32x4.mem[31][3] ),
    .S(net628),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(_0472_),
    .A1(_0473_),
    .S(net687),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _1553_ (.A0(_0471_),
    .A1(_0474_),
    .S(net645),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(\Inst_RegFile_32x4.mem[16][3] ),
    .A1(\Inst_RegFile_32x4.mem[17][3] ),
    .S(net626),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _1555_ (.A0(\Inst_RegFile_32x4.mem[18][3] ),
    .A1(\Inst_RegFile_32x4.mem[19][3] ),
    .S(net626),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _1556_ (.A0(_0476_),
    .A1(_0477_),
    .S(net688),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _1557_ (.A0(\Inst_RegFile_32x4.mem[20][3] ),
    .A1(\Inst_RegFile_32x4.mem[21][3] ),
    .S(net626),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(\Inst_RegFile_32x4.mem[22][3] ),
    .A1(\Inst_RegFile_32x4.mem[23][3] ),
    .S(net626),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _1559_ (.A0(_0479_),
    .A1(_0480_),
    .S(net688),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _1560_ (.A0(_0478_),
    .A1(_0481_),
    .S(net645),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _1561_ (.A0(_0475_),
    .A1(_0482_),
    .S(_0394_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _1562_ (.A0(\Inst_RegFile_32x4.mem[10][3] ),
    .A1(\Inst_RegFile_32x4.mem[11][3] ),
    .S(net623),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _1563_ (.A0(\Inst_RegFile_32x4.mem[8][3] ),
    .A1(\Inst_RegFile_32x4.mem[9][3] ),
    .S(net623),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _1564_ (.A0(_0485_),
    .A1(_0484_),
    .S(net685),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _1565_ (.A0(\Inst_RegFile_32x4.mem[12][3] ),
    .A1(\Inst_RegFile_32x4.mem[13][3] ),
    .S(net621),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _1566_ (.A0(\Inst_RegFile_32x4.mem[14][3] ),
    .A1(\Inst_RegFile_32x4.mem[15][3] ),
    .S(net621),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(_0487_),
    .A1(_0488_),
    .S(net686),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_2 _1568_ (.A0(_0486_),
    .A1(_0489_),
    .S(net643),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _1569_ (.A0(\Inst_RegFile_32x4.mem[0][3] ),
    .A1(\Inst_RegFile_32x4.mem[1][3] ),
    .S(net625),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _1570_ (.A0(\Inst_RegFile_32x4.mem[2][3] ),
    .A1(\Inst_RegFile_32x4.mem[3][3] ),
    .S(net622),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _1571_ (.A0(_0491_),
    .A1(_0492_),
    .S(net686),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _1572_ (.A0(\Inst_RegFile_32x4.mem[4][3] ),
    .A1(\Inst_RegFile_32x4.mem[5][3] ),
    .S(net620),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _1573_ (.A0(\Inst_RegFile_32x4.mem[6][3] ),
    .A1(\Inst_RegFile_32x4.mem[7][3] ),
    .S(net620),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _1574_ (.A0(_0494_),
    .A1(_0495_),
    .S(net686),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _1575_ (.A0(_0493_),
    .A1(_0496_),
    .S(net644),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_4 _1576_ (.A0(_0490_),
    .A1(_0497_),
    .S(_0394_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_4 _1577_ (.A0(_0498_),
    .A1(_0483_),
    .S(_0409_),
    .X(\Inst_RegFile_32x4.BD_comb[3] ));
 sky130_fd_sc_hd__mux2_4 _1578_ (.A0(\Inst_RegFile_32x4.BD_comb[3] ),
    .A1(\Inst_RegFile_32x4.BD_reg[3] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD3));
 sky130_fd_sc_hd__mux2_1 _1579_ (.A0(\Inst_RegFile_32x4.mem[26][2] ),
    .A1(\Inst_RegFile_32x4.mem[27][2] ),
    .S(net628),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _1580_ (.A0(\Inst_RegFile_32x4.mem[24][2] ),
    .A1(\Inst_RegFile_32x4.mem[25][2] ),
    .S(net628),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _1581_ (.A0(_0500_),
    .A1(_0499_),
    .S(net688),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _1582_ (.A0(\Inst_RegFile_32x4.mem[28][2] ),
    .A1(\Inst_RegFile_32x4.mem[29][2] ),
    .S(net624),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _1583_ (.A0(\Inst_RegFile_32x4.mem[30][2] ),
    .A1(\Inst_RegFile_32x4.mem[31][2] ),
    .S(net624),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _1584_ (.A0(_0502_),
    .A1(_0503_),
    .S(net687),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _1585_ (.A0(_0501_),
    .A1(_0504_),
    .S(net644),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _1586_ (.A0(\Inst_RegFile_32x4.mem[16][2] ),
    .A1(\Inst_RegFile_32x4.mem[17][2] ),
    .S(net626),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _1587_ (.A0(\Inst_RegFile_32x4.mem[18][2] ),
    .A1(\Inst_RegFile_32x4.mem[19][2] ),
    .S(net627),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _1588_ (.A0(_0506_),
    .A1(_0507_),
    .S(net688),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _1589_ (.A0(\Inst_RegFile_32x4.mem[20][2] ),
    .A1(\Inst_RegFile_32x4.mem[21][2] ),
    .S(net626),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _1590_ (.A0(\Inst_RegFile_32x4.mem[22][2] ),
    .A1(\Inst_RegFile_32x4.mem[23][2] ),
    .S(net626),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _1591_ (.A0(_0509_),
    .A1(_0510_),
    .S(net688),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _1592_ (.A0(_0508_),
    .A1(_0511_),
    .S(net645),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_4 _1593_ (.A0(_0505_),
    .A1(_0512_),
    .S(_0394_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _1594_ (.A0(\Inst_RegFile_32x4.mem[8][2] ),
    .A1(\Inst_RegFile_32x4.mem[9][2] ),
    .S(net623),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _1595_ (.A0(\Inst_RegFile_32x4.mem[10][2] ),
    .A1(\Inst_RegFile_32x4.mem[11][2] ),
    .S(net623),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _1596_ (.A0(_0514_),
    .A1(_0515_),
    .S(net685),
    .X(_0516_));
 sky130_fd_sc_hd__and2b_1 _1597_ (.A_N(net643),
    .B(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__and2b_1 _1598_ (.A_N(net622),
    .B(\Inst_RegFile_32x4.mem[14][2] ),
    .X(_0518_));
 sky130_fd_sc_hd__a21bo_1 _1599_ (.A1(\Inst_RegFile_32x4.mem[15][2] ),
    .A2(net622),
    .B1_N(net685),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _1600_ (.A0(\Inst_RegFile_32x4.mem[12][2] ),
    .A1(\Inst_RegFile_32x4.mem[13][2] ),
    .S(net621),
    .X(_0520_));
 sky130_fd_sc_hd__o221a_1 _1601_ (.A1(_0518_),
    .A2(_0519_),
    .B1(_0520_),
    .B2(net685),
    .C1(net644),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _1602_ (.A0(\Inst_RegFile_32x4.mem[2][2] ),
    .A1(\Inst_RegFile_32x4.mem[3][2] ),
    .S(net622),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _1603_ (.A0(\Inst_RegFile_32x4.mem[0][2] ),
    .A1(\Inst_RegFile_32x4.mem[1][2] ),
    .S(net622),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _1604_ (.A0(_0523_),
    .A1(_0522_),
    .S(net685),
    .X(_0524_));
 sky130_fd_sc_hd__and2b_1 _1605_ (.A_N(net643),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _1606_ (.A0(\Inst_RegFile_32x4.mem[4][2] ),
    .A1(\Inst_RegFile_32x4.mem[5][2] ),
    .S(net620),
    .X(_0526_));
 sky130_fd_sc_hd__or2_1 _1607_ (.A(net686),
    .B(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _1608_ (.A0(\Inst_RegFile_32x4.mem[6][2] ),
    .A1(\Inst_RegFile_32x4.mem[7][2] ),
    .S(net620),
    .X(_0528_));
 sky130_fd_sc_hd__inv_1 _1609_ (.A(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2_1 _1610_ (.A(net686),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__a31o_1 _1611_ (.A1(_0527_),
    .A2(net643),
    .A3(_0530_),
    .B1(_0393_),
    .X(_0531_));
 sky130_fd_sc_hd__o32a_4 _1612_ (.A1(net397),
    .A2(_0517_),
    .A3(_0521_),
    .B1(_0531_),
    .B2(_0525_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_4 _1613_ (.A0(_0532_),
    .A1(_0513_),
    .S(_0409_),
    .X(\Inst_RegFile_32x4.BD_comb[2] ));
 sky130_fd_sc_hd__mux2_4 _1614_ (.A0(\Inst_RegFile_32x4.BD_comb[2] ),
    .A1(\Inst_RegFile_32x4.BD_reg[2] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD2));
 sky130_fd_sc_hd__mux4_1 _1615_ (.A0(net692),
    .A1(net673),
    .A2(net659),
    .A3(net655),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0533_));
 sky130_fd_sc_hd__or2_1 _1616_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .B(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__mux4_2 _1617_ (.A0(net648),
    .A1(net428),
    .A2(net667),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0535_));
 sky130_fd_sc_hd__o21a_1 _1618_ (.A1(_0968_),
    .A2(_0535_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0536_));
 sky130_fd_sc_hd__mux4_1 _1619_ (.A0(net418),
    .A1(net67),
    .A2(net85),
    .A3(net2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0537_));
 sky130_fd_sc_hd__mux4_1 _1620_ (.A0(net10),
    .A1(net87),
    .A2(net95),
    .A3(net115),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _1621_ (.A0(_0537_),
    .A1(_0538_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0539_));
 sky130_fd_sc_hd__a22o_4 _1622_ (.A1(_0534_),
    .A2(_0536_),
    .B1(_0539_),
    .B2(_0969_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG4 ));
 sky130_fd_sc_hd__mux4_2 _1623_ (.A0(net81),
    .A1(net23),
    .A2(net109),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_0540_));
 sky130_fd_sc_hd__mux4_2 _1624_ (.A0(net69),
    .A1(net12),
    .A2(net97),
    .A3(net136),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_4 _1625_ (.A0(_0541_),
    .A1(_0540_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _1626_ (.A0(net104),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _1627_ (.A0(net76),
    .A1(net19),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0544_));
 sky130_fd_sc_hd__and2b_1 _1628_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__a211o_1 _1629_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ),
    .A2(_0543_),
    .B1(_0545_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _1630_ (.A0(net77),
    .A1(net20),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_0547_));
 sky130_fd_sc_hd__inv_1 _1631_ (.A(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__mux2_1 _1632_ (.A0(net105),
    .A1(net133),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_0549_));
 sky130_fd_sc_hd__nand2_1 _1633_ (.A(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__o211a_1 _1634_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ),
    .A2(_0548_),
    .B1(_0550_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .X(_0551_));
 sky130_fd_sc_hd__nor2_1 _1635_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__a22o_4 _1636_ (.A1(_0542_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ),
    .B1(_0546_),
    .B2(_0552_),
    .X(B_ADR0));
 sky130_fd_sc_hd__mux4_2 _1637_ (.A0(net691),
    .A1(net670),
    .A2(net657),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0553_));
 sky130_fd_sc_hd__mux4_2 _1638_ (.A0(net681),
    .A1(net634),
    .A2(net665),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_4 _1639_ (.A0(_0553_),
    .A1(_0554_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0555_));
 sky130_fd_sc_hd__mux4_1 _1640_ (.A0(net66),
    .A1(net78),
    .A2(net784),
    .A3(net9),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0556_));
 sky130_fd_sc_hd__mux4_1 _1641_ (.A0(net782),
    .A1(net94),
    .A2(net122),
    .A3(net139),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _1642_ (.A0(_0556_),
    .A1(_0557_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_4 _1643_ (.A0(_0558_),
    .A1(_0555_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ),
    .X(\Inst_RegFile_switch_matrix.JN2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1644_ (.A0(net69),
    .A1(net97),
    .A2(net25),
    .A3(net125),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ),
    .X(_0559_));
 sky130_fd_sc_hd__mux4_2 _1645_ (.A0(net81),
    .A1(net8),
    .A2(net121),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_4 _1646_ (.A0(_0559_),
    .A1(_0560_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_0561_));
 sky130_fd_sc_hd__mux4_1 _1647_ (.A0(net76),
    .A1(net19),
    .A2(net132),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ),
    .X(_0562_));
 sky130_fd_sc_hd__mux4_2 _1648_ (.A0(net77),
    .A1(net20),
    .A2(net105),
    .A3(net133),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _1649_ (.A0(_0562_),
    .A1(_0563_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_4 _1650_ (.A0(_0564_),
    .A1(_0561_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ),
    .X(A_ADR0));
 sky130_fd_sc_hd__mux4_1 _1651_ (.A0(net135),
    .A1(net672),
    .A2(net658),
    .A3(net648),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0565_));
 sky130_fd_sc_hd__mux4_2 _1652_ (.A0(net683),
    .A1(net636),
    .A2(net667),
    .A3(net641),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_4 _1653_ (.A0(_0565_),
    .A1(_0566_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0567_));
 sky130_fd_sc_hd__mux4_1 _1654_ (.A0(net59),
    .A1(net65),
    .A2(net84),
    .A3(net8),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0568_));
 sky130_fd_sc_hd__mux4_1 _1655_ (.A0(net22),
    .A1(net93),
    .A2(net109),
    .A3(net121),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _1656_ (.A0(_0568_),
    .A1(_0569_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_4 _1657_ (.A0(_0570_),
    .A1(_0567_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ),
    .X(\Inst_RegFile_switch_matrix.JW2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1658_ (.A0(net690),
    .A1(net670),
    .A2(net661),
    .A3(net647),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0571_));
 sky130_fd_sc_hd__mux4_2 _1659_ (.A0(net681),
    .A1(net634),
    .A2(net665),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_4 _1660_ (.A0(_0571_),
    .A1(_0572_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .X(_0573_));
 sky130_fd_sc_hd__mux4_1 _1661_ (.A0(net65),
    .A1(net8),
    .A2(net2),
    .A3(net25),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0574_));
 sky130_fd_sc_hd__mux4_1 _1662_ (.A0(net781),
    .A1(net93),
    .A2(net109),
    .A3(net121),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _1663_ (.A0(_0574_),
    .A1(_0575_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_4 _1664_ (.A0(_0576_),
    .A1(_0573_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ),
    .X(\Inst_RegFile_switch_matrix.JS2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1665_ (.A0(net690),
    .A1(net670),
    .A2(net657),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0577_));
 sky130_fd_sc_hd__mux4_2 _1666_ (.A0(net680),
    .A1(net633),
    .A2(net666),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_4 _1667_ (.A0(_0577_),
    .A1(_0578_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0579_));
 sky130_fd_sc_hd__mux4_1 _1668_ (.A0(net59),
    .A1(net65),
    .A2(net81),
    .A3(net8),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0580_));
 sky130_fd_sc_hd__mux4_1 _1669_ (.A0(net781),
    .A1(net93),
    .A2(net112),
    .A3(net121),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _1670_ (.A0(_0580_),
    .A1(_0581_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_4 _1671_ (.A0(_0582_),
    .A1(_0579_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ),
    .X(\Inst_RegFile_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1672_ (.A0(net690),
    .A1(net673),
    .A2(net658),
    .A3(net649),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0583_));
 sky130_fd_sc_hd__or2_1 _1673_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .B(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__mux4_2 _1674_ (.A0(net684),
    .A1(net636),
    .A2(net668),
    .A3(net642),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .X(_0585_));
 sky130_fd_sc_hd__o21a_1 _1675_ (.A1(_0585_),
    .A2(_1007_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0586_));
 sky130_fd_sc_hd__mux4_1 _1676_ (.A0(net65),
    .A1(net2),
    .A2(net81),
    .A3(net8),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .X(_0587_));
 sky130_fd_sc_hd__mux4_1 _1677_ (.A0(net781),
    .A1(net93),
    .A2(net121),
    .A3(net138),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _1678_ (.A0(_0587_),
    .A1(_0588_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .X(_0589_));
 sky130_fd_sc_hd__a22o_4 _1679_ (.A1(_0586_),
    .A2(_0584_),
    .B1(_0589_),
    .B2(_1008_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1680_ (.A0(net691),
    .A1(net414),
    .A2(net407),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0590_));
 sky130_fd_sc_hd__nor2_1 _1681_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__mux4_2 _1682_ (.A0(net680),
    .A1(net427),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0592_));
 sky130_fd_sc_hd__o21ai_2 _1683_ (.A1(_0592_),
    .A2(_1009_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0593_));
 sky130_fd_sc_hd__mux4_1 _1684_ (.A0(net58),
    .A1(net7),
    .A2(net64),
    .A3(net782),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0594_));
 sky130_fd_sc_hd__nor2_1 _1685_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .B(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__mux4_1 _1686_ (.A0(net92),
    .A1(net108),
    .A2(net111),
    .A3(net120),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0596_));
 sky130_fd_sc_hd__nor2_1 _1687_ (.A(_1009_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__o32a_4 _1688_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0595_),
    .A3(_0597_),
    .B1(_0593_),
    .B2(_0591_),
    .X(_0598_));
 sky130_fd_sc_hd__inv_2 _1689_ (.A(_0598_),
    .Y(\Inst_RegFile_switch_matrix.JW2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1690_ (.A0(net691),
    .A1(net670),
    .A2(net407),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0599_));
 sky130_fd_sc_hd__or2_1 _1691_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .B(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__mux4_2 _1692_ (.A0(net680),
    .A1(net427),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0601_));
 sky130_fd_sc_hd__o21a_1 _1693_ (.A1(_1011_),
    .A2(_0601_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0602_));
 sky130_fd_sc_hd__mux4_1 _1694_ (.A0(net64),
    .A1(net7),
    .A2(net1),
    .A3(net782),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0603_));
 sky130_fd_sc_hd__mux4_1 _1695_ (.A0(net92),
    .A1(net108),
    .A2(net120),
    .A3(net137),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _1696_ (.A0(_0603_),
    .A1(_0604_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0605_));
 sky130_fd_sc_hd__a22o_1 _1697_ (.A1(_0602_),
    .A2(_0600_),
    .B1(_0605_),
    .B2(_1012_),
    .X(\Inst_RegFile_switch_matrix.JS2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1698_ (.A0(net134),
    .A1(net671),
    .A2(net653),
    .A3(net647),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0606_));
 sky130_fd_sc_hd__or2_1 _1699_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ),
    .B(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__mux4_2 _1700_ (.A0(net682),
    .A1(net635),
    .A2(net666),
    .A3(net640),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0608_));
 sky130_fd_sc_hd__o21a_1 _1701_ (.A1(_0608_),
    .A2(_1013_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0609_));
 sky130_fd_sc_hd__mux4_1 _1702_ (.A0(net7),
    .A1(net92),
    .A2(net782),
    .A3(net120),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0610_));
 sky130_fd_sc_hd__mux4_1 _1703_ (.A0(net58),
    .A1(net64),
    .A2(net80),
    .A3(net83),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(_0610_),
    .A1(_0611_),
    .S(_1013_),
    .X(_0612_));
 sky130_fd_sc_hd__a22o_4 _1705_ (.A1(_0609_),
    .A2(_0607_),
    .B1(_0612_),
    .B2(_1014_),
    .X(\Inst_RegFile_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1706_ (.A0(net680),
    .A1(net633),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0613_));
 sky130_fd_sc_hd__or2_4 _1707_ (.A(_1015_),
    .B(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__mux4_1 _1708_ (.A0(net691),
    .A1(net670),
    .A2(net652),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0615_));
 sky130_fd_sc_hd__o21a_1 _1709_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .A2(_0615_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0616_));
 sky130_fd_sc_hd__mux4_1 _1710_ (.A0(net64),
    .A1(net1),
    .A2(net80),
    .A3(net7),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0617_));
 sky130_fd_sc_hd__mux4_1 _1711_ (.A0(net24),
    .A1(net782),
    .A2(net92),
    .A3(net120),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _1712_ (.A0(_0617_),
    .A1(_0618_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0619_));
 sky130_fd_sc_hd__a22o_4 _1713_ (.A1(_0614_),
    .A2(_0616_),
    .B1(_0619_),
    .B2(_1016_),
    .X(\Inst_RegFile_switch_matrix.JN2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1714_ (.A0(net136),
    .A1(net673),
    .A2(net659),
    .A3(net655),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_0620_));
 sky130_fd_sc_hd__mux4_1 _1715_ (.A0(net649),
    .A1(net684),
    .A2(net668),
    .A3(net637),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_2 _1716_ (.A0(_0620_),
    .A1(_0621_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .X(_0622_));
 sky130_fd_sc_hd__mux4_1 _1717_ (.A0(net86),
    .A1(net90),
    .A2(net88),
    .A3(net114),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_0623_));
 sky130_fd_sc_hd__mux4_1 _1718_ (.A0(net58),
    .A1(net1),
    .A2(net62),
    .A3(net5),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _1719_ (.A0(_0624_),
    .A1(_0623_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_4 _1720_ (.A0(_0625_),
    .A1(_0622_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.JW2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1721_ (.A0(net690),
    .A1(net652),
    .A2(net657),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0626_));
 sky130_fd_sc_hd__mux4_2 _1722_ (.A0(net680),
    .A1(net633),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_4 _1723_ (.A0(_0626_),
    .A1(_0627_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0628_));
 sky130_fd_sc_hd__mux4_1 _1724_ (.A0(net61),
    .A1(net63),
    .A2(net6),
    .A3(net781),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0629_));
 sky130_fd_sc_hd__mux4_1 _1725_ (.A0(net91),
    .A1(net107),
    .A2(net110),
    .A3(net119),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _1726_ (.A0(_0629_),
    .A1(_0630_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_4 _1727_ (.A0(_0631_),
    .A1(_0628_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_RegFile_switch_matrix.JW2BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1728_ (.A0(net693),
    .A1(net414),
    .A2(net415),
    .A3(net407),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0632_));
 sky130_fd_sc_hd__mux4_1 _1729_ (.A0(net646),
    .A1(net680),
    .A2(net665),
    .A3(net427),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_4 _1730_ (.A0(_0632_),
    .A1(_0633_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0634_));
 sky130_fd_sc_hd__mux4_1 _1731_ (.A0(net86),
    .A1(net90),
    .A2(net110),
    .A3(net114),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0635_));
 sky130_fd_sc_hd__mux4_1 _1732_ (.A0(net58),
    .A1(net1),
    .A2(net62),
    .A3(net5),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _1733_ (.A0(_0636_),
    .A1(_0635_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_4 _1734_ (.A0(_0637_),
    .A1(_0634_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.JS2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1735_ (.A0(net690),
    .A1(net652),
    .A2(net415),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0638_));
 sky130_fd_sc_hd__mux4_2 _1736_ (.A0(net680),
    .A1(net633),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_4 _1737_ (.A0(_0638_),
    .A1(_0639_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0640_));
 sky130_fd_sc_hd__mux4_1 _1738_ (.A0(net91),
    .A1(net119),
    .A2(net107),
    .A3(net136),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0641_));
 sky130_fd_sc_hd__mux4_1 _1739_ (.A0(net63),
    .A1(net6),
    .A2(net783),
    .A3(net781),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _1740_ (.A0(_0642_),
    .A1(_0641_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_4 _1741_ (.A0(_0643_),
    .A1(_0640_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ),
    .X(\Inst_RegFile_switch_matrix.JS2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1742_ (.A0(net648),
    .A1(net683),
    .A2(net431),
    .A3(net637),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_0644_));
 sky130_fd_sc_hd__mux4_1 _1743_ (.A0(net114),
    .A1(net672),
    .A2(net658),
    .A3(net419),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_0645_));
 sky130_fd_sc_hd__or2_1 _1744_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__o21a_1 _1745_ (.A1(_1017_),
    .A2(_0644_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_0647_));
 sky130_fd_sc_hd__mux4_1 _1746_ (.A0(net23),
    .A1(net88),
    .A2(net86),
    .A3(net90),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_0648_));
 sky130_fd_sc_hd__mux4_1 _1747_ (.A0(net58),
    .A1(net1),
    .A2(net62),
    .A3(net5),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _1748_ (.A0(_0648_),
    .A1(_0649_),
    .S(_1017_),
    .X(_0650_));
 sky130_fd_sc_hd__a22o_1 _1749_ (.A1(_0646_),
    .A2(_0647_),
    .B1(_0650_),
    .B2(_1018_),
    .X(\Inst_RegFile_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1750_ (.A0(net690),
    .A1(net407),
    .A2(net415),
    .A3(net647),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0651_));
 sky130_fd_sc_hd__or2_1 _1751_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__mux4_2 _1752_ (.A0(net680),
    .A1(net427),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0653_));
 sky130_fd_sc_hd__o21a_1 _1753_ (.A1(_0653_),
    .A2(_1019_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0654_));
 sky130_fd_sc_hd__mux4_1 _1754_ (.A0(net61),
    .A1(net63),
    .A2(net79),
    .A3(net82),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0655_));
 sky130_fd_sc_hd__mux4_1 _1755_ (.A0(net6),
    .A1(net91),
    .A2(net781),
    .A3(net119),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _1756_ (.A0(_0655_),
    .A1(_0656_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_0657_));
 sky130_fd_sc_hd__a22o_1 _1757_ (.A1(_0654_),
    .A2(_0652_),
    .B1(_0657_),
    .B2(_1020_),
    .X(\Inst_RegFile_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1758_ (.A0(net693),
    .A1(net673),
    .A2(net659),
    .A3(net654),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0658_));
 sky130_fd_sc_hd__mux4_1 _1759_ (.A0(net649),
    .A1(net684),
    .A2(net668),
    .A3(net637),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_4 _1760_ (.A0(_0658_),
    .A1(_0659_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_0660_));
 sky130_fd_sc_hd__nand2_4 _1761_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__mux4_1 _1762_ (.A0(net58),
    .A1(net62),
    .A2(net82),
    .A3(net1),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0662_));
 sky130_fd_sc_hd__mux4_1 _1763_ (.A0(net5),
    .A1(net90),
    .A2(net86),
    .A3(net114),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _1764_ (.A0(_0662_),
    .A1(_0663_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_0664_));
 sky130_fd_sc_hd__nand2b_1 _1765_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand2_2 _1766_ (.A(_0661_),
    .B(_0665_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1767_ (.A0(net690),
    .A1(net652),
    .A2(net415),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_0666_));
 sky130_fd_sc_hd__mux4_2 _1768_ (.A0(net680),
    .A1(net633),
    .A2(net665),
    .A3(net638),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_4 _1769_ (.A0(_0666_),
    .A1(_0667_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .X(_0668_));
 sky130_fd_sc_hd__mux4_1 _1770_ (.A0(net63),
    .A1(net79),
    .A2(net783),
    .A3(net6),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0669_));
 sky130_fd_sc_hd__mux4_1 _1771_ (.A0(net23),
    .A1(net781),
    .A2(net91),
    .A3(net119),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _1772_ (.A0(_0669_),
    .A1(_0670_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_4 _1773_ (.A0(_0671_),
    .A1(_0668_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ),
    .X(\Inst_RegFile_switch_matrix.JN2BEG0 ));
 sky130_fd_sc_hd__nand2b_1 _1774_ (.A_N(net784),
    .B(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .Y(_0672_));
 sky130_fd_sc_hd__o21ba_1 _1775_ (.A1(net84),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _1776_ (.A0(net112),
    .A1(net693),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0674_));
 sky130_fd_sc_hd__a221o_1 _1777_ (.A1(_0672_),
    .A2(_0673_),
    .B1(_0674_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _1778_ (.A0(net672),
    .A1(net659),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0676_));
 sky130_fd_sc_hd__inv_1 _1779_ (.A(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__mux2_1 _1780_ (.A0(net419),
    .A1(net649),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0678_));
 sky130_fd_sc_hd__o21ai_1 _1781_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .A2(_0677_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .Y(_0679_));
 sky130_fd_sc_hd__a21o_1 _1782_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .A2(_0678_),
    .B1(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__mux4_2 _1783_ (.A0(_0998_),
    .A1(_0983_),
    .A2(_0979_),
    .A3(_0138_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0681_));
 sky130_fd_sc_hd__inv_2 _1784_ (.A(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__mux4_2 _1785_ (.A0(net74),
    .A1(net102),
    .A2(net17),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0683_));
 sky130_fd_sc_hd__a21oi_1 _1786_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_0683_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .Y(_0684_));
 sky130_fd_sc_hd__o21a_1 _1787_ (.A1(_0681_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .B1(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__nand2_1 _1788_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .B(net403),
    .Y(_0686_));
 sky130_fd_sc_hd__o211a_1 _1789_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(net434),
    .B1(_0686_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_0687_));
 sky130_fd_sc_hd__o21ai_2 _1790_ (.A1(_0687_),
    .A2(_0685_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .Y(_0688_));
 sky130_fd_sc_hd__mux4_1 _1791_ (.A0(net683),
    .A1(net428),
    .A2(net667),
    .A3(net447),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0689_));
 sky130_fd_sc_hd__o211a_1 _1792_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .A2(_0689_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ),
    .C1(_0688_),
    .X(_0690_));
 sky130_fd_sc_hd__a31o_4 _1793_ (.A1(_1021_),
    .A2(_0675_),
    .A3(_0680_),
    .B1(_0690_),
    .X(\Inst_RegFile_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1794_ (.A0(net419),
    .A1(net648),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _1795_ (.A0(net672),
    .A1(net658),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0692_));
 sky130_fd_sc_hd__and2b_1 _1796_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .B(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__a21bo_1 _1797_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_0691_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_0694_));
 sky130_fd_sc_hd__mux4_1 _1798_ (.A0(net83),
    .A1(net4),
    .A2(net111),
    .A3(net692),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .X(_0695_));
 sky130_fd_sc_hd__o22a_1 _1799_ (.A1(_0693_),
    .A2(_0694_),
    .B1(_0695_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_0696_));
 sky130_fd_sc_hd__mux4_2 _1800_ (.A0(net73),
    .A1(net16),
    .A2(net101),
    .A3(net129),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0697_));
 sky130_fd_sc_hd__mux4_2 _1801_ (.A0(net73),
    .A1(net16),
    .A2(net101),
    .A3(net129),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _1802_ (.A0(_1044_),
    .A1(net689),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _1803_ (.A0(_0697_),
    .A1(_0698_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0700_));
 sky130_fd_sc_hd__and2b_1 _1804_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .B(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__a21bo_1 _1805_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_0699_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_0702_));
 sky130_fd_sc_hd__mux4_2 _1806_ (.A0(net683),
    .A1(net636),
    .A2(net667),
    .A3(net447),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0703_));
 sky130_fd_sc_hd__o22a_1 _1807_ (.A1(_0701_),
    .A2(_0702_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ),
    .B2(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_4 _1808_ (.A0(_0696_),
    .A1(_0704_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ),
    .X(\Inst_RegFile_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1809_ (.A0(net418),
    .A1(net87),
    .A2(net115),
    .A3(net672),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ),
    .X(_0705_));
 sky130_fd_sc_hd__mux4_2 _1810_ (.A0(net66),
    .A1(net94),
    .A2(net23),
    .A3(net122),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ),
    .X(_0706_));
 sky130_fd_sc_hd__mux4_2 _1811_ (.A0(net683),
    .A1(_1073_),
    .A2(net402),
    .A3(_0706_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_4 _1812_ (.A0(_0705_),
    .A1(_0707_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ),
    .X(\Inst_RegFile_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1813_ (.A0(net66),
    .A1(net9),
    .A2(net112),
    .A3(net122),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _1814_ (.A0(net689),
    .A1(_0708_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_0709_));
 sky130_fd_sc_hd__nand2_1 _1815_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__nor2_1 _1816_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .B(net638),
    .Y(_0711_));
 sky130_fd_sc_hd__a211o_1 _1817_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_1045_),
    .B1(_0711_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .X(_0712_));
 sky130_fd_sc_hd__and3_1 _1818_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ),
    .B(_0710_),
    .C(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__mux4_1 _1819_ (.A0(net58),
    .A1(net86),
    .A2(net114),
    .A3(net646),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .X(_0714_));
 sky130_fd_sc_hd__o21ba_1 _1820_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_0714_),
    .B1_N(_0713_),
    .X(\Inst_RegFile_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1821_ (.A0(net61),
    .A1(net89),
    .A2(net692),
    .A3(net419),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ),
    .X(_0715_));
 sky130_fd_sc_hd__mux4_2 _1822_ (.A0(net634),
    .A1(_0682_),
    .A2(_0683_),
    .A3(_0140_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_4 _1823_ (.A0(_0715_),
    .A1(_0716_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ),
    .X(\Inst_RegFile_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__o21ai_1 _1824_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0698_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ),
    .Y(_0717_));
 sky130_fd_sc_hd__a21oi_1 _1825_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0366_),
    .B1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__mux2_1 _1826_ (.A0(net667),
    .A1(_0697_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .X(_0719_));
 sky130_fd_sc_hd__inv_1 _1827_ (.A(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__o21ai_1 _1828_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ),
    .A2(_0720_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ),
    .Y(_0721_));
 sky130_fd_sc_hd__mux4_1 _1829_ (.A0(net60),
    .A1(net88),
    .A2(net693),
    .A3(net658),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ),
    .X(_0722_));
 sky130_fd_sc_hd__o22a_1 _1830_ (.A1(_0718_),
    .A2(_0721_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ),
    .B2(_0722_),
    .X(\Inst_RegFile_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1831_ (.A0(net418),
    .A1(net2),
    .A2(net115),
    .A3(net414),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .X(_0723_));
 sky130_fd_sc_hd__or2_1 _1832_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .B(net681),
    .X(_0724_));
 sky130_fd_sc_hd__a21oi_1 _1833_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(_1072_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .Y(_0725_));
 sky130_fd_sc_hd__mux4_2 _1834_ (.A0(net62),
    .A1(net90),
    .A2(net5),
    .A3(net139),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_2 _1835_ (.A0(_0352_),
    .A1(_0726_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_0727_));
 sky130_fd_sc_hd__a22o_1 _1836_ (.A1(_0724_),
    .A2(_0725_),
    .B1(_0727_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_2 _1837_ (.A0(_0723_),
    .A1(_0728_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ),
    .X(\Inst_RegFile_switch_matrix.SS4BEG3 ));
 sky130_fd_sc_hd__mux2_1 _1838_ (.A0(net689),
    .A1(_0191_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_0729_));
 sky130_fd_sc_hd__nand2_1 _1839_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__nor2_1 _1840_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .B(net640),
    .Y(_0731_));
 sky130_fd_sc_hd__a211o_1 _1841_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_1045_),
    .B1(_0731_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_0732_));
 sky130_fd_sc_hd__nor2_1 _1842_ (.A(net58),
    .B(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .Y(_0733_));
 sky130_fd_sc_hd__a211o_1 _1843_ (.A1(_1010_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .C1(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _1844_ (.A0(net114),
    .A1(net647),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_0735_));
 sky130_fd_sc_hd__a21oi_1 _1845_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .A2(_0735_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ),
    .Y(_0736_));
 sky130_fd_sc_hd__a32oi_1 _1846_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(_0730_),
    .A3(_0732_),
    .B1(_0734_),
    .B2(_0736_),
    .Y(\Inst_RegFile_switch_matrix.SS4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1847_ (.A0(net61),
    .A1(net783),
    .A2(net692),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .X(_0737_));
 sky130_fd_sc_hd__or2_1 _1848_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .B(net635),
    .X(_0738_));
 sky130_fd_sc_hd__a21oi_2 _1849_ (.A1(_0681_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .Y(_0739_));
 sky130_fd_sc_hd__mux2_4 _1850_ (.A0(_0683_),
    .A1(_0153_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .X(_0740_));
 sky130_fd_sc_hd__a22o_1 _1851_ (.A1(_0739_),
    .A2(_0738_),
    .B1(_0740_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_4 _1852_ (.A0(_0737_),
    .A1(_0741_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ),
    .X(\Inst_RegFile_switch_matrix.SS4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1853_ (.A0(_0698_),
    .A1(_0378_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .X(_0742_));
 sky130_fd_sc_hd__nand2_1 _1854_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__mux2_1 _1855_ (.A0(net666),
    .A1(_0697_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .X(_0744_));
 sky130_fd_sc_hd__inv_1 _1856_ (.A(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__o211a_1 _1857_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ),
    .A2(_0745_),
    .B1(_0743_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ),
    .X(_0746_));
 sky130_fd_sc_hd__mux4_1 _1858_ (.A0(net60),
    .A1(net3),
    .A2(net693),
    .A3(net661),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ),
    .X(_0747_));
 sky130_fd_sc_hd__o21ba_4 _1859_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ),
    .A2(_0747_),
    .B1_N(_0746_),
    .X(\Inst_RegFile_switch_matrix.SS4BEG0 ));
 sky130_fd_sc_hd__nand2b_1 _1860_ (.A_N(net784),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .Y(_0748_));
 sky130_fd_sc_hd__o21ba_1 _1861_ (.A1(net85),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _1862_ (.A0(net113),
    .A1(net693),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0750_));
 sky130_fd_sc_hd__a221o_1 _1863_ (.A1(_0748_),
    .A2(_0749_),
    .B1(_0750_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _1864_ (.A0(net674),
    .A1(net660),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0752_));
 sky130_fd_sc_hd__and2b_1 _1865_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .B(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _1866_ (.A0(net413),
    .A1(net405),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0754_));
 sky130_fd_sc_hd__a211o_1 _1867_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .A2(_0754_),
    .B1(_0753_),
    .C1(_1022_),
    .X(_0755_));
 sky130_fd_sc_hd__mux4_2 _1868_ (.A0(_0682_),
    .A1(_0683_),
    .A2(_1073_),
    .A3(net402),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .X(_0756_));
 sky130_fd_sc_hd__mux4_1 _1869_ (.A0(net684),
    .A1(net398),
    .A2(net668),
    .A3(net404),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0757_));
 sky130_fd_sc_hd__or2_1 _1870_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .B(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__o211a_1 _1871_ (.A1(_0756_),
    .A2(_1022_),
    .B1(_0758_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0759_));
 sky130_fd_sc_hd__a31o_4 _1872_ (.A1(_1023_),
    .A2(_0751_),
    .A3(_0755_),
    .B1(_0759_),
    .X(\Inst_RegFile_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1873_ (.A0(net655),
    .A1(net650),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_1 _1874_ (.A0(net674),
    .A1(net660),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0761_));
 sky130_fd_sc_hd__and2b_1 _1875_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .B(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__a21bo_1 _1876_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_0760_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_0763_));
 sky130_fd_sc_hd__mux4_1 _1877_ (.A0(net82),
    .A1(net110),
    .A2(net783),
    .A3(net692),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0764_));
 sky130_fd_sc_hd__o22a_1 _1878_ (.A1(_0762_),
    .A2(_0763_),
    .B1(_0764_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _1879_ (.A0(_1044_),
    .A1(net689),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _1880_ (.A0(_0697_),
    .A1(_0698_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0767_));
 sky130_fd_sc_hd__and2b_1 _1881_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .B(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__a21bo_1 _1882_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_0766_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_0769_));
 sky130_fd_sc_hd__mux4_1 _1883_ (.A0(net684),
    .A1(net398),
    .A2(net668),
    .A3(net642),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0770_));
 sky130_fd_sc_hd__o22a_1 _1884_ (.A1(_0768_),
    .A2(_0769_),
    .B1(_0770_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_1 _1885_ (.A0(_0765_),
    .A1(_0771_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ),
    .X(\Inst_RegFile_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1886_ (.A0(net418),
    .A1(net2),
    .A2(net87),
    .A3(net674),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0772_));
 sky130_fd_sc_hd__nor2_1 _1887_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .B(net684),
    .Y(_0773_));
 sky130_fd_sc_hd__a211oi_1 _1888_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(net434),
    .B1(_0773_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .Y(_0774_));
 sky130_fd_sc_hd__mux4_1 _1889_ (.A0(net68),
    .A1(net11),
    .A2(net113),
    .A3(net124),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _1890_ (.A0(net402),
    .A1(_0775_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .X(_0776_));
 sky130_fd_sc_hd__a21bo_1 _1891_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .A2(_0776_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ),
    .X(_0777_));
 sky130_fd_sc_hd__o22a_1 _1892_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(_0772_),
    .B1(_0774_),
    .B2(_0777_),
    .X(\Inst_RegFile_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1893_ (.A0(net85),
    .A1(net11),
    .A2(net96),
    .A3(net124),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _1894_ (.A0(net689),
    .A1(_0778_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_0779_));
 sky130_fd_sc_hd__nand2_1 _1895_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__nor2_4 _1896_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .B(net404),
    .Y(_0781_));
 sky130_fd_sc_hd__a211o_1 _1897_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(_1045_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .C1(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__nor2_1 _1898_ (.A(net58),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .Y(_0783_));
 sky130_fd_sc_hd__a211o_1 _1899_ (.A1(_1010_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .C1(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _1900_ (.A0(net86),
    .A1(net405),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_0785_));
 sky130_fd_sc_hd__a21oi_1 _1901_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .A2(_0785_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ),
    .Y(_0786_));
 sky130_fd_sc_hd__a32oi_1 _1902_ (.A1(_0782_),
    .A2(_0780_),
    .A3(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ),
    .B1(_0784_),
    .B2(_0786_),
    .Y(\Inst_RegFile_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__nor2_1 _1903_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .B(net398),
    .Y(_0787_));
 sky130_fd_sc_hd__a211oi_1 _1904_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .A2(_0681_),
    .B1(_0787_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .Y(_0788_));
 sky130_fd_sc_hd__mux2_1 _1905_ (.A0(_0683_),
    .A1(_0559_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .X(_0789_));
 sky130_fd_sc_hd__mux4_1 _1906_ (.A0(net61),
    .A1(net783),
    .A2(net89),
    .A3(net413),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .X(_0790_));
 sky130_fd_sc_hd__a21bo_1 _1907_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .A2(_0789_),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ),
    .X(_0791_));
 sky130_fd_sc_hd__o22a_4 _1908_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ),
    .A2(_0790_),
    .B1(_0791_),
    .B2(_0788_),
    .X(\Inst_RegFile_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1909_ (.A0(_0698_),
    .A1(_0541_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .X(_0792_));
 sky130_fd_sc_hd__nand2_1 _1910_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__mux2_1 _1911_ (.A0(net668),
    .A1(_0697_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .X(_0794_));
 sky130_fd_sc_hd__inv_1 _1912_ (.A(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__o211a_1 _1913_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .A2(_0795_),
    .B1(_0793_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _1914_ (.A0(net60),
    .A1(net784),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .X(_0797_));
 sky130_fd_sc_hd__nand2b_1 _1915_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__mux2_2 _1916_ (.A0(net88),
    .A1(net660),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .X(_0799_));
 sky130_fd_sc_hd__a21oi_2 _1917_ (.A1(_0799_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ),
    .Y(_0800_));
 sky130_fd_sc_hd__a21oi_1 _1918_ (.A1(_0798_),
    .A2(_0800_),
    .B1(_0796_),
    .Y(\Inst_RegFile_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1919_ (.A0(net418),
    .A1(net2),
    .A2(net115),
    .A3(net673),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0801_));
 sky130_fd_sc_hd__or2_1 _1920_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .B(net683),
    .X(_0802_));
 sky130_fd_sc_hd__a21oi_1 _1921_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_1072_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ),
    .Y(_0803_));
 sky130_fd_sc_hd__mux4_2 _1922_ (.A0(net82),
    .A1(net92),
    .A2(net7),
    .A3(net120),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_2 _1923_ (.A0(net402),
    .A1(_0804_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_0805_));
 sky130_fd_sc_hd__a22o_1 _1924_ (.A1(_0802_),
    .A2(_0803_),
    .B1(_0805_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _1925_ (.A0(_0801_),
    .A1(_0806_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.NN4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1926_ (.A0(net64),
    .A1(net92),
    .A2(net7),
    .A3(net138),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _1927_ (.A0(net689),
    .A1(_0807_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_0808_));
 sky130_fd_sc_hd__nand2_1 _1928_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .B(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__nor2_1 _1929_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .B(net404),
    .Y(_0810_));
 sky130_fd_sc_hd__a211o_1 _1930_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_1045_),
    .B1(_0810_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_0811_));
 sky130_fd_sc_hd__nor2_1 _1931_ (.A(net58),
    .B(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .Y(_0812_));
 sky130_fd_sc_hd__a211o_1 _1932_ (.A1(_1010_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .C1(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _1933_ (.A0(net114),
    .A1(net648),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_0814_));
 sky130_fd_sc_hd__a21oi_1 _1934_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .A2(_0814_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ),
    .Y(_0815_));
 sky130_fd_sc_hd__a32oi_1 _1935_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ),
    .A2(_0809_),
    .A3(_0811_),
    .B1(_0813_),
    .B2(_0815_),
    .Y(\Inst_RegFile_switch_matrix.NN4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1936_ (.A0(net61),
    .A1(net783),
    .A2(net692),
    .A3(net413),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .X(_0816_));
 sky130_fd_sc_hd__or2_1 _1937_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .B(net398),
    .X(_0817_));
 sky130_fd_sc_hd__a21oi_2 _1938_ (.A1(_0681_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .Y(_0818_));
 sky130_fd_sc_hd__mux2_2 _1939_ (.A0(_0683_),
    .A1(_1060_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .X(_0819_));
 sky130_fd_sc_hd__a22o_1 _1940_ (.A1(_0818_),
    .A2(_0817_),
    .B1(_0819_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_4 _1941_ (.A0(_0816_),
    .A1(_0820_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ),
    .X(\Inst_RegFile_switch_matrix.NN4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1942_ (.A0(_0698_),
    .A1(_0341_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .X(_0821_));
 sky130_fd_sc_hd__nand2_1 _1943_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ),
    .B(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__mux2_1 _1944_ (.A0(net668),
    .A1(_0697_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .X(_0823_));
 sky130_fd_sc_hd__inv_1 _1945_ (.A(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__o211a_1 _1946_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ),
    .A2(_0824_),
    .B1(_0822_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ),
    .X(_0825_));
 sky130_fd_sc_hd__mux4_2 _1947_ (.A0(net60),
    .A1(net784),
    .A2(net693),
    .A3(net660),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ),
    .X(_0826_));
 sky130_fd_sc_hd__o21ba_4 _1948_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(_0826_),
    .B1_N(_0825_),
    .X(\Inst_RegFile_switch_matrix.NN4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1949_ (.A0(net85),
    .A1(net109),
    .A2(net136),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_0827_));
 sky130_fd_sc_hd__mux4_2 _1950_ (.A0(net414),
    .A1(_0407_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .A3(_0827_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1951_ (.A0(net638),
    .A1(net689),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .A3(_0377_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1952_ (.A0(net427),
    .A1(_0563_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .A3(net396),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1953_ (.A0(net80),
    .A1(net125),
    .A2(net7),
    .A3(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_0828_));
 sky130_fd_sc_hd__mux4_2 _1954_ (.A0(net71),
    .A1(net14),
    .A2(net99),
    .A3(net127),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ),
    .X(_0829_));
 sky130_fd_sc_hd__mux4_2 _1955_ (.A0(net406),
    .A1(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .A2(_0829_),
    .A3(_0828_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1956_ (.A0(net91),
    .A1(net691),
    .A2(net106),
    .A3(net647),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1957_ (.A0(net90),
    .A1(net690),
    .A2(net109),
    .A3(net653),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1958_ (.A0(net782),
    .A1(net93),
    .A2(net108),
    .A3(net661),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1959_ (.A0(net781),
    .A1(net107),
    .A2(net92),
    .A3(net671),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1960_ (.A0(net640),
    .A1(_0407_),
    .A2(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .A3(_0827_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1961_ (.A0(net635),
    .A1(net689),
    .A2(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .A3(_0377_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1962_ (.A0(net666),
    .A1(_0563_),
    .A2(\Inst_RegFile_switch_matrix.E2BEG0 ),
    .A3(net396),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1963_ (.A0(net682),
    .A1(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .A2(_0829_),
    .A3(_0828_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1964_ (.A0(net635),
    .A1(_0407_),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .A3(_0827_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1965_ (.A0(net406),
    .A1(net689),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .A3(_0377_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1966_ (.A0(net682),
    .A1(_0563_),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .A3(net396),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1967_ (.A0(net647),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .A2(_0829_),
    .A3(_0828_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1968_ (.A0(net63),
    .A1(net78),
    .A2(net691),
    .A3(net639),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1969_ (.A0(net62),
    .A1(net690),
    .A2(net81),
    .A3(net428),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1970_ (.A0(net65),
    .A1(net80),
    .A2(net782),
    .A3(net667),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1971_ (.A0(net64),
    .A1(net79),
    .A2(net781),
    .A3(net681),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1972_ (.A0(net667),
    .A1(_0407_),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .A3(_0827_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1973_ (.A0(net680),
    .A1(net689),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .A3(_0377_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1974_ (.A0(net646),
    .A1(_0563_),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .A3(net396),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1975_ (.A0(net407),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .A2(_0829_),
    .A3(_0828_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__a21o_1 _1976_ (.A1(_0661_),
    .A2(_0665_),
    .B1(_1028_),
    .X(_0830_));
 sky130_fd_sc_hd__a21oi_1 _1977_ (.A1(_1028_),
    .A2(_0726_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .Y(_0831_));
 sky130_fd_sc_hd__mux2_1 _1978_ (.A0(\Inst_RegFile_switch_matrix.JW2BEG7 ),
    .A1(\Inst_RegFile_switch_matrix.JS2BEG7 ),
    .S(_1028_),
    .X(_0832_));
 sky130_fd_sc_hd__a2bb2o_1 _1979_ (.A1_N(_1029_),
    .A2_N(_0832_),
    .B1(_0831_),
    .B2(_0830_),
    .X(_0833_));
 sky130_fd_sc_hd__a211o_1 _1980_ (.A1(_1039_),
    .A2(_1040_),
    .B1(_1042_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0834_));
 sky130_fd_sc_hd__o211a_1 _1981_ (.A1(_1028_),
    .A2(_0128_),
    .B1(_0834_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _1982_ (.A0(net62),
    .A1(net90),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0836_));
 sky130_fd_sc_hd__a21o_1 _1983_ (.A1(_1029_),
    .A2(_0836_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0837_));
 sky130_fd_sc_hd__a2bb2o_4 _1984_ (.A1_N(_0835_),
    .A2_N(_0837_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ),
    .B2(_0833_),
    .X(_0838_));
 sky130_fd_sc_hd__o21ai_1 _1985_ (.A1(_0991_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ),
    .Y(_0839_));
 sky130_fd_sc_hd__a21o_1 _1986_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .B1(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _1987_ (.A0(net78),
    .A1(net110),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0841_));
 sky130_fd_sc_hd__o21a_1 _1988_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ),
    .A2(_0841_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0842_));
 sky130_fd_sc_hd__a22o_1 _1989_ (.A1(_1027_),
    .A2(_0191_),
    .B1(_0840_),
    .B2(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__mux4_2 _1990_ (.A0(net70),
    .A1(net126),
    .A2(net98),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_4 _1991_ (.A0(_0829_),
    .A1(_0844_),
    .S(_1027_),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_4 _1992_ (.A0(_0845_),
    .A1(_0843_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ),
    .X(_0846_));
 sky130_fd_sc_hd__and2b_2 _1993_ (.A_N(_0838_),
    .B(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__mux4_2 _1994_ (.A0(net75),
    .A1(net18),
    .A2(net103),
    .A3(net131),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_4 _1995_ (.A0(_0683_),
    .A1(_0848_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0849_));
 sky130_fd_sc_hd__and2b_1 _1996_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .B(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__mux4_1 _1997_ (.A0(net83),
    .A1(net24),
    .A2(net107),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_2 _1998_ (.A0(_0708_),
    .A1(_0851_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0852_));
 sky130_fd_sc_hd__a21oi_4 _1999_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .A2(_0852_),
    .B1(_0850_),
    .Y(_0853_));
 sky130_fd_sc_hd__a21o_4 _2000_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .A2(_0852_),
    .B1(_0850_),
    .X(_0854_));
 sky130_fd_sc_hd__nand2_8 _2001_ (.A(net437),
    .B(_0847_),
    .Y(_0855_));
 sky130_fd_sc_hd__mux2_1 _2002_ (.A0(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .A1(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .S(_1030_),
    .X(_0856_));
 sky130_fd_sc_hd__a21o_1 _2003_ (.A1(_1030_),
    .A2(_0378_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ),
    .X(_0857_));
 sky130_fd_sc_hd__a21o_1 _2004_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .B1(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__o21ai_1 _2005_ (.A1(_1031_),
    .A2(_0856_),
    .B1(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__mux4_1 _2006_ (.A0(_0970_),
    .A1(_0974_),
    .A2(_0989_),
    .A3(net435),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0860_));
 sky130_fd_sc_hd__nor2_1 _2007_ (.A(_1030_),
    .B(_0848_),
    .Y(_0861_));
 sky130_fd_sc_hd__a211o_1 _2008_ (.A1(_1030_),
    .A2(_0860_),
    .B1(_0861_),
    .C1(_1031_),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _2009_ (.A0(net65),
    .A1(net93),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .X(_0863_));
 sky130_fd_sc_hd__a21oi_1 _2010_ (.A1(_1031_),
    .A2(_0863_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_0864_));
 sky130_fd_sc_hd__a22o_1 _2011_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ),
    .A2(_0859_),
    .B1(_0862_),
    .B2(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__mux4_2 _2012_ (.A0(net8),
    .A1(net113),
    .A2(net138),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ),
    .X(_0866_));
 sky130_fd_sc_hd__mux2_4 _2013_ (.A0(_0778_),
    .A1(_0866_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _2014_ (.A0(net132),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _2015_ (.A0(net19),
    .A1(net104),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_0869_));
 sky130_fd_sc_hd__and2b_1 _2016_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ),
    .B(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__a211o_1 _2017_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ),
    .A2(_0868_),
    .B1(_0870_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _2018_ (.A0(net77),
    .A1(net20),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0872_));
 sky130_fd_sc_hd__inv_1 _2019_ (.A(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__mux2_1 _2020_ (.A0(net105),
    .A1(net133),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_1 _2021_ (.A(\Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__o211a_1 _2022_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ),
    .A2(_0873_),
    .B1(_0875_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0876_));
 sky130_fd_sc_hd__nor2_1 _2023_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ),
    .B(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__a22o_4 _2024_ (.A1(_0867_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ),
    .B1(_0871_),
    .B2(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__or2_4 _2025_ (.A(_0878_),
    .B(_0865_),
    .X(_0879_));
 sky130_fd_sc_hd__or2_1 _2026_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .B(_0860_),
    .X(_0880_));
 sky130_fd_sc_hd__a21oi_2 _2027_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0698_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .Y(_0881_));
 sky130_fd_sc_hd__nand2_1 _2028_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .B(_0828_),
    .Y(_0882_));
 sky130_fd_sc_hd__nand2b_1 _2029_ (.A_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .B(_0807_),
    .Y(_0883_));
 sky130_fd_sc_hd__a32oi_4 _2030_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0882_),
    .A3(_0883_),
    .B1(_0880_),
    .B2(_0881_),
    .Y(_0884_));
 sky130_fd_sc_hd__a32o_1 _2031_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0882_),
    .A3(_0883_),
    .B1(_0880_),
    .B2(_0881_),
    .X(_0885_));
 sky130_fd_sc_hd__nor2_8 _2032_ (.A(_0884_),
    .B(_0879_),
    .Y(_0886_));
 sky130_fd_sc_hd__or2_4 _2033_ (.A(_0884_),
    .B(_0879_),
    .X(_0887_));
 sky130_fd_sc_hd__nor2_8 _2034_ (.A(_0887_),
    .B(_0855_),
    .Y(_0888_));
 sky130_fd_sc_hd__mux2_4 _2035_ (.A0(_0775_),
    .A1(_0827_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .X(_0889_));
 sky130_fd_sc_hd__mux4_1 _2036_ (.A0(net76),
    .A1(net104),
    .A2(net132),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _2037_ (.A0(net77),
    .A1(net20),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0891_));
 sky130_fd_sc_hd__or2_1 _2038_ (.A(\Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ),
    .B(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_1 _2039_ (.A0(net105),
    .A1(net133),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_0893_));
 sky130_fd_sc_hd__o211a_1 _2040_ (.A1(_1025_),
    .A2(_0893_),
    .B1(_0892_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .X(_0894_));
 sky130_fd_sc_hd__a21o_1 _2041_ (.A1(_1026_),
    .A2(_0890_),
    .B1(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_2 _2042_ (.A0(_0895_),
    .A1(_0889_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_4 _2043_ (.A0(net471),
    .A1(net610),
    .S(_0888_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _2044_ (.A0(_0406_),
    .A1(_0697_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_0897_));
 sky130_fd_sc_hd__mux4_1 _2045_ (.A0(net25),
    .A1(net125),
    .A2(net108),
    .A3(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _2046_ (.A0(_0804_),
    .A1(_0898_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_2 _2047_ (.A0(_0897_),
    .A1(_0899_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_4 _2048_ (.A0(net507),
    .A1(net606),
    .S(_0888_),
    .X(_0001_));
 sky130_fd_sc_hd__mux4_2 _2049_ (.A0(net79),
    .A1(net690),
    .A2(net781),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_0901_));
 sky130_fd_sc_hd__mux4_2 _2050_ (.A0(_0682_),
    .A1(_0706_),
    .A2(_0407_),
    .A3(_0901_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_4 _2051_ (.A0(net485),
    .A1(net631),
    .S(_0888_),
    .X(_0002_));
 sky130_fd_sc_hd__nand2_1 _2052_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .B(_0598_),
    .Y(_0903_));
 sky130_fd_sc_hd__o211a_1 _2053_ (.A1(net106),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ),
    .C1(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _2054_ (.A0(net78),
    .A1(net782),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0905_));
 sky130_fd_sc_hd__inv_1 _2055_ (.A(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__o21ai_1 _2056_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_0906_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .Y(_0907_));
 sky130_fd_sc_hd__o221a_1 _2057_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0726_),
    .B1(_0904_),
    .B2(_0907_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _2058_ (.A0(net98),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_0909_));
 sky130_fd_sc_hd__nand2_1 _2059_ (.A(_0986_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .Y(_0910_));
 sky130_fd_sc_hd__o21ba_1 _2060_ (.A1(net70),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .B1_N(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_0911_));
 sky130_fd_sc_hd__a221o_1 _2061_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ),
    .A2(_0909_),
    .B1(_0910_),
    .B2(_0911_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _2062_ (.A0(net71),
    .A1(net14),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0913_));
 sky130_fd_sc_hd__inv_1 _2063_ (.A(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__mux2_1 _2064_ (.A0(net99),
    .A1(net127),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0915_));
 sky130_fd_sc_hd__o21ai_1 _2065_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_0914_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .Y(_0916_));
 sky130_fd_sc_hd__a21o_1 _2066_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_0915_),
    .B1(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__a31o_2 _2067_ (.A1(_1024_),
    .A2(_0912_),
    .A3(_0917_),
    .B1(_0908_),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_4 _2068_ (.A0(net536),
    .A1(net602),
    .S(_0888_),
    .X(_0003_));
 sky130_fd_sc_hd__nand2b_1 _2069_ (.A_N(_0865_),
    .B(_0878_),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_4 _2070_ (.A(_0884_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__or2_4 _2071_ (.A(_0884_),
    .B(_0919_),
    .X(_0921_));
 sky130_fd_sc_hd__nor2_8 _2072_ (.A(_0921_),
    .B(_0855_),
    .Y(_0922_));
 sky130_fd_sc_hd__mux2_4 _2073_ (.A0(net532),
    .A1(net610),
    .S(_0922_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_4 _2074_ (.A0(net551),
    .A1(net606),
    .S(_0922_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_4 _2075_ (.A0(net564),
    .A1(net631),
    .S(_0922_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_4 _2076_ (.A0(net571),
    .A1(net602),
    .S(_0922_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_8 _2077_ (.A(_0885_),
    .B(_0879_),
    .Y(_0923_));
 sky130_fd_sc_hd__or2_4 _2078_ (.A(_0885_),
    .B(_0879_),
    .X(_0924_));
 sky130_fd_sc_hd__nor2_8 _2079_ (.A(_0924_),
    .B(_0855_),
    .Y(_0925_));
 sky130_fd_sc_hd__mux2_4 _2080_ (.A0(net469),
    .A1(net610),
    .S(_0925_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_4 _2081_ (.A0(net484),
    .A1(net606),
    .S(_0925_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_4 _2082_ (.A0(net472),
    .A1(net631),
    .S(_0925_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_4 _2083_ (.A0(net489),
    .A1(net602),
    .S(_0925_),
    .X(_0011_));
 sky130_fd_sc_hd__nor2_2 _2084_ (.A(_0885_),
    .B(_0919_),
    .Y(_0926_));
 sky130_fd_sc_hd__or2_4 _2085_ (.A(_0885_),
    .B(_0919_),
    .X(_0927_));
 sky130_fd_sc_hd__nor2_8 _2086_ (.A(_0927_),
    .B(_0855_),
    .Y(_0928_));
 sky130_fd_sc_hd__mux2_4 _2087_ (.A0(net556),
    .A1(net610),
    .S(_0928_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_4 _2088_ (.A0(net539),
    .A1(net606),
    .S(_0928_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_4 _2089_ (.A0(net550),
    .A1(net631),
    .S(_0928_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_4 _2090_ (.A0(net572),
    .A1(net602),
    .S(_0928_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_4 _2091_ (.A(_0847_),
    .B(_0854_),
    .X(_0929_));
 sky130_fd_sc_hd__nand2_8 _2092_ (.A(_0854_),
    .B(_0847_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2_8 _2093_ (.A(_0886_),
    .B(_0929_),
    .Y(_0931_));
 sky130_fd_sc_hd__mux2_4 _2094_ (.A0(net609),
    .A1(net488),
    .S(_0931_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_4 _2095_ (.A0(net604),
    .A1(net483),
    .S(_0931_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_4 _2096_ (.A0(net630),
    .A1(net475),
    .S(_0931_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_4 _2097_ (.A0(net600),
    .A1(net522),
    .S(_0931_),
    .X(_0019_));
 sky130_fd_sc_hd__nand2b_4 _2098_ (.A_N(_0846_),
    .B(_0838_),
    .Y(_0932_));
 sky130_fd_sc_hd__nor2_8 _2099_ (.A(_0932_),
    .B(_0854_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand2_8 _2100_ (.A(_0923_),
    .B(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__mux2_4 _2101_ (.A0(net611),
    .A1(net502),
    .S(_0934_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_4 _2102_ (.A0(net605),
    .A1(net482),
    .S(_0934_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_4 _2103_ (.A0(net629),
    .A1(net513),
    .S(_0934_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_4 _2104_ (.A0(net601),
    .A1(net462),
    .S(_0934_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_8 _2105_ (.A(_0930_),
    .B(_0924_),
    .Y(_0935_));
 sky130_fd_sc_hd__mux2_4 _2106_ (.A0(net559),
    .A1(net609),
    .S(_0935_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_4 _2107_ (.A0(net506),
    .A1(net606),
    .S(_0935_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_4 _2108_ (.A0(net464),
    .A1(net630),
    .S(_0935_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_4 _2109_ (.A0(net493),
    .A1(net602),
    .S(_0935_),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_4 _2110_ (.A(_0838_),
    .B(_0846_),
    .Y(_0936_));
 sky130_fd_sc_hd__nor2_8 _2111_ (.A(_0936_),
    .B(_0854_),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_8 _2112_ (.A(_0920_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__mux2_4 _2113_ (.A0(net609),
    .A1(net562),
    .S(_0938_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_4 _2114_ (.A0(net605),
    .A1(net549),
    .S(_0938_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_4 _2115_ (.A0(net629),
    .A1(net494),
    .S(_0938_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_4 _2116_ (.A0(net601),
    .A1(net526),
    .S(_0938_),
    .X(_0031_));
 sky130_fd_sc_hd__nor2_8 _2117_ (.A(_0936_),
    .B(net437),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_8 _2118_ (.A(_0920_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__mux2_4 _2119_ (.A0(net608),
    .A1(net568),
    .S(_0940_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_4 _2120_ (.A0(net604),
    .A1(net576),
    .S(_0940_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_4 _2121_ (.A0(net630),
    .A1(net546),
    .S(_0940_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_4 _2122_ (.A0(net600),
    .A1(net567),
    .S(_0940_),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_8 _2123_ (.A(_0838_),
    .B(_0846_),
    .Y(_0941_));
 sky130_fd_sc_hd__nand2_8 _2124_ (.A(_0941_),
    .B(net437),
    .Y(_0942_));
 sky130_fd_sc_hd__nor2_8 _2125_ (.A(_0942_),
    .B(_0921_),
    .Y(_0943_));
 sky130_fd_sc_hd__mux2_4 _2126_ (.A0(net560),
    .A1(net610),
    .S(_0943_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_4 _2127_ (.A0(net528),
    .A1(net606),
    .S(_0943_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_4 _2128_ (.A0(net565),
    .A1(net631),
    .S(_0943_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_4 _2129_ (.A0(net575),
    .A1(net602),
    .S(_0943_),
    .X(_0039_));
 sky130_fd_sc_hd__nand2_8 _2130_ (.A(_0941_),
    .B(_0854_),
    .Y(_0944_));
 sky130_fd_sc_hd__nor2_8 _2131_ (.A(_0944_),
    .B(_0924_),
    .Y(_0945_));
 sky130_fd_sc_hd__mux2_4 _2132_ (.A0(net519),
    .A1(net611),
    .S(_0945_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_4 _2133_ (.A0(net458),
    .A1(net607),
    .S(_0945_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_4 _2134_ (.A0(net542),
    .A1(net632),
    .S(_0945_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_4 _2135_ (.A0(net541),
    .A1(net603),
    .S(_0945_),
    .X(_0043_));
 sky130_fd_sc_hd__nor2_8 _2136_ (.A(_0927_),
    .B(_0944_),
    .Y(_0946_));
 sky130_fd_sc_hd__mux2_4 _2137_ (.A0(net573),
    .A1(net611),
    .S(_0946_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_2 _2138_ (.A0(net511),
    .A1(net607),
    .S(_0946_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_4 _2139_ (.A0(net577),
    .A1(net632),
    .S(_0946_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_4 _2140_ (.A0(net574),
    .A1(net603),
    .S(_0946_),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_8 _2141_ (.A(_0939_),
    .B(_0923_),
    .Y(_0947_));
 sky130_fd_sc_hd__mux2_4 _2142_ (.A0(net608),
    .A1(net478),
    .S(_0947_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_4 _2143_ (.A0(net604),
    .A1(net534),
    .S(_0947_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_4 _2144_ (.A0(net629),
    .A1(net455),
    .S(_0947_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_4 _2145_ (.A0(net600),
    .A1(net514),
    .S(_0947_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_8 _2146_ (.A(_0926_),
    .B(_0939_),
    .Y(_0948_));
 sky130_fd_sc_hd__mux2_4 _2147_ (.A0(net608),
    .A1(net516),
    .S(_0948_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_4 _2148_ (.A0(net604),
    .A1(net558),
    .S(_0948_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_4 _2149_ (.A0(net629),
    .A1(net579),
    .S(_0948_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_4 _2150_ (.A0(net600),
    .A1(net529),
    .S(_0948_),
    .X(_0055_));
 sky130_fd_sc_hd__nor2_8 _2151_ (.A(_0942_),
    .B(_0887_),
    .Y(_0949_));
 sky130_fd_sc_hd__mux2_4 _2152_ (.A0(net480),
    .A1(net610),
    .S(_0949_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_4 _2153_ (.A0(net487),
    .A1(net606),
    .S(_0949_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_4 _2154_ (.A0(net474),
    .A1(net631),
    .S(_0949_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_4 _2155_ (.A0(net554),
    .A1(net602),
    .S(_0949_),
    .X(_0059_));
 sky130_fd_sc_hd__nor2_8 _2156_ (.A(_0942_),
    .B(_0924_),
    .Y(_0950_));
 sky130_fd_sc_hd__mux2_4 _2157_ (.A0(net459),
    .A1(net610),
    .S(_0950_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_4 _2158_ (.A0(net463),
    .A1(net606),
    .S(_0950_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_4 _2159_ (.A0(net466),
    .A1(net631),
    .S(_0950_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_4 _2160_ (.A0(net457),
    .A1(net602),
    .S(_0950_),
    .X(_0063_));
 sky130_fd_sc_hd__nand2_4 _2161_ (.A(_0920_),
    .B(_0933_),
    .Y(_0951_));
 sky130_fd_sc_hd__mux2_4 _2162_ (.A0(net609),
    .A1(net524),
    .S(_0951_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_2 _2163_ (.A0(net605),
    .A1(net518),
    .S(_0951_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_4 _2164_ (.A0(net629),
    .A1(net517),
    .S(_0951_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_2 _2165_ (.A0(net601),
    .A1(net530),
    .S(_0951_),
    .X(_0067_));
 sky130_fd_sc_hd__nor2_8 _2166_ (.A(_0944_),
    .B(_0887_),
    .Y(_0952_));
 sky130_fd_sc_hd__mux2_4 _2167_ (.A0(net452),
    .A1(net610),
    .S(_0952_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_4 _2168_ (.A0(net473),
    .A1(net607),
    .S(_0952_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_4 _2169_ (.A0(net499),
    .A1(net631),
    .S(_0952_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_4 _2170_ (.A0(net495),
    .A1(net603),
    .S(_0952_),
    .X(_0071_));
 sky130_fd_sc_hd__nor2_8 _2171_ (.A(_0944_),
    .B(_0921_),
    .Y(_0953_));
 sky130_fd_sc_hd__mux2_4 _2172_ (.A0(net537),
    .A1(net610),
    .S(_0953_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_4 _2173_ (.A0(net578),
    .A1(net607),
    .S(_0953_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_4 _2174_ (.A0(net561),
    .A1(net631),
    .S(_0953_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_4 _2175_ (.A0(net566),
    .A1(net603),
    .S(_0953_),
    .X(_0075_));
 sky130_fd_sc_hd__nor2_8 _2176_ (.A(_0942_),
    .B(_0927_),
    .Y(_0954_));
 sky130_fd_sc_hd__mux2_4 _2177_ (.A0(net548),
    .A1(net610),
    .S(_0954_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_4 _2178_ (.A0(net555),
    .A1(net606),
    .S(_0954_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_4 _2179_ (.A0(net545),
    .A1(net631),
    .S(_0954_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_4 _2180_ (.A0(net569),
    .A1(net602),
    .S(_0954_),
    .X(_0079_));
 sky130_fd_sc_hd__nand2_8 _2181_ (.A(_0920_),
    .B(_0929_),
    .Y(_0955_));
 sky130_fd_sc_hd__mux2_4 _2182_ (.A0(net609),
    .A1(net557),
    .S(_0955_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_4 _2183_ (.A0(net604),
    .A1(net553),
    .S(_0955_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_4 _2184_ (.A0(net630),
    .A1(net540),
    .S(_0955_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_4 _2185_ (.A0(net600),
    .A1(net563),
    .S(_0955_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_8 _2186_ (.A(_0927_),
    .B(_0930_),
    .Y(_0956_));
 sky130_fd_sc_hd__mux2_2 _2187_ (.A0(net523),
    .A1(net609),
    .S(_0956_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_4 _2188_ (.A0(net544),
    .A1(net606),
    .S(_0956_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_2 _2189_ (.A0(net501),
    .A1(net632),
    .S(_0956_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_2 _2190_ (.A0(net531),
    .A1(net602),
    .S(_0956_),
    .X(_0087_));
 sky130_fd_sc_hd__nand2_4 _2191_ (.A(_0926_),
    .B(_0933_),
    .Y(_0957_));
 sky130_fd_sc_hd__mux2_2 _2192_ (.A0(net609),
    .A1(net503),
    .S(_0957_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_4 _2193_ (.A0(net605),
    .A1(net515),
    .S(_0957_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_4 _2194_ (.A0(net629),
    .A1(net527),
    .S(_0957_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_2 _2195_ (.A0(net601),
    .A1(net461),
    .S(_0957_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_8 _2196_ (.A(_0932_),
    .B(net437),
    .Y(_0958_));
 sky130_fd_sc_hd__nand2_8 _2197_ (.A(_0958_),
    .B(_0886_),
    .Y(_0959_));
 sky130_fd_sc_hd__mux2_4 _2198_ (.A0(net608),
    .A1(net490),
    .S(_0959_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_4 _2199_ (.A0(net604),
    .A1(net521),
    .S(_0959_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_4 _2200_ (.A0(net630),
    .A1(net453),
    .S(_0959_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_4 _2201_ (.A0(net600),
    .A1(net456),
    .S(_0959_),
    .X(_0095_));
 sky130_fd_sc_hd__nand2_8 _2202_ (.A(_0920_),
    .B(_0958_),
    .Y(_0960_));
 sky130_fd_sc_hd__mux2_4 _2203_ (.A0(net608),
    .A1(net504),
    .S(_0960_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_4 _2204_ (.A0(net604),
    .A1(net533),
    .S(_0960_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_4 _2205_ (.A0(net630),
    .A1(net497),
    .S(_0960_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_4 _2206_ (.A0(net600),
    .A1(net505),
    .S(_0960_),
    .X(_0099_));
 sky130_fd_sc_hd__nand2_8 _2207_ (.A(_0923_),
    .B(net439),
    .Y(_0961_));
 sky130_fd_sc_hd__mux2_4 _2208_ (.A0(net608),
    .A1(net525),
    .S(_0961_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_4 _2209_ (.A0(net604),
    .A1(net538),
    .S(_0961_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_4 _2210_ (.A0(net630),
    .A1(net460),
    .S(_0961_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_4 _2211_ (.A0(net600),
    .A1(net500),
    .S(_0961_),
    .X(_0103_));
 sky130_fd_sc_hd__nand2_8 _2212_ (.A(_0926_),
    .B(_0958_),
    .Y(_0962_));
 sky130_fd_sc_hd__mux2_4 _2213_ (.A0(net608),
    .A1(net492),
    .S(_0962_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_4 _2214_ (.A0(net604),
    .A1(net509),
    .S(_0962_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_4 _2215_ (.A0(net630),
    .A1(net491),
    .S(_0962_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_4 _2216_ (.A0(net600),
    .A1(net535),
    .S(_0962_),
    .X(_0107_));
 sky130_fd_sc_hd__nand2_8 _2217_ (.A(_0886_),
    .B(_0937_),
    .Y(_0963_));
 sky130_fd_sc_hd__mux2_4 _2218_ (.A0(net609),
    .A1(net477),
    .S(_0963_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_4 _2219_ (.A0(net605),
    .A1(net512),
    .S(_0963_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_4 _2220_ (.A0(net629),
    .A1(net467),
    .S(_0963_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_4 _2221_ (.A0(net601),
    .A1(net481),
    .S(_0963_),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_8 _2222_ (.A(_0933_),
    .B(_0886_),
    .Y(_0964_));
 sky130_fd_sc_hd__mux2_4 _2223_ (.A0(net609),
    .A1(net476),
    .S(_0964_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_4 _2224_ (.A0(net605),
    .A1(net520),
    .S(_0964_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_4 _2225_ (.A0(net629),
    .A1(net498),
    .S(_0964_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_4 _2226_ (.A0(net601),
    .A1(net486),
    .S(_0964_),
    .X(_0115_));
 sky130_fd_sc_hd__nand2_8 _2227_ (.A(_0923_),
    .B(_0937_),
    .Y(_0965_));
 sky130_fd_sc_hd__mux2_4 _2228_ (.A0(net608),
    .A1(net470),
    .S(_0965_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_4 _2229_ (.A0(net605),
    .A1(net552),
    .S(_0965_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_4 _2230_ (.A0(net629),
    .A1(net465),
    .S(_0965_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_4 _2231_ (.A0(net601),
    .A1(net468),
    .S(_0965_),
    .X(_0119_));
 sky130_fd_sc_hd__nand2_8 _2232_ (.A(_0926_),
    .B(_0937_),
    .Y(_0966_));
 sky130_fd_sc_hd__mux2_4 _2233_ (.A0(net608),
    .A1(net510),
    .S(_0966_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_4 _2234_ (.A0(net605),
    .A1(net547),
    .S(_0966_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_4 _2235_ (.A0(net629),
    .A1(net508),
    .S(_0966_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_4 _2236_ (.A0(net601),
    .A1(net570),
    .S(_0966_),
    .X(_0123_));
 sky130_fd_sc_hd__nand2_4 _2237_ (.A(_0939_),
    .B(_0886_),
    .Y(_0967_));
 sky130_fd_sc_hd__mux2_2 _2238_ (.A0(net608),
    .A1(net479),
    .S(_0967_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_4 _2239_ (.A0(net604),
    .A1(net543),
    .S(_0967_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_2 _2240_ (.A0(net630),
    .A1(net454),
    .S(_0967_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_2 _2241_ (.A0(net600),
    .A1(net496),
    .S(_0967_),
    .X(_0127_));
 sky130_fd_sc_hd__dfxtp_1 _2242_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0000_),
    .Q(\Inst_RegFile_32x4.mem[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2243_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0001_),
    .Q(\Inst_RegFile_32x4.mem[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2244_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0002_),
    .Q(\Inst_RegFile_32x4.mem[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2245_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0003_),
    .Q(\Inst_RegFile_32x4.mem[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2246_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0004_),
    .Q(\Inst_RegFile_32x4.mem[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2247_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0005_),
    .Q(\Inst_RegFile_32x4.mem[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2248_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0006_),
    .Q(\Inst_RegFile_32x4.mem[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2249_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0007_),
    .Q(\Inst_RegFile_32x4.mem[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2250_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0008_),
    .Q(\Inst_RegFile_32x4.mem[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2251_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0009_),
    .Q(\Inst_RegFile_32x4.mem[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2252_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0010_),
    .Q(\Inst_RegFile_32x4.mem[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2253_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0011_),
    .Q(\Inst_RegFile_32x4.mem[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2254_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0012_),
    .Q(\Inst_RegFile_32x4.mem[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2255_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0013_),
    .Q(\Inst_RegFile_32x4.mem[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2256_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0014_),
    .Q(\Inst_RegFile_32x4.mem[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2257_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0015_),
    .Q(\Inst_RegFile_32x4.mem[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2258_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0016_),
    .Q(\Inst_RegFile_32x4.mem[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2259_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0017_),
    .Q(\Inst_RegFile_32x4.mem[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2260_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0018_),
    .Q(\Inst_RegFile_32x4.mem[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2261_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0019_),
    .Q(\Inst_RegFile_32x4.mem[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2262_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0020_),
    .Q(\Inst_RegFile_32x4.mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2263_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0021_),
    .Q(\Inst_RegFile_32x4.mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2264_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0022_),
    .Q(\Inst_RegFile_32x4.mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2265_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0023_),
    .Q(\Inst_RegFile_32x4.mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2266_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0024_),
    .Q(\Inst_RegFile_32x4.mem[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2267_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0025_),
    .Q(\Inst_RegFile_32x4.mem[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2268_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0026_),
    .Q(\Inst_RegFile_32x4.mem[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2269_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0027_),
    .Q(\Inst_RegFile_32x4.mem[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2270_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0028_),
    .Q(\Inst_RegFile_32x4.mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2271_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0029_),
    .Q(\Inst_RegFile_32x4.mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2272_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0030_),
    .Q(\Inst_RegFile_32x4.mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2273_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0031_),
    .Q(\Inst_RegFile_32x4.mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2274_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0032_),
    .Q(\Inst_RegFile_32x4.mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2275_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0033_),
    .Q(\Inst_RegFile_32x4.mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2276_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0034_),
    .Q(\Inst_RegFile_32x4.mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2277_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0035_),
    .Q(\Inst_RegFile_32x4.mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2278_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0036_),
    .Q(\Inst_RegFile_32x4.mem[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2279_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0037_),
    .Q(\Inst_RegFile_32x4.mem[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2280_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0038_),
    .Q(\Inst_RegFile_32x4.mem[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2281_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0039_),
    .Q(\Inst_RegFile_32x4.mem[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2282_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0040_),
    .Q(\Inst_RegFile_32x4.mem[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2283_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0041_),
    .Q(\Inst_RegFile_32x4.mem[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2284_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0042_),
    .Q(\Inst_RegFile_32x4.mem[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2285_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0043_),
    .Q(\Inst_RegFile_32x4.mem[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2286_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0044_),
    .Q(\Inst_RegFile_32x4.mem[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2287_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0045_),
    .Q(\Inst_RegFile_32x4.mem[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2288_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0046_),
    .Q(\Inst_RegFile_32x4.mem[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2289_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0047_),
    .Q(\Inst_RegFile_32x4.mem[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2290_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0048_),
    .Q(\Inst_RegFile_32x4.mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2291_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0049_),
    .Q(\Inst_RegFile_32x4.mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2292_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0050_),
    .Q(\Inst_RegFile_32x4.mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2293_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0051_),
    .Q(\Inst_RegFile_32x4.mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2294_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0052_),
    .Q(\Inst_RegFile_32x4.mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2295_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0053_),
    .Q(\Inst_RegFile_32x4.mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2296_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0054_),
    .Q(\Inst_RegFile_32x4.mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2297_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0055_),
    .Q(\Inst_RegFile_32x4.mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2298_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0056_),
    .Q(\Inst_RegFile_32x4.mem[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2299_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0057_),
    .Q(\Inst_RegFile_32x4.mem[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2300_ (.CLK(clknet_4_14_0_UserCLK_regs),
    .D(_0058_),
    .Q(\Inst_RegFile_32x4.mem[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2301_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0059_),
    .Q(\Inst_RegFile_32x4.mem[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2302_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0060_),
    .Q(\Inst_RegFile_32x4.mem[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2303_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0061_),
    .Q(\Inst_RegFile_32x4.mem[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2304_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0062_),
    .Q(\Inst_RegFile_32x4.mem[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2305_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0063_),
    .Q(\Inst_RegFile_32x4.mem[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2306_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0064_),
    .Q(\Inst_RegFile_32x4.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2307_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0065_),
    .Q(\Inst_RegFile_32x4.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2308_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0066_),
    .Q(\Inst_RegFile_32x4.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2309_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0067_),
    .Q(\Inst_RegFile_32x4.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2310_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0068_),
    .Q(\Inst_RegFile_32x4.mem[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2311_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0069_),
    .Q(\Inst_RegFile_32x4.mem[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2312_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0070_),
    .Q(\Inst_RegFile_32x4.mem[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2313_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0071_),
    .Q(\Inst_RegFile_32x4.mem[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2314_ (.CLK(clknet_4_10_0_UserCLK_regs),
    .D(_0072_),
    .Q(\Inst_RegFile_32x4.mem[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2315_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0073_),
    .Q(\Inst_RegFile_32x4.mem[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2316_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0074_),
    .Q(\Inst_RegFile_32x4.mem[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2317_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(_0075_),
    .Q(\Inst_RegFile_32x4.mem[21][3] ));
 sky130_fd_sc_hd__dlxtp_1 _2318_ (.D(net757),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2319_ (.D(net754),
    .GATE(net734),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2320_ (.D(net753),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2321_ (.D(net752),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2322_ (.D(net751),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2323_ (.D(net749),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2324_ (.D(net748),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2325_ (.D(net747),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2326_ (.D(net779),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2327_ (.D(net778),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2328_ (.D(net777),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2329_ (.D(net776),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2330_ (.D(net775),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2331_ (.D(net774),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2332_ (.D(net773),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2333_ (.D(net772),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2334_ (.D(net771),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2335_ (.D(net770),
    .GATE(net733),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2336_ (.D(net39),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2337_ (.D(net40),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2338_ (.D(net766),
    .GATE(net732),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2339_ (.D(net42),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2340_ (.D(net43),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2341_ (.D(net44),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2342_ (.D(net761),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2343_ (.D(net760),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2344_ (.D(net759),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2345_ (.D(net758),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2346_ (.D(net756),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2347_ (.D(net50),
    .GATE(net731),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2348_ (.D(net780),
    .GATE(net57),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2349_ (.D(net769),
    .GATE(net57),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2350_ (.D(net757),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2351_ (.D(net754),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2352_ (.D(net753),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2353_ (.D(net752),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2354_ (.D(net54),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2355_ (.D(net750),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2356_ (.D(net748),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2357_ (.D(net56),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2358_ (.D(net779),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2359_ (.D(net29),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2360_ (.D(net30),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2361_ (.D(net31),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2362_ (.D(net32),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2363_ (.D(net33),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2364_ (.D(net773),
    .GATE(net738),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2365_ (.D(net772),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2366_ (.D(net771),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2367_ (.D(net770),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2368_ (.D(net768),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2369_ (.D(net767),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2370_ (.D(net766),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2371_ (.D(net765),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2372_ (.D(net764),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2373_ (.D(net763),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2374_ (.D(net761),
    .GATE(net736),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2375_ (.D(net760),
    .GATE(net737),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2376_ (.D(net759),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2377_ (.D(net758),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2378_ (.D(net756),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2379_ (.D(net755),
    .GATE(net735),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2380_ (.D(net780),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2381_ (.D(net38),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2382_ (.D(net48),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2383_ (.D(net51),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2384_ (.D(net52),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2385_ (.D(net53),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2386_ (.D(net54),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2387_ (.D(net750),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2388_ (.D(net55),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2389_ (.D(net56),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2390_ (.D(net779),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2391_ (.D(net778),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2392_ (.D(net30),
    .GATE(net742),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2393_ (.D(net31),
    .GATE(net742),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2394_ (.D(net32),
    .GATE(net742),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2395_ (.D(net33),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2396_ (.D(net773),
    .GATE(net741),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2397_ (.D(net35),
    .GATE(net742),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2398_ (.D(net36),
    .GATE(net742),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2399_ (.D(net37),
    .GATE(net742),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2400_ (.D(net768),
    .GATE(net742),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2401_ (.D(net767),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2402_ (.D(net766),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2403_ (.D(net765),
    .GATE(net740),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2404_ (.D(net764),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2405_ (.D(net763),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2406_ (.D(net762),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2407_ (.D(net760),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2408_ (.D(net759),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2409_ (.D(net758),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2410_ (.D(net756),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2411_ (.D(net755),
    .GATE(net739),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2412_ (.D(net780),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2413_ (.D(net769),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2414_ (.D(net757),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2415_ (.D(net754),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2416_ (.D(net753),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2417_ (.D(net752),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2418_ (.D(net751),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2419_ (.D(net749),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2420_ (.D(net748),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2421_ (.D(net747),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2422_ (.D(net779),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2423_ (.D(net778),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2424_ (.D(net777),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2425_ (.D(net776),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2426_ (.D(net775),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2427_ (.D(net774),
    .GATE(net694),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2428_ (.D(net773),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2429_ (.D(net772),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2430_ (.D(net771),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2431_ (.D(net770),
    .GATE(net695),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2432_ (.D(net768),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2433_ (.D(net767),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2434_ (.D(net766),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2435_ (.D(net765),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2436_ (.D(net764),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2437_ (.D(net763),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2438_ (.D(net762),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2439_ (.D(net760),
    .GATE(net696),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2440_ (.D(net46),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2441_ (.D(net47),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2442_ (.D(net756),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2443_ (.D(net755),
    .GATE(net697),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2444_ (.D(net780),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2445_ (.D(net769),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2446_ (.D(net757),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2447_ (.D(net754),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2448_ (.D(net52),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2449_ (.D(net53),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2450_ (.D(net751),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2451_ (.D(net750),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2452_ (.D(net748),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2453_ (.D(net747),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2454_ (.D(net28),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2455_ (.D(net778),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2456_ (.D(net777),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2457_ (.D(net776),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2458_ (.D(net775),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2459_ (.D(net774),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2460_ (.D(net773),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2461_ (.D(net772),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2462_ (.D(net36),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2463_ (.D(net770),
    .GATE(net699),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2464_ (.D(net768),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2465_ (.D(net40),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2466_ (.D(net766),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2467_ (.D(net765),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2468_ (.D(net764),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2469_ (.D(net763),
    .GATE(net700),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2470_ (.D(net761),
    .GATE(net701),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2471_ (.D(net760),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2472_ (.D(net46),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2473_ (.D(net758),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2474_ (.D(net756),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2475_ (.D(net755),
    .GATE(net698),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2476_ (.D(net27),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2477_ (.D(net38),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2478_ (.D(net48),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2479_ (.D(net51),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2480_ (.D(net52),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2481_ (.D(net53),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2482_ (.D(net751),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2483_ (.D(net749),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2484_ (.D(net748),
    .GATE(net705),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2485_ (.D(net747),
    .GATE(net705),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2486_ (.D(net28),
    .GATE(net706),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2487_ (.D(net29),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2488_ (.D(net777),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2489_ (.D(net776),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2490_ (.D(net775),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2491_ (.D(net774),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2492_ (.D(net34),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2493_ (.D(net35),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2494_ (.D(net771),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2495_ (.D(net37),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2496_ (.D(net768),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2497_ (.D(net767),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2498_ (.D(net766),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2499_ (.D(net765),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2500_ (.D(net764),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2501_ (.D(net763),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2502_ (.D(net761),
    .GATE(net705),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2503_ (.D(net760),
    .GATE(net703),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2504_ (.D(net46),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2505_ (.D(net47),
    .GATE(net704),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2506_ (.D(net756),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2507_ (.D(net755),
    .GATE(net702),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2508_ (.D(net780),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2509_ (.D(net769),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2510_ (.D(net757),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2511_ (.D(net754),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2512_ (.D(net753),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2513_ (.D(net752),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2514_ (.D(net751),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2515_ (.D(net749),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2516_ (.D(net55),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2517_ (.D(net747),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2518_ (.D(net779),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2519_ (.D(net778),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2520_ (.D(net30),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2521_ (.D(net31),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2522_ (.D(net32),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2523_ (.D(net33),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2524_ (.D(net34),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2525_ (.D(net772),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2526_ (.D(net771),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2527_ (.D(net770),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2528_ (.D(net768),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2529_ (.D(net767),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2530_ (.D(net766),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2531_ (.D(net765),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2532_ (.D(net764),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2533_ (.D(net763),
    .GATE(net710),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2534_ (.D(net762),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2535_ (.D(net760),
    .GATE(net707),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2536_ (.D(net759),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2537_ (.D(net758),
    .GATE(net709),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2538_ (.D(net756),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2539_ (.D(net755),
    .GATE(net708),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2540_ (.D(net27),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2541_ (.D(net769),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2542_ (.D(net48),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2543_ (.D(net51),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2544_ (.D(net753),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2545_ (.D(net752),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2546_ (.D(net751),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2547_ (.D(net749),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2548_ (.D(net748),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2549_ (.D(net747),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2550_ (.D(net28),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2551_ (.D(net29),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2552_ (.D(net777),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2553_ (.D(net776),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2554_ (.D(net775),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2555_ (.D(net774),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2556_ (.D(net34),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2557_ (.D(net35),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2558_ (.D(net36),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2559_ (.D(net37),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2560_ (.D(net768),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2561_ (.D(net767),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2562_ (.D(net766),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2563_ (.D(net765),
    .GATE(net712),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2564_ (.D(net43),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2565_ (.D(net44),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2566_ (.D(net762),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2567_ (.D(net45),
    .GATE(net714),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2568_ (.D(net759),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2569_ (.D(net758),
    .GATE(net713),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2570_ (.D(net756),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2571_ (.D(net755),
    .GATE(net711),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2572_ (.D(net780),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2573_ (.D(net769),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2574_ (.D(net757),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2575_ (.D(net754),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2576_ (.D(net753),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2577_ (.D(net752),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2578_ (.D(net751),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2579_ (.D(net749),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2580_ (.D(net748),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2581_ (.D(net747),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2582_ (.D(net779),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2583_ (.D(net778),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2584_ (.D(net777),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2585_ (.D(net776),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2586_ (.D(net775),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2587_ (.D(net774),
    .GATE(net715),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2588_ (.D(net773),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2589_ (.D(net772),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2590_ (.D(net771),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2591_ (.D(net770),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2592_ (.D(net39),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2593_ (.D(net40),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2594_ (.D(net41),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2595_ (.D(net42),
    .GATE(net718),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2596_ (.D(net764),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2597_ (.D(net763),
    .GATE(net716),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2598_ (.D(net761),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2599_ (.D(net45),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2600_ (.D(net759),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2601_ (.D(net758),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2602_ (.D(net49),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2603_ (.D(net50),
    .GATE(net717),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2604_ (.D(net780),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2605_ (.D(net769),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2606_ (.D(net757),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2607_ (.D(net754),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2608_ (.D(net753),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2609_ (.D(net752),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2610_ (.D(net54),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2611_ (.D(net749),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2612_ (.D(net748),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2613_ (.D(net747),
    .GATE(net719),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2614_ (.D(net779),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2615_ (.D(net778),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2616_ (.D(net777),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2617_ (.D(net776),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2618_ (.D(net775),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2619_ (.D(net774),
    .GATE(net720),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2620_ (.D(net773),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2621_ (.D(net772),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2622_ (.D(net771),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2623_ (.D(net770),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2624_ (.D(net39),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2625_ (.D(net40),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2626_ (.D(net766),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2627_ (.D(net765),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2628_ (.D(net43),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2629_ (.D(net763),
    .GATE(net722),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2630_ (.D(net761),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2631_ (.D(net760),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2632_ (.D(net759),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2633_ (.D(net758),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2634_ (.D(net49),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2635_ (.D(net50),
    .GATE(net721),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2636_ (.D(net780),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2637_ (.D(net769),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2638_ (.D(net757),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2639_ (.D(net754),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2640_ (.D(net753),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2641_ (.D(net752),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2642_ (.D(net751),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2643_ (.D(net749),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2644_ (.D(net748),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2645_ (.D(net747),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2646_ (.D(net779),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2647_ (.D(net778),
    .GATE(net726),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2648_ (.D(net777),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2649_ (.D(net776),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2650_ (.D(net775),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2651_ (.D(net774),
    .GATE(net724),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2652_ (.D(net773),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2653_ (.D(net772),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2654_ (.D(net771),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2655_ (.D(net770),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2656_ (.D(net768),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2657_ (.D(net767),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2658_ (.D(net41),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2659_ (.D(net42),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2660_ (.D(net43),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2661_ (.D(net44),
    .GATE(net725),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2662_ (.D(net761),
    .GATE(net726),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2663_ (.D(net45),
    .GATE(net726),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2664_ (.D(net759),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2665_ (.D(net758),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2666_ (.D(net756),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2667_ (.D(net755),
    .GATE(net723),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2668_ (.D(net780),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2669_ (.D(net769),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2670_ (.D(net757),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2671_ (.D(net754),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2672_ (.D(net753),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2673_ (.D(net752),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2674_ (.D(net751),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2675_ (.D(net749),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2676_ (.D(net748),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2677_ (.D(net747),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2678_ (.D(net779),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2679_ (.D(net778),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2680_ (.D(net777),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2681_ (.D(net776),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2682_ (.D(net775),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2683_ (.D(net774),
    .GATE(net730),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2684_ (.D(net773),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2685_ (.D(net772),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2686_ (.D(net771),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2687_ (.D(net770),
    .GATE(net727),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2688_ (.D(net768),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2689_ (.D(net767),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2690_ (.D(net41),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2691_ (.D(net42),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2692_ (.D(net764),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2693_ (.D(net763),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2694_ (.D(net761),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2695_ (.D(net45),
    .GATE(net728),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2696_ (.D(net759),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2697_ (.D(net758),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2698_ (.D(net49),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2699_ (.D(net50),
    .GATE(net729),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2700_ (.D(net780),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2701_ (.D(net769),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2702_ (.D(net48),
    .GATE(net744),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2703_ (.D(net51),
    .GATE(net744),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2704_ (.D(net753),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2705_ (.D(net752),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2706_ (.D(net751),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2707_ (.D(net749),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2708_ (.D(net55),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2709_ (.D(net56),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2710_ (.D(net28),
    .GATE(net744),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2711_ (.D(net29),
    .GATE(net744),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2712_ (.D(net30),
    .GATE(net746),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2713_ (.D(net31),
    .GATE(net744),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2714_ (.D(net775),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2715_ (.D(net774),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2716_ (.D(net34),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2717_ (.D(net35),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2718_ (.D(net36),
    .GATE(net744),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2719_ (.D(net37),
    .GATE(net744),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2720_ (.D(net768),
    .GATE(net746),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2721_ (.D(net767),
    .GATE(net746),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2722_ (.D(net766),
    .GATE(net744),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2723_ (.D(net765),
    .GATE(net744),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2724_ (.D(net764),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2725_ (.D(net44),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2726_ (.D(net761),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2727_ (.D(net760),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2728_ (.D(net759),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2729_ (.D(net47),
    .GATE(net745),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2730_ (.D(net756),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2731_ (.D(net755),
    .GATE(net743),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dfxtp_1 _2732_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.BD_comb[0] ),
    .Q(\Inst_RegFile_32x4.BD_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2733_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.BD_comb[1] ),
    .Q(\Inst_RegFile_32x4.BD_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2734_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.BD_comb[2] ),
    .Q(\Inst_RegFile_32x4.BD_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2735_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.BD_comb[3] ),
    .Q(\Inst_RegFile_32x4.BD_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2736_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.AD_comb[0] ),
    .Q(\Inst_RegFile_32x4.AD_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2737_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.AD_comb[1] ),
    .Q(\Inst_RegFile_32x4.AD_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2738_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.AD_comb[2] ),
    .Q(\Inst_RegFile_32x4.AD_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2739_ (.CLK(clknet_4_8_0_UserCLK_regs),
    .D(\Inst_RegFile_32x4.AD_comb[3] ),
    .Q(\Inst_RegFile_32x4.AD_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2740_ (.CLK(clknet_4_11_0_UserCLK_regs),
    .D(_0076_),
    .Q(\Inst_RegFile_32x4.mem[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2741_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0077_),
    .Q(\Inst_RegFile_32x4.mem[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2742_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0078_),
    .Q(\Inst_RegFile_32x4.mem[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2743_ (.CLK(clknet_4_15_0_UserCLK_regs),
    .D(_0079_),
    .Q(\Inst_RegFile_32x4.mem[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2744_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0080_),
    .Q(\Inst_RegFile_32x4.mem[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2745_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0081_),
    .Q(\Inst_RegFile_32x4.mem[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2746_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0082_),
    .Q(\Inst_RegFile_32x4.mem[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2747_ (.CLK(clknet_4_9_0_UserCLK_regs),
    .D(_0083_),
    .Q(\Inst_RegFile_32x4.mem[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2748_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0084_),
    .Q(\Inst_RegFile_32x4.mem[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2749_ (.CLK(clknet_4_13_0_UserCLK_regs),
    .D(_0085_),
    .Q(\Inst_RegFile_32x4.mem[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2750_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0086_),
    .Q(\Inst_RegFile_32x4.mem[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2751_ (.CLK(clknet_4_12_0_UserCLK_regs),
    .D(_0087_),
    .Q(\Inst_RegFile_32x4.mem[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2752_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0088_),
    .Q(\Inst_RegFile_32x4.mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2753_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0089_),
    .Q(\Inst_RegFile_32x4.mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2754_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0090_),
    .Q(\Inst_RegFile_32x4.mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2755_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0091_),
    .Q(\Inst_RegFile_32x4.mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2756_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0092_),
    .Q(\Inst_RegFile_32x4.mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2757_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0093_),
    .Q(\Inst_RegFile_32x4.mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2758_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0094_),
    .Q(\Inst_RegFile_32x4.mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2759_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0095_),
    .Q(\Inst_RegFile_32x4.mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2760_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0096_),
    .Q(\Inst_RegFile_32x4.mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2761_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0097_),
    .Q(\Inst_RegFile_32x4.mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2762_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0098_),
    .Q(\Inst_RegFile_32x4.mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2763_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0099_),
    .Q(\Inst_RegFile_32x4.mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2764_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0100_),
    .Q(\Inst_RegFile_32x4.mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2765_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0101_),
    .Q(\Inst_RegFile_32x4.mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2766_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0102_),
    .Q(\Inst_RegFile_32x4.mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2767_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0103_),
    .Q(\Inst_RegFile_32x4.mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2768_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0104_),
    .Q(\Inst_RegFile_32x4.mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2769_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0105_),
    .Q(\Inst_RegFile_32x4.mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2770_ (.CLK(clknet_4_0_0_UserCLK_regs),
    .D(_0106_),
    .Q(\Inst_RegFile_32x4.mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2771_ (.CLK(clknet_4_2_0_UserCLK_regs),
    .D(_0107_),
    .Q(\Inst_RegFile_32x4.mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2772_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0108_),
    .Q(\Inst_RegFile_32x4.mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2773_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0109_),
    .Q(\Inst_RegFile_32x4.mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2774_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0110_),
    .Q(\Inst_RegFile_32x4.mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2775_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0111_),
    .Q(\Inst_RegFile_32x4.mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2776_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0112_),
    .Q(\Inst_RegFile_32x4.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2777_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0113_),
    .Q(\Inst_RegFile_32x4.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2778_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0114_),
    .Q(\Inst_RegFile_32x4.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2779_ (.CLK(clknet_4_6_0_UserCLK_regs),
    .D(_0115_),
    .Q(\Inst_RegFile_32x4.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2780_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0116_),
    .Q(\Inst_RegFile_32x4.mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2781_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0117_),
    .Q(\Inst_RegFile_32x4.mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2782_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0118_),
    .Q(\Inst_RegFile_32x4.mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2783_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0119_),
    .Q(\Inst_RegFile_32x4.mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2784_ (.CLK(clknet_4_4_0_UserCLK_regs),
    .D(_0120_),
    .Q(\Inst_RegFile_32x4.mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2785_ (.CLK(clknet_4_7_0_UserCLK_regs),
    .D(_0121_),
    .Q(\Inst_RegFile_32x4.mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2786_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0122_),
    .Q(\Inst_RegFile_32x4.mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2787_ (.CLK(clknet_4_5_0_UserCLK_regs),
    .D(_0123_),
    .Q(\Inst_RegFile_32x4.mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2788_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0124_),
    .Q(\Inst_RegFile_32x4.mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2789_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0125_),
    .Q(\Inst_RegFile_32x4.mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2790_ (.CLK(clknet_4_1_0_UserCLK_regs),
    .D(_0126_),
    .Q(\Inst_RegFile_32x4.mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2791_ (.CLK(clknet_4_3_0_UserCLK_regs),
    .D(_0127_),
    .Q(\Inst_RegFile_32x4.mem[12][3] ));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(net433),
    .X(net434));
 sky130_fd_sc_hd__buf_6 _2793_ (.A(\Inst_RegFile_switch_matrix.E1BEG1 ),
    .X(net141));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer11 (.A(net402),
    .X(net403));
 sky130_fd_sc_hd__buf_6 rebuffer41 (.A(_1072_),
    .X(net433));
 sky130_fd_sc_hd__buf_6 _2796_ (.A(\Inst_RegFile_switch_matrix.E2BEG0 ),
    .X(net144));
 sky130_fd_sc_hd__buf_6 _2797_ (.A(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .X(net145));
 sky130_fd_sc_hd__buf_6 _2798_ (.A(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .X(net146));
 sky130_fd_sc_hd__buf_1 _2799_ (.A(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .X(net147));
 sky130_fd_sc_hd__buf_6 rebuffer43 (.A(_0334_),
    .X(net435));
 sky130_fd_sc_hd__buf_1 _2801_ (.A(\Inst_RegFile_switch_matrix.E2BEG5 ),
    .X(net149));
 sky130_fd_sc_hd__buf_12 rebuffer45 (.A(_0853_),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 _2803_ (.A(\Inst_RegFile_switch_matrix.E2BEG7 ),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 _2804_ (.A(net13),
    .X(net152));
 sky130_fd_sc_hd__buf_1 _2805_ (.A(net14),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 _2806_ (.A(net15),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 _2807_ (.A(net16),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 _2808_ (.A(net17),
    .X(net156));
 sky130_fd_sc_hd__buf_1 _2809_ (.A(net18),
    .X(net157));
 sky130_fd_sc_hd__buf_1 _2810_ (.A(net19),
    .X(net158));
 sky130_fd_sc_hd__buf_1 _2811_ (.A(net20),
    .X(net159));
 sky130_fd_sc_hd__buf_1 _2812_ (.A(E6END[2]),
    .X(net160));
 sky130_fd_sc_hd__buf_1 _2813_ (.A(E6END[3]),
    .X(net163));
 sky130_fd_sc_hd__buf_1 _2814_ (.A(E6END[4]),
    .X(net164));
 sky130_fd_sc_hd__buf_1 _2815_ (.A(E6END[5]),
    .X(net165));
 sky130_fd_sc_hd__buf_1 _2816_ (.A(E6END[6]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 _2817_ (.A(E6END[7]),
    .X(net167));
 sky130_fd_sc_hd__buf_1 _2818_ (.A(E6END[8]),
    .X(net168));
 sky130_fd_sc_hd__buf_1 _2819_ (.A(E6END[9]),
    .X(net169));
 sky130_fd_sc_hd__buf_1 _2820_ (.A(E6END[10]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 _2821_ (.A(E6END[11]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 _2822_ (.A(\Inst_RegFile_switch_matrix.E6BEG0 ),
    .X(net161));
 sky130_fd_sc_hd__mux2_4 clone3 (.A0(_0564_),
    .A1(_0561_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ),
    .X(net395));
 sky130_fd_sc_hd__buf_1 _2824_ (.A(EE4END[4]),
    .X(net172));
 sky130_fd_sc_hd__buf_1 _2825_ (.A(EE4END[5]),
    .X(net179));
 sky130_fd_sc_hd__buf_1 _2826_ (.A(EE4END[6]),
    .X(net180));
 sky130_fd_sc_hd__buf_1 _2827_ (.A(EE4END[7]),
    .X(net181));
 sky130_fd_sc_hd__buf_1 _2828_ (.A(EE4END[8]),
    .X(net182));
 sky130_fd_sc_hd__buf_1 _2829_ (.A(EE4END[9]),
    .X(net183));
 sky130_fd_sc_hd__buf_1 _2830_ (.A(EE4END[10]),
    .X(net184));
 sky130_fd_sc_hd__buf_1 _2831_ (.A(EE4END[11]),
    .X(net185));
 sky130_fd_sc_hd__buf_1 _2832_ (.A(EE4END[12]),
    .X(net186));
 sky130_fd_sc_hd__buf_1 _2833_ (.A(EE4END[13]),
    .X(net187));
 sky130_fd_sc_hd__buf_1 _2834_ (.A(EE4END[14]),
    .X(net173));
 sky130_fd_sc_hd__buf_1 _2835_ (.A(EE4END[15]),
    .X(net174));
 sky130_fd_sc_hd__buf_4 _2836_ (.A(\Inst_RegFile_switch_matrix.EE4BEG0 ),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 clone54 (.A(net679),
    .X(net446));
 sky130_fd_sc_hd__buf_4 _2838_ (.A(\Inst_RegFile_switch_matrix.EE4BEG2 ),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 _2839_ (.A(\Inst_RegFile_switch_matrix.EE4BEG3 ),
    .X(net178));
 sky130_fd_sc_hd__buf_1 _2840_ (.A(net27),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 _2841_ (.A(net38),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 _2842_ (.A(net757),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 _2843_ (.A(net754),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 _2844_ (.A(net52),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 _2845_ (.A(net53),
    .X(net215));
 sky130_fd_sc_hd__buf_4 _2846_ (.A(net54),
    .X(net216));
 sky130_fd_sc_hd__buf_4 _2847_ (.A(net750),
    .X(net217));
 sky130_fd_sc_hd__buf_1 _2848_ (.A(net55),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 _2849_ (.A(net56),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 _2850_ (.A(net779),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 _2851_ (.A(net778),
    .X(net190));
 sky130_fd_sc_hd__buf_4 _2852_ (.A(net777),
    .X(net191));
 sky130_fd_sc_hd__buf_4 _2853_ (.A(net776),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 _2854_ (.A(net32),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 _2855_ (.A(net33),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 _2856_ (.A(net773),
    .X(net195));
 sky130_fd_sc_hd__buf_1 _2857_ (.A(net772),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 _2858_ (.A(net771),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 _2859_ (.A(net770),
    .X(net198));
 sky130_fd_sc_hd__buf_1 _2860_ (.A(net39),
    .X(net200));
 sky130_fd_sc_hd__buf_1 _2861_ (.A(net767),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 _2862_ (.A(net41),
    .X(net202));
 sky130_fd_sc_hd__buf_1 _2863_ (.A(net765),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 _2864_ (.A(net764),
    .X(net204));
 sky130_fd_sc_hd__buf_4 _2865_ (.A(net763),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 _2866_ (.A(net761),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 _2867_ (.A(net760),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 _2868_ (.A(net46),
    .X(net208));
 sky130_fd_sc_hd__buf_1 _2869_ (.A(net47),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 _2870_ (.A(net49),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 _2871_ (.A(net755),
    .X(net212));
 sky130_fd_sc_hd__buf_2 _2872_ (.A(net746),
    .X(net220));
 sky130_fd_sc_hd__buf_2 _2873_ (.A(net730),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 _2874_ (.A(net726),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 _2875_ (.A(net722),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 _2876_ (.A(net718),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 _2877_ (.A(net714),
    .X(net235));
 sky130_fd_sc_hd__buf_1 _2878_ (.A(net710),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 _2879_ (.A(net705),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 _2880_ (.A(net701),
    .X(net238));
 sky130_fd_sc_hd__buf_1 _2881_ (.A(net697),
    .X(net239));
 sky130_fd_sc_hd__buf_4 _2882_ (.A(FrameStrobe[10]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 _2883_ (.A(net738),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 _2884_ (.A(net734),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 _2885_ (.A(FrameStrobe[13]),
    .X(net224));
 sky130_fd_sc_hd__buf_1 _2886_ (.A(FrameStrobe[14]),
    .X(net225));
 sky130_fd_sc_hd__buf_1 _2887_ (.A(FrameStrobe[15]),
    .X(net226));
 sky130_fd_sc_hd__buf_1 _2888_ (.A(FrameStrobe[16]),
    .X(net227));
 sky130_fd_sc_hd__buf_1 _2889_ (.A(FrameStrobe[17]),
    .X(net228));
 sky130_fd_sc_hd__buf_1 _2890_ (.A(FrameStrobe[18]),
    .X(net229));
 sky130_fd_sc_hd__buf_1 _2891_ (.A(FrameStrobe[19]),
    .X(net230));
 sky130_fd_sc_hd__buf_6 _2892_ (.A(\Inst_RegFile_switch_matrix.N1BEG0 ),
    .X(net240));
 sky130_fd_sc_hd__buf_6 _2893_ (.A(\Inst_RegFile_switch_matrix.N1BEG1 ),
    .X(net241));
 sky130_fd_sc_hd__buf_6 _2894_ (.A(\Inst_RegFile_switch_matrix.N1BEG2 ),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 clone40 (.A(net625),
    .X(net432));
 sky130_fd_sc_hd__buf_8 _2896_ (.A(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .X(net244));
 sky130_fd_sc_hd__buf_8 _2897_ (.A(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .X(net245));
 sky130_fd_sc_hd__buf_6 _2898_ (.A(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 _2899_ (.A(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .X(net247));
 sky130_fd_sc_hd__buf_6 _2900_ (.A(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .X(net248));
 sky130_fd_sc_hd__buf_1 _2901_ (.A(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .X(net249));
 sky130_fd_sc_hd__buf_8 clone52 (.A(net677),
    .X(net444));
 sky130_fd_sc_hd__buf_6 _2903_ (.A(\Inst_RegFile_switch_matrix.JN2BEG7 ),
    .X(net251));
 sky130_fd_sc_hd__buf_4 _2904_ (.A(net70),
    .X(net252));
 sky130_fd_sc_hd__buf_4 _2905_ (.A(net71),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 _2906_ (.A(net72),
    .X(net254));
 sky130_fd_sc_hd__buf_1 _2907_ (.A(net73),
    .X(net255));
 sky130_fd_sc_hd__buf_1 _2908_ (.A(net74),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 _2909_ (.A(net75),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 _2910_ (.A(net76),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 _2911_ (.A(net77),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 _2912_ (.A(N4END[4]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 _2913_ (.A(N4END[5]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 _2914_ (.A(N4END[6]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 _2915_ (.A(N4END[7]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 _2916_ (.A(N4END[8]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 _2917_ (.A(N4END[9]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 _2918_ (.A(N4END[10]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 _2919_ (.A(N4END[11]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 _2920_ (.A(N4END[12]),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 _2921_ (.A(N4END[13]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 _2922_ (.A(N4END[14]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 _2923_ (.A(N4END[15]),
    .X(net262));
 sky130_fd_sc_hd__buf_6 _2924_ (.A(\Inst_RegFile_switch_matrix.N4BEG0 ),
    .X(net263));
 sky130_fd_sc_hd__buf_1 _2925_ (.A(\Inst_RegFile_switch_matrix.N4BEG1 ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\Inst_RegFile_32x4.mem[4][3] ),
    .X(net456));
 sky130_fd_sc_hd__buf_4 _2927_ (.A(\Inst_RegFile_switch_matrix.N4BEG3 ),
    .X(net266));
 sky130_fd_sc_hd__buf_1 _2928_ (.A(NN4END[4]),
    .X(net276));
 sky130_fd_sc_hd__buf_1 _2929_ (.A(NN4END[5]),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 _2930_ (.A(NN4END[6]),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 _2931_ (.A(NN4END[7]),
    .X(net285));
 sky130_fd_sc_hd__buf_1 _2932_ (.A(NN4END[8]),
    .X(net286));
 sky130_fd_sc_hd__buf_1 _2933_ (.A(NN4END[9]),
    .X(net287));
 sky130_fd_sc_hd__buf_1 _2934_ (.A(NN4END[10]),
    .X(net288));
 sky130_fd_sc_hd__buf_1 _2935_ (.A(NN4END[11]),
    .X(net289));
 sky130_fd_sc_hd__buf_1 _2936_ (.A(NN4END[12]),
    .X(net290));
 sky130_fd_sc_hd__buf_1 _2937_ (.A(NN4END[13]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_2 _2938_ (.A(NN4END[14]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 _2939_ (.A(NN4END[15]),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\Inst_RegFile_32x4.mem[12][2] ),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 clone55 (.A(net642),
    .X(net447));
 sky130_fd_sc_hd__buf_4 _2942_ (.A(\Inst_RegFile_switch_matrix.NN4BEG2 ),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 _2943_ (.A(\Inst_RegFile_switch_matrix.NN4BEG3 ),
    .X(net282));
 sky130_fd_sc_hd__buf_6 _2944_ (.A(\Inst_RegFile_switch_matrix.S1BEG0 ),
    .X(net292));
 sky130_fd_sc_hd__buf_8 clone36 (.A(net637),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(_0352_),
    .X(net402));
 sky130_fd_sc_hd__buf_6 clone35 (.A(net635),
    .X(net427));
 sky130_fd_sc_hd__buf_6 _2948_ (.A(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 _2949_ (.A(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .X(net297));
 sky130_fd_sc_hd__buf_6 _2950_ (.A(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .X(net298));
 sky130_fd_sc_hd__buf_6 _2951_ (.A(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .X(net299));
 sky130_fd_sc_hd__buf_6 _2952_ (.A(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\Inst_RegFile_32x4.mem[20][0] ),
    .X(net452));
 sky130_fd_sc_hd__buf_1 _2954_ (.A(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .X(net302));
 sky130_fd_sc_hd__buf_6 _2955_ (.A(\Inst_RegFile_switch_matrix.JS2BEG7 ),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 _2956_ (.A(net98),
    .X(net304));
 sky130_fd_sc_hd__buf_1 _2957_ (.A(net99),
    .X(net305));
 sky130_fd_sc_hd__buf_1 _2958_ (.A(net100),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 _2959_ (.A(net101),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 _2960_ (.A(net102),
    .X(net308));
 sky130_fd_sc_hd__buf_1 _2961_ (.A(net103),
    .X(net309));
 sky130_fd_sc_hd__buf_1 _2962_ (.A(net104),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_2 _2963_ (.A(net105),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_2 _2964_ (.A(S4END[4]),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 _2965_ (.A(S4END[5]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_2 _2966_ (.A(S4END[6]),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 _2967_ (.A(S4END[7]),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 _2968_ (.A(S4END[8]),
    .X(net322));
 sky130_fd_sc_hd__buf_2 _2969_ (.A(S4END[9]),
    .X(net323));
 sky130_fd_sc_hd__buf_2 _2970_ (.A(S4END[10]),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 _2971_ (.A(S4END[11]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 _2972_ (.A(S4END[12]),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 _2973_ (.A(S4END[13]),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 _2974_ (.A(S4END[14]),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 _2975_ (.A(S4END[15]),
    .X(net314));
 sky130_fd_sc_hd__buf_4 _2976_ (.A(\Inst_RegFile_switch_matrix.S4BEG0 ),
    .X(net315));
 sky130_fd_sc_hd__buf_4 _2977_ (.A(\Inst_RegFile_switch_matrix.S4BEG1 ),
    .X(net316));
 sky130_fd_sc_hd__buf_6 _2978_ (.A(\Inst_RegFile_switch_matrix.S4BEG2 ),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 _2979_ (.A(\Inst_RegFile_switch_matrix.S4BEG3 ),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 _2980_ (.A(SS4END[4]),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_2 _2981_ (.A(SS4END[5]),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_2 _2982_ (.A(SS4END[6]),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_2 _2983_ (.A(SS4END[7]),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 _2984_ (.A(SS4END[8]),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 _2985_ (.A(SS4END[9]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_2 _2986_ (.A(SS4END[10]),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 _2987_ (.A(SS4END[11]),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_2 _2988_ (.A(SS4END[12]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 _2989_ (.A(SS4END[13]),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 _2990_ (.A(SS4END[14]),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 _2991_ (.A(SS4END[15]),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\Inst_RegFile_32x4.mem[4][2] ),
    .X(net453));
 sky130_fd_sc_hd__buf_8 _2993_ (.A(\Inst_RegFile_switch_matrix.SS4BEG1 ),
    .X(net332));
 sky130_fd_sc_hd__buf_4 _2994_ (.A(\Inst_RegFile_switch_matrix.SS4BEG2 ),
    .X(net333));
 sky130_fd_sc_hd__buf_6 _2995_ (.A(\Inst_RegFile_switch_matrix.SS4BEG3 ),
    .X(net334));
 sky130_fd_sc_hd__buf_2 _2996_ (.A(clknet_1_0__leaf_UserCLK),
    .X(net344));
 sky130_fd_sc_hd__buf_6 _2997_ (.A(\Inst_RegFile_switch_matrix.W1BEG0 ),
    .X(net345));
 sky130_fd_sc_hd__buf_6 rebuffer39 (.A(net669),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_2 rebuffer5 (.A(_0394_),
    .X(net397));
 sky130_fd_sc_hd__buf_6 _3000_ (.A(\Inst_RegFile_switch_matrix.W1BEG3 ),
    .X(net348));
 sky130_fd_sc_hd__buf_6 _3001_ (.A(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .X(net349));
 sky130_fd_sc_hd__buf_6 _3002_ (.A(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .X(net350));
 sky130_fd_sc_hd__buf_6 _3003_ (.A(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .X(net351));
 sky130_fd_sc_hd__buf_1 _3004_ (.A(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .X(net352));
 sky130_fd_sc_hd__buf_6 _3005_ (.A(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .X(net353));
 sky130_fd_sc_hd__buf_6 rebuffer44 (.A(_1071_),
    .X(net436));
 sky130_fd_sc_hd__buf_1 _3007_ (.A(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .X(net355));
 sky130_fd_sc_hd__buf_6 _3008_ (.A(\Inst_RegFile_switch_matrix.JW2BEG7 ),
    .X(net356));
 sky130_fd_sc_hd__buf_1 _3009_ (.A(net126),
    .X(net357));
 sky130_fd_sc_hd__buf_1 _3010_ (.A(net127),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_2 _3011_ (.A(net128),
    .X(net359));
 sky130_fd_sc_hd__buf_1 _3012_ (.A(net129),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 _3013_ (.A(net130),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 _3014_ (.A(net131),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_2 _3015_ (.A(net132),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 _3016_ (.A(net133),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 _3017_ (.A(W6END[2]),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 _3018_ (.A(W6END[3]),
    .X(net368));
 sky130_fd_sc_hd__buf_2 _3019_ (.A(W6END[4]),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_2 _3020_ (.A(W6END[5]),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 _3021_ (.A(W6END[6]),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 _3022_ (.A(W6END[7]),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 _3023_ (.A(W6END[8]),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 _3024_ (.A(W6END[9]),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 _3025_ (.A(W6END[10]),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_2 _3026_ (.A(W6END[11]),
    .X(net376));
 sky130_fd_sc_hd__buf_8 rebuffer47 (.A(_0958_),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_1 clone53 (.A(net677),
    .X(net445));
 sky130_fd_sc_hd__buf_2 _3029_ (.A(WW4END[4]),
    .X(net377));
 sky130_fd_sc_hd__buf_2 _3030_ (.A(WW4END[5]),
    .X(net384));
 sky130_fd_sc_hd__buf_4 _3031_ (.A(WW4END[6]),
    .X(net385));
 sky130_fd_sc_hd__buf_4 _3032_ (.A(WW4END[7]),
    .X(net386));
 sky130_fd_sc_hd__buf_4 _3033_ (.A(WW4END[8]),
    .X(net387));
 sky130_fd_sc_hd__buf_4 _3034_ (.A(WW4END[9]),
    .X(net388));
 sky130_fd_sc_hd__buf_4 _3035_ (.A(WW4END[10]),
    .X(net389));
 sky130_fd_sc_hd__buf_4 _3036_ (.A(WW4END[11]),
    .X(net390));
 sky130_fd_sc_hd__buf_2 _3037_ (.A(WW4END[12]),
    .X(net391));
 sky130_fd_sc_hd__buf_2 _3038_ (.A(WW4END[13]),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_2 _3039_ (.A(WW4END[14]),
    .X(net378));
 sky130_fd_sc_hd__buf_2 _3040_ (.A(WW4END[15]),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\Inst_RegFile_32x4.mem[14][2] ),
    .X(net455));
 sky130_fd_sc_hd__buf_6 clone2 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_2 _3043_ (.A(\Inst_RegFile_switch_matrix.WW4BEG2 ),
    .X(net382));
 sky130_fd_sc_hd__buf_6 clone6 (.A(BD2),
    .X(net398));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_885 ();
 sky130_fd_sc_hd__clkbuf_2 fanout600 (.A(_0918_),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_2 fanout601 (.A(_0918_),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_2 fanout602 (.A(net603),
    .X(net602));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout603 (.A(_0918_),
    .X(net603));
 sky130_fd_sc_hd__buf_2 fanout604 (.A(_0900_),
    .X(net604));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout605 (.A(_0900_),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_2 fanout606 (.A(net607),
    .X(net606));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout607 (.A(_0900_),
    .X(net607));
 sky130_fd_sc_hd__buf_4 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__buf_6 fanout609 (.A(net611),
    .X(net609));
 sky130_fd_sc_hd__buf_2 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__buf_6 fanout611 (.A(_0896_),
    .X(net611));
 sky130_fd_sc_hd__buf_8 fanout612 (.A(A_ADR0),
    .X(net612));
 sky130_fd_sc_hd__buf_6 clone1 (.A(_0169_),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_4 fanout614 (.A(net616),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_4 fanout615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__buf_2 fanout616 (.A(A_ADR0),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_4 fanout617 (.A(A_ADR0),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_2 fanout618 (.A(net619),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_4 fanout619 (.A(A_ADR0),
    .X(net619));
 sky130_fd_sc_hd__buf_8 fanout620 (.A(net625),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_2 fanout621 (.A(net625),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_4 fanout622 (.A(net624),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_2 fanout623 (.A(net624),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_4 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__buf_6 fanout625 (.A(B_ADR0),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_4 fanout626 (.A(B_ADR0),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_2 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_4 fanout628 (.A(B_ADR0),
    .X(net628));
 sky130_fd_sc_hd__buf_2 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_4 fanout630 (.A(net632),
    .X(net630));
 sky130_fd_sc_hd__buf_2 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_2 fanout632 (.A(_0902_),
    .X(net632));
 sky130_fd_sc_hd__buf_8 fanout633 (.A(net635),
    .X(net633));
 sky130_fd_sc_hd__buf_8 fanout634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__buf_8 fanout635 (.A(BD2),
    .X(net635));
 sky130_fd_sc_hd__buf_8 fanout636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__buf_8 fanout637 (.A(BD2),
    .X(net637));
 sky130_fd_sc_hd__buf_6 fanout638 (.A(net640),
    .X(net638));
 sky130_fd_sc_hd__buf_4 fanout639 (.A(net640),
    .X(net639));
 sky130_fd_sc_hd__buf_6 fanout640 (.A(BD3),
    .X(net640));
 sky130_fd_sc_hd__buf_8 fanout641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__buf_8 fanout642 (.A(BD3),
    .X(net642));
 sky130_fd_sc_hd__buf_8 fanout643 (.A(net644),
    .X(net643));
 sky130_fd_sc_hd__buf_8 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_6 fanout645 (.A(_0368_),
    .X(net645));
 sky130_fd_sc_hd__buf_4 fanout646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__buf_2 fanout647 (.A(AD3),
    .X(net647));
 sky130_fd_sc_hd__buf_8 fanout648 (.A(net650),
    .X(net648));
 sky130_fd_sc_hd__buf_8 fanout649 (.A(net650),
    .X(net649));
 sky130_fd_sc_hd__buf_8 fanout650 (.A(AD3),
    .X(net650));
 sky130_fd_sc_hd__buf_6 fanout651 (.A(_0169_),
    .X(net651));
 sky130_fd_sc_hd__buf_8 fanout652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__buf_8 fanout653 (.A(net656),
    .X(net653));
 sky130_fd_sc_hd__buf_8 fanout654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__buf_8 fanout655 (.A(net656),
    .X(net655));
 sky130_fd_sc_hd__buf_8 fanout656 (.A(AD2),
    .X(net656));
 sky130_fd_sc_hd__buf_8 fanout657 (.A(net661),
    .X(net657));
 sky130_fd_sc_hd__buf_6 fanout658 (.A(net660),
    .X(net658));
 sky130_fd_sc_hd__buf_4 fanout659 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__buf_4 fanout660 (.A(net661),
    .X(net660));
 sky130_fd_sc_hd__buf_8 fanout661 (.A(AD1),
    .X(net661));
 sky130_fd_sc_hd__buf_8 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__buf_8 fanout663 (.A(net664),
    .X(net663));
 sky130_fd_sc_hd__buf_8 fanout664 (.A(_0142_),
    .X(net664));
 sky130_fd_sc_hd__buf_8 fanout665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__buf_12 fanout666 (.A(net669),
    .X(net666));
 sky130_fd_sc_hd__buf_2 fanout667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__buf_2 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__buf_8 fanout669 (.A(BD1),
    .X(net669));
 sky130_fd_sc_hd__buf_8 fanout670 (.A(net671),
    .X(net670));
 sky130_fd_sc_hd__buf_8 fanout671 (.A(AD0),
    .X(net671));
 sky130_fd_sc_hd__buf_2 fanout672 (.A(net674),
    .X(net672));
 sky130_fd_sc_hd__buf_2 fanout673 (.A(net674),
    .X(net673));
 sky130_fd_sc_hd__buf_2 fanout674 (.A(AD0),
    .X(net674));
 sky130_fd_sc_hd__buf_8 fanout675 (.A(net677),
    .X(net675));
 sky130_fd_sc_hd__buf_8 fanout676 (.A(net677),
    .X(net676));
 sky130_fd_sc_hd__buf_8 fanout677 (.A(net679),
    .X(net677));
 sky130_fd_sc_hd__buf_4 fanout678 (.A(net679),
    .X(net678));
 sky130_fd_sc_hd__buf_6 fanout679 (.A(_1062_),
    .X(net679));
 sky130_fd_sc_hd__buf_2 fanout680 (.A(net682),
    .X(net680));
 sky130_fd_sc_hd__buf_6 fanout681 (.A(net682),
    .X(net681));
 sky130_fd_sc_hd__buf_8 fanout682 (.A(BD0),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_4 fanout683 (.A(net684),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_4 fanout684 (.A(BD0),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_4 fanout685 (.A(net686),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_4 fanout686 (.A(net687),
    .X(net686));
 sky130_fd_sc_hd__buf_2 fanout687 (.A(_0343_),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_4 fanout688 (.A(_0343_),
    .X(net688));
 sky130_fd_sc_hd__buf_4 fanout689 (.A(_0324_),
    .X(net689));
 sky130_fd_sc_hd__buf_2 fanout690 (.A(net135),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_4 fanout691 (.A(net134),
    .X(net691));
 sky130_fd_sc_hd__buf_2 fanout692 (.A(net117),
    .X(net692));
 sky130_fd_sc_hd__buf_4 fanout693 (.A(net116),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_2 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_2 fanout695 (.A(net696),
    .X(net695));
 sky130_fd_sc_hd__buf_2 fanout696 (.A(net697),
    .X(net696));
 sky130_fd_sc_hd__buf_2 fanout697 (.A(FrameStrobe[9]),
    .X(net697));
 sky130_fd_sc_hd__buf_2 fanout698 (.A(net700),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_2 fanout699 (.A(net700),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_2 fanout700 (.A(net701),
    .X(net700));
 sky130_fd_sc_hd__buf_2 fanout701 (.A(FrameStrobe[8]),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_2 fanout702 (.A(net706),
    .X(net702));
 sky130_fd_sc_hd__buf_2 fanout703 (.A(net704),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_2 fanout704 (.A(net705),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_2 fanout705 (.A(net706),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_2 fanout706 (.A(FrameStrobe[7]),
    .X(net706));
 sky130_fd_sc_hd__buf_2 fanout707 (.A(net708),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_2 fanout708 (.A(net709),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_2 fanout709 (.A(net710),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_2 fanout710 (.A(FrameStrobe[6]),
    .X(net710));
 sky130_fd_sc_hd__buf_2 fanout711 (.A(FrameStrobe[5]),
    .X(net711));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout712 (.A(FrameStrobe[5]),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_2 fanout713 (.A(net714),
    .X(net713));
 sky130_fd_sc_hd__buf_2 fanout714 (.A(FrameStrobe[5]),
    .X(net714));
 sky130_fd_sc_hd__buf_2 fanout715 (.A(net718),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_2 fanout716 (.A(net717),
    .X(net716));
 sky130_fd_sc_hd__buf_2 fanout717 (.A(net718),
    .X(net717));
 sky130_fd_sc_hd__buf_2 fanout718 (.A(FrameStrobe[4]),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_2 fanout719 (.A(FrameStrobe[3]),
    .X(net719));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout720 (.A(FrameStrobe[3]),
    .X(net720));
 sky130_fd_sc_hd__buf_2 fanout721 (.A(net722),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_4 fanout722 (.A(FrameStrobe[3]),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_2 fanout723 (.A(net724),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_2 fanout724 (.A(net726),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_2 fanout725 (.A(net726),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_2 fanout726 (.A(FrameStrobe[2]),
    .X(net726));
 sky130_fd_sc_hd__buf_2 fanout727 (.A(net730),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_2 fanout728 (.A(net729),
    .X(net728));
 sky130_fd_sc_hd__buf_2 fanout729 (.A(net730),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_2 fanout730 (.A(FrameStrobe[1]),
    .X(net730));
 sky130_fd_sc_hd__buf_2 fanout731 (.A(net732),
    .X(net731));
 sky130_fd_sc_hd__buf_2 fanout732 (.A(net734),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_4 fanout733 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__buf_1 fanout734 (.A(FrameStrobe[12]),
    .X(net734));
 sky130_fd_sc_hd__buf_2 fanout735 (.A(net57),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_2 fanout736 (.A(net737),
    .X(net736));
 sky130_fd_sc_hd__buf_2 fanout737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_2 fanout738 (.A(net57),
    .X(net738));
 sky130_fd_sc_hd__buf_2 fanout739 (.A(FrameStrobe[10]),
    .X(net739));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout740 (.A(FrameStrobe[10]),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_2 fanout741 (.A(net742),
    .X(net741));
 sky130_fd_sc_hd__buf_2 fanout742 (.A(FrameStrobe[10]),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_2 fanout743 (.A(net744),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_2 fanout744 (.A(net746),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_2 fanout745 (.A(net746),
    .X(net745));
 sky130_fd_sc_hd__buf_1 fanout746 (.A(FrameStrobe[0]),
    .X(net746));
 sky130_fd_sc_hd__buf_4 fanout747 (.A(net56),
    .X(net747));
 sky130_fd_sc_hd__buf_4 fanout748 (.A(net55),
    .X(net748));
 sky130_fd_sc_hd__buf_2 fanout749 (.A(net750),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_2 fanout750 (.A(FrameData[7]),
    .X(net750));
 sky130_fd_sc_hd__buf_2 fanout751 (.A(net54),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_4 fanout752 (.A(net53),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_4 fanout753 (.A(net52),
    .X(net753));
 sky130_fd_sc_hd__buf_4 fanout754 (.A(net51),
    .X(net754));
 sky130_fd_sc_hd__buf_4 fanout755 (.A(net50),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 fanout756 (.A(net49),
    .X(net756));
 sky130_fd_sc_hd__buf_4 fanout757 (.A(net48),
    .X(net757));
 sky130_fd_sc_hd__buf_4 fanout758 (.A(net47),
    .X(net758));
 sky130_fd_sc_hd__buf_4 fanout759 (.A(net46),
    .X(net759));
 sky130_fd_sc_hd__buf_4 fanout760 (.A(net45),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_4 fanout761 (.A(net762),
    .X(net761));
 sky130_fd_sc_hd__buf_2 fanout762 (.A(FrameData[26]),
    .X(net762));
 sky130_fd_sc_hd__buf_4 fanout763 (.A(net44),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_4 fanout764 (.A(net43),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_4 fanout765 (.A(net42),
    .X(net765));
 sky130_fd_sc_hd__buf_4 fanout766 (.A(net41),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_4 fanout767 (.A(net40),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_4 fanout768 (.A(net39),
    .X(net768));
 sky130_fd_sc_hd__buf_4 fanout769 (.A(net38),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_4 fanout770 (.A(net37),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_4 fanout771 (.A(net36),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_4 fanout772 (.A(net35),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_4 fanout773 (.A(net34),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_4 fanout774 (.A(net33),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_4 fanout775 (.A(net32),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_4 fanout776 (.A(net31),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_4 fanout777 (.A(net30),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_4 fanout778 (.A(net29),
    .X(net778));
 sky130_fd_sc_hd__buf_4 fanout779 (.A(net28),
    .X(net779));
 sky130_fd_sc_hd__buf_4 fanout780 (.A(net27),
    .X(net780));
 sky130_fd_sc_hd__buf_2 fanout781 (.A(net22),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_4 fanout782 (.A(net21),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_4 fanout783 (.A(net4),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_4 fanout784 (.A(net3),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(E1END[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input2 (.A(E1END[1]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(E1END[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(E1END[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(E2END[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(E2END[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(E2END[2]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(E2END[3]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(E2END[4]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(E2END[5]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(E2END[6]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(E2END[7]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(E2MID[0]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(E2MID[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(E2MID[2]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(E2MID[3]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(E2MID[4]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(E2MID[5]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(E2MID[6]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(E2MID[7]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(E6END[0]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(E6END[1]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(EE4END[0]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(EE4END[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(EE4END[2]),
    .X(net25));
 sky130_fd_sc_hd__buf_6 input26 (.A(EE4END[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(FrameData[0]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(FrameData[10]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(FrameData[11]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(FrameData[12]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(FrameData[13]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(FrameData[14]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(FrameData[15]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(FrameData[16]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(FrameData[17]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(FrameData[18]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(FrameData[19]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(FrameData[1]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(FrameData[20]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(FrameData[21]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(FrameData[22]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(FrameData[23]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(FrameData[24]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(FrameData[25]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(FrameData[27]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(FrameData[28]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(FrameData[29]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(FrameData[2]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(FrameData[30]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(FrameData[31]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(FrameData[3]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(FrameData[4]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(FrameData[5]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(FrameData[6]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(FrameData[8]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(FrameData[9]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(FrameStrobe[11]),
    .X(net57));
 sky130_fd_sc_hd__buf_4 input58 (.A(N1END[0]),
    .X(net58));
 sky130_fd_sc_hd__buf_12 input59 (.A(N1END[1]),
    .X(net59));
 sky130_fd_sc_hd__buf_4 input60 (.A(N1END[2]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(N1END[3]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(N2END[0]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(N2END[1]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(N2END[2]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(N2END[3]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(N2END[4]),
    .X(net66));
 sky130_fd_sc_hd__buf_6 input67 (.A(N2END[5]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(N2END[6]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input69 (.A(N2END[7]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(N2MID[0]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(N2MID[1]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input72 (.A(N2MID[2]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(N2MID[3]),
    .X(net73));
 sky130_fd_sc_hd__buf_2 input74 (.A(N2MID[4]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(N2MID[5]),
    .X(net75));
 sky130_fd_sc_hd__buf_2 input76 (.A(N2MID[6]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(N2MID[7]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(N4END[0]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(N4END[1]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input80 (.A(N4END[2]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(N4END[3]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 input82 (.A(NN4END[0]),
    .X(net82));
 sky130_fd_sc_hd__buf_2 input83 (.A(NN4END[1]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(NN4END[2]),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input85 (.A(NN4END[3]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 input86 (.A(S1END[0]),
    .X(net86));
 sky130_fd_sc_hd__buf_4 input87 (.A(S1END[1]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(S1END[2]),
    .X(net88));
 sky130_fd_sc_hd__buf_6 input89 (.A(S1END[3]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(S2END[0]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(S2END[1]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(S2END[2]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(S2END[3]),
    .X(net93));
 sky130_fd_sc_hd__buf_2 input94 (.A(S2END[4]),
    .X(net94));
 sky130_fd_sc_hd__buf_6 input95 (.A(S2END[5]),
    .X(net95));
 sky130_fd_sc_hd__dlymetal6s2s_1 input96 (.A(S2END[6]),
    .X(net96));
 sky130_fd_sc_hd__buf_2 input97 (.A(S2END[7]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(S2MID[0]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input99 (.A(S2MID[1]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(S2MID[2]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(S2MID[3]),
    .X(net101));
 sky130_fd_sc_hd__dlymetal6s2s_1 input102 (.A(S2MID[4]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(S2MID[5]),
    .X(net103));
 sky130_fd_sc_hd__dlymetal6s2s_1 input104 (.A(S2MID[6]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(S2MID[7]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 input106 (.A(S4END[0]),
    .X(net106));
 sky130_fd_sc_hd__buf_2 input107 (.A(S4END[1]),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(S4END[2]),
    .X(net108));
 sky130_fd_sc_hd__buf_2 input109 (.A(S4END[3]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 input110 (.A(SS4END[0]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 input111 (.A(SS4END[1]),
    .X(net111));
 sky130_fd_sc_hd__buf_2 input112 (.A(SS4END[2]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(SS4END[3]),
    .X(net113));
 sky130_fd_sc_hd__buf_4 input114 (.A(W1END[0]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(W1END[1]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(W1END[2]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(W1END[3]),
    .X(net117));
 sky130_fd_sc_hd__dlymetal6s2s_1 input118 (.A(W2END[0]),
    .X(net118));
 sky130_fd_sc_hd__buf_2 input119 (.A(W2END[1]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 input120 (.A(W2END[2]),
    .X(net120));
 sky130_fd_sc_hd__buf_2 input121 (.A(W2END[3]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 input122 (.A(W2END[4]),
    .X(net122));
 sky130_fd_sc_hd__buf_2 input123 (.A(W2END[5]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(W2END[6]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(W2END[7]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(W2MID[0]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(W2MID[1]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(W2MID[2]),
    .X(net128));
 sky130_fd_sc_hd__buf_2 input129 (.A(W2MID[3]),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input130 (.A(W2MID[4]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(W2MID[5]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(W2MID[6]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(W2MID[7]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input134 (.A(W6END[0]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(W6END[1]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 input136 (.A(WW4END[0]),
    .X(net136));
 sky130_fd_sc_hd__buf_2 input137 (.A(WW4END[1]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input138 (.A(WW4END[2]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 input139 (.A(WW4END[3]),
    .X(net139));
 sky130_fd_sc_hd__buf_6 output140 (.A(\Inst_RegFile_switch_matrix.E1BEG0 ),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__buf_8 output141 (.A(net141),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__buf_8 output142 (.A(\Inst_RegFile_switch_matrix.E1BEG2 ),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__buf_8 output143 (.A(\Inst_RegFile_switch_matrix.E1BEG3 ),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__buf_8 output144 (.A(net144),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__buf_8 output145 (.A(net145),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__buf_8 output146 (.A(net146),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__buf_6 output147 (.A(net147),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__buf_8 output148 (.A(\Inst_RegFile_switch_matrix.E2BEG4 ),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net149),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__buf_8 output150 (.A(\Inst_RegFile_switch_matrix.E2BEG6 ),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__buf_4 output151 (.A(net151),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__buf_6 output161 (.A(net161),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__buf_6 output162 (.A(\Inst_RegFile_switch_matrix.E6BEG1 ),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__buf_6 output175 (.A(net175),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__buf_6 output176 (.A(\Inst_RegFile_switch_matrix.EE4BEG1 ),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__buf_8 output177 (.A(net177),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__buf_6 output178 (.A(net178),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net226),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net232),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_6 output240 (.A(net240),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__buf_8 output241 (.A(net241),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__buf_8 output242 (.A(net242),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_6 output243 (.A(\Inst_RegFile_switch_matrix.N1BEG3 ),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_8 output244 (.A(net244),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_8 output245 (.A(net245),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_8 output246 (.A(net246),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_8 output248 (.A(net248),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_4 output249 (.A(net249),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_8 output250 (.A(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_8 output251 (.A(net251),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_6 output263 (.A(net263),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_6 output265 (.A(\Inst_RegFile_switch_matrix.N4BEG2 ),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_6 output266 (.A(net266),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_6 output279 (.A(\Inst_RegFile_switch_matrix.NN4BEG0 ),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__buf_8 output280 (.A(\Inst_RegFile_switch_matrix.NN4BEG1 ),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_8 output281 (.A(net281),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_6 output282 (.A(net282),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_6 output292 (.A(net292),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_6 output293 (.A(\Inst_RegFile_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__buf_6 output294 (.A(\Inst_RegFile_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_8 output295 (.A(\Inst_RegFile_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_8 output296 (.A(net296),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_6 output297 (.A(net297),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_8 output298 (.A(net298),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_8 output299 (.A(net299),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_8 output300 (.A(net300),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__buf_8 output301 (.A(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__buf_8 output303 (.A(net303),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__buf_4 output315 (.A(net315),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__buf_6 output316 (.A(net316),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__buf_8 output317 (.A(net317),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_4 output318 (.A(net318),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__buf_6 output331 (.A(\Inst_RegFile_switch_matrix.SS4BEG0 ),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__buf_8 output332 (.A(net332),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__buf_4 output333 (.A(net333),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__buf_6 output334 (.A(net334),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__buf_2 output335 (.A(net335),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__buf_2 output336 (.A(net336),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__buf_1 output344 (.A(net344),
    .X(UserCLKo));
 sky130_fd_sc_hd__buf_6 output345 (.A(net345),
    .X(W1BEG[0]));
 sky130_fd_sc_hd__buf_6 output346 (.A(\Inst_RegFile_switch_matrix.W1BEG1 ),
    .X(W1BEG[1]));
 sky130_fd_sc_hd__buf_6 output347 (.A(\Inst_RegFile_switch_matrix.W1BEG2 ),
    .X(W1BEG[2]));
 sky130_fd_sc_hd__buf_6 output348 (.A(net348),
    .X(W1BEG[3]));
 sky130_fd_sc_hd__buf_8 output349 (.A(net349),
    .X(W2BEG[0]));
 sky130_fd_sc_hd__buf_8 output350 (.A(net350),
    .X(W2BEG[1]));
 sky130_fd_sc_hd__buf_8 output351 (.A(net351),
    .X(W2BEG[2]));
 sky130_fd_sc_hd__buf_2 output352 (.A(net352),
    .X(W2BEG[3]));
 sky130_fd_sc_hd__buf_8 output353 (.A(net353),
    .X(W2BEG[4]));
 sky130_fd_sc_hd__buf_6 output354 (.A(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .X(W2BEG[5]));
 sky130_fd_sc_hd__buf_4 output355 (.A(net355),
    .X(W2BEG[6]));
 sky130_fd_sc_hd__buf_6 output356 (.A(net356),
    .X(W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .X(W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .X(W6BEG[0]));
 sky130_fd_sc_hd__buf_8 output366 (.A(\Inst_RegFile_switch_matrix.W6BEG0 ),
    .X(W6BEG[10]));
 sky130_fd_sc_hd__buf_8 output367 (.A(\Inst_RegFile_switch_matrix.W6BEG1 ),
    .X(W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .X(W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .X(W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .X(W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .X(W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net375),
    .X(W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .X(W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output377 (.A(net377),
    .X(WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net378),
    .X(WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(WW4BEG[11]));
 sky130_fd_sc_hd__buf_6 output380 (.A(\Inst_RegFile_switch_matrix.WW4BEG0 ),
    .X(WW4BEG[12]));
 sky130_fd_sc_hd__buf_8 output381 (.A(\Inst_RegFile_switch_matrix.WW4BEG1 ),
    .X(WW4BEG[13]));
 sky130_fd_sc_hd__buf_6 output382 (.A(net382),
    .X(WW4BEG[14]));
 sky130_fd_sc_hd__buf_8 output383 (.A(\Inst_RegFile_switch_matrix.WW4BEG3 ),
    .X(WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output384 (.A(net384),
    .X(WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .X(WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .X(WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output387 (.A(net387),
    .X(WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output388 (.A(net388),
    .X(WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output389 (.A(net389),
    .X(WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net390),
    .X(WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output391 (.A(net391),
    .X(WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .X(WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_UserCLK (.A(UserCLK),
    .X(UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK_regs (.A(UserCLK_regs),
    .X(clknet_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_0_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_1_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_2_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_3_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_4_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_5_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_6_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_7_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_8_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_9_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_10_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_11_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_12_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_13_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_14_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_4_15_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_4_0_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_4_1_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_4_2_0_UserCLK_regs));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_4_3_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_4_4_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload5 (.A(clknet_4_5_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload6 (.A(clknet_4_6_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_4 clkload7 (.A(clknet_4_8_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_4 clkload8 (.A(clknet_4_9_0_UserCLK_regs));
 sky130_fd_sc_hd__bufinv_16 clkload9 (.A(clknet_4_10_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_4_11_0_UserCLK_regs));
 sky130_fd_sc_hd__bufinv_16 clkload11 (.A(clknet_4_12_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_4 clkload12 (.A(clknet_4_14_0_UserCLK_regs));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_4_15_0_UserCLK_regs));
 sky130_fd_sc_hd__buf_6 rebuffer4 (.A(_0139_),
    .X(net396));
 sky130_fd_sc_hd__buf_8 clone12 (.A(net412),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 clone13 (.A(AD3),
    .X(net405));
 sky130_fd_sc_hd__buf_8 clone14 (.A(net669),
    .X(net406));
 sky130_fd_sc_hd__buf_8 clone15 (.A(net653),
    .X(net407));
 sky130_fd_sc_hd__buf_6 rebuffer20 (.A(BD3),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 clone21 (.A(net656),
    .X(net413));
 sky130_fd_sc_hd__buf_8 clone22 (.A(net671),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 clone23 (.A(net661),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_1 clone24 (.A(net663),
    .X(net416));
 sky130_fd_sc_hd__buf_6 clone25 (.A(net644),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_1 clone26 (.A(N1END[1]),
    .X(net418));
 sky130_fd_sc_hd__dlymetal6s2s_1 clone27 (.A(net655),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\Inst_RegFile_32x4.mem[18][3] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\Inst_RegFile_32x4.mem[22][1] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\Inst_RegFile_32x4.mem[18][0] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\Inst_RegFile_32x4.mem[6][2] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\Inst_RegFile_32x4.mem[3][3] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\Inst_RegFile_32x4.mem[2][3] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\Inst_RegFile_32x4.mem[18][1] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\Inst_RegFile_32x4.mem[30][2] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\Inst_RegFile_32x4.mem[10][2] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\Inst_RegFile_32x4.mem[18][2] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\Inst_RegFile_32x4.mem[8][2] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\Inst_RegFile_32x4.mem[10][3] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\Inst_RegFile_32x4.mem[26][0] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\Inst_RegFile_32x4.mem[10][0] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\Inst_RegFile_32x4.mem[24][0] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\Inst_RegFile_32x4.mem[26][2] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\Inst_RegFile_32x4.mem[20][1] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\Inst_RegFile_32x4.mem[16][2] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\Inst_RegFile_32x4.mem[28][2] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\Inst_RegFile_32x4.mem[0][0] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\Inst_RegFile_32x4.mem[8][0] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\Inst_RegFile_32x4.mem[14][0] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\Inst_RegFile_32x4.mem[12][0] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\Inst_RegFile_32x4.mem[16][0] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\Inst_RegFile_32x4.mem[8][3] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\Inst_RegFile_32x4.mem[2][1] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\Inst_RegFile_32x4.mem[28][1] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\Inst_RegFile_32x4.mem[26][1] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\Inst_RegFile_32x4.mem[24][2] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\Inst_RegFile_32x4.mem[0][3] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\Inst_RegFile_32x4.mem[16][1] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\Inst_RegFile_32x4.mem[28][0] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\Inst_RegFile_32x4.mem[26][3] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\Inst_RegFile_32x4.mem[4][0] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\Inst_RegFile_32x4.mem[7][2] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\Inst_RegFile_32x4.mem[7][0] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\Inst_RegFile_32x4.mem[30][3] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\Inst_RegFile_32x4.mem[9][2] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\Inst_RegFile_32x4.mem[20][3] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\Inst_RegFile_32x4.mem[12][3] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\Inst_RegFile_32x4.mem[5][2] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\Inst_RegFile_32x4.mem[0][2] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\Inst_RegFile_32x4.mem[20][2] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\Inst_RegFile_32x4.mem[6][3] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\Inst_RegFile_32x4.mem[31][2] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\Inst_RegFile_32x4.mem[2][0] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\Inst_RegFile_32x4.mem[3][0] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\Inst_RegFile_32x4.mem[5][0] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\Inst_RegFile_32x4.mem[5][3] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\Inst_RegFile_32x4.mem[30][1] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\Inst_RegFile_32x4.mem[24][1] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\Inst_RegFile_32x4.mem[11][2] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\Inst_RegFile_32x4.mem[7][1] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\Inst_RegFile_32x4.mem[11][0] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\Inst_RegFile_32x4.mem[23][1] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\Inst_RegFile_32x4.mem[8][1] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\Inst_RegFile_32x4.mem[2][2] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\Inst_RegFile_32x4.mem[14][3] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\Inst_RegFile_32x4.mem[3][1] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\Inst_RegFile_32x4.mem[15][0] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\Inst_RegFile_32x4.mem[1][2] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\Inst_RegFile_32x4.mem[1][1] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\Inst_RegFile_32x4.mem[22][0] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\Inst_RegFile_32x4.mem[0][1] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\Inst_RegFile_32x4.mem[4][1] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\Inst_RegFile_32x4.mem[28][3] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\Inst_RegFile_32x4.mem[31][0] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\Inst_RegFile_32x4.mem[1][0] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\Inst_RegFile_32x4.mem[6][0] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\Inst_RegFile_32x4.mem[9][3] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\Inst_RegFile_32x4.mem[3][2] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\Inst_RegFile_32x4.mem[17][1] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\Inst_RegFile_32x4.mem[15][3] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\Inst_RegFile_32x4.mem[1][3] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\Inst_RegFile_32x4.mem[31][3] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\Inst_RegFile_32x4.mem[25][0] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\Inst_RegFile_32x4.mem[5][1] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\Inst_RegFile_32x4.mem[14][1] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\Inst_RegFile_32x4.mem[7][3] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\Inst_RegFile_32x4.mem[24][3] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\Inst_RegFile_32x4.mem[21][0] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\Inst_RegFile_32x4.mem[6][1] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\Inst_RegFile_32x4.mem[27][1] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\Inst_RegFile_32x4.mem[29][2] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\Inst_RegFile_32x4.mem[22][3] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\Inst_RegFile_32x4.mem[22][2] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\Inst_RegFile_32x4.mem[12][1] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\Inst_RegFile_32x4.mem[31][1] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\Inst_RegFile_32x4.mem[19][2] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\Inst_RegFile_32x4.mem[13][2] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\Inst_RegFile_32x4.mem[11][1] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\Inst_RegFile_32x4.mem[19][0] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\Inst_RegFile_32x4.mem[9][1] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\Inst_RegFile_32x4.mem[27][2] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\Inst_RegFile_32x4.mem[25][1] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\Inst_RegFile_32x4.mem[10][1] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\Inst_RegFile_32x4.mem[29][1] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\Inst_RegFile_32x4.mem[16][3] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\Inst_RegFile_32x4.mem[19][1] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\Inst_RegFile_32x4.mem[27][0] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\Inst_RegFile_32x4.mem[29][0] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\Inst_RegFile_32x4.mem[15][1] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\Inst_RegFile_32x4.mem[30][0] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\Inst_RegFile_32x4.mem[17][0] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\Inst_RegFile_32x4.mem[21][2] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\Inst_RegFile_32x4.mem[9][0] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\Inst_RegFile_32x4.mem[29][3] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\Inst_RegFile_32x4.mem[25][2] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\Inst_RegFile_32x4.mem[17][2] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\Inst_RegFile_32x4.mem[21][3] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\Inst_RegFile_32x4.mem[13][3] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\Inst_RegFile_32x4.mem[13][0] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\Inst_RegFile_32x4.mem[19][3] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\Inst_RegFile_32x4.mem[11][3] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\Inst_RegFile_32x4.mem[25][3] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\Inst_RegFile_32x4.mem[27][3] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\Inst_RegFile_32x4.mem[23][0] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\Inst_RegFile_32x4.mem[23][3] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\Inst_RegFile_32x4.mem[17][3] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\Inst_RegFile_32x4.mem[13][1] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\Inst_RegFile_32x4.mem[23][2] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\Inst_RegFile_32x4.mem[21][1] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\Inst_RegFile_32x4.mem[15][2] ),
    .X(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(E6END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(E6END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(E6END[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(E6END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(E6END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(E6END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(E6END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(E6END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(EE4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(EE4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(EE4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(EE4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(EE4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(EE4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(EE4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(EE4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(EE4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(EE4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(EE4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(FrameData[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(FrameStrobe[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(FrameStrobe[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(FrameStrobe[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(FrameStrobe[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(FrameStrobe[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(FrameStrobe[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(FrameStrobe[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(FrameStrobe[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(FrameStrobe[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(FrameStrobe[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(FrameStrobe[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(N4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(N4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(N4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(N4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(N4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(N4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(N4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(N4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(N4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(N4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(N4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(N4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(NN4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(NN4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(NN4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(NN4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(NN4END[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(NN4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(NN4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(NN4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(NN4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(NN4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(NN4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(NN4END[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(W2END[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net760));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(EE4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(EE4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(\Inst_RegFile_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(\Inst_RegFile_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(W2MID[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net747));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net111));
 sky130_fd_sc_hd__decap_3 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_471 ();
endmodule
