module W_term_single (UserCLK,
    UserCLKo,
    E1BEG,
    E2BEG,
    E2BEGb,
    E6BEG,
    EE4BEG,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    W1END,
    W2END,
    W2MID,
    W6END,
    WW4END);
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 output [11:0] E6BEG;
 output [15:0] EE4BEG;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] W1END;
 input [7:0] W2END;
 input [7:0] W2MID;
 input [11:0] W6END;
 input [15:0] WW4END;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;

 sky130_fd_sc_hd__buf_1 _000_ (.A(W1END[3]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 _001_ (.A(W1END[2]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 _002_ (.A(W1END[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 _003_ (.A(W1END[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 _004_ (.A(W2MID[7]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 _005_ (.A(W2MID[6]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 _006_ (.A(W2MID[5]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 _007_ (.A(W2MID[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 _008_ (.A(W2MID[3]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 _009_ (.A(W2MID[2]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 _010_ (.A(W2MID[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 _011_ (.A(W2MID[0]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 _012_ (.A(W2END[7]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 _013_ (.A(W2END[6]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 _014_ (.A(W2END[5]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 _015_ (.A(W2END[4]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 _016_ (.A(W2END[3]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 _017_ (.A(W2END[2]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 _018_ (.A(W2END[1]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 _019_ (.A(W2END[0]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 _020_ (.A(W6END[11]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 _021_ (.A(W6END[10]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 _022_ (.A(W6END[9]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 _023_ (.A(W6END[8]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 _024_ (.A(W6END[7]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 _025_ (.A(W6END[6]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 _026_ (.A(W6END[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 _027_ (.A(W6END[4]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 _028_ (.A(W6END[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 _029_ (.A(W6END[2]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 _030_ (.A(W6END[1]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 _031_ (.A(W6END[0]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 _032_ (.A(WW4END[15]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 _033_ (.A(WW4END[14]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 _034_ (.A(WW4END[13]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 _035_ (.A(WW4END[12]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _036_ (.A(WW4END[11]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 _037_ (.A(WW4END[10]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 _038_ (.A(WW4END[9]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 _039_ (.A(WW4END[8]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 _040_ (.A(WW4END[7]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 _041_ (.A(WW4END[6]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 _042_ (.A(WW4END[5]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 _043_ (.A(WW4END[4]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 _044_ (.A(WW4END[3]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 _045_ (.A(WW4END[2]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 _046_ (.A(WW4END[1]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 _047_ (.A(WW4END[0]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 _048_ (.A(FrameData[0]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _049_ (.A(FrameData[1]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 _050_ (.A(FrameData[2]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _051_ (.A(FrameData[3]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _052_ (.A(FrameData[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _053_ (.A(FrameData[5]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _054_ (.A(FrameData[6]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _055_ (.A(FrameData[7]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 _056_ (.A(FrameData[8]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _057_ (.A(FrameData[9]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 _058_ (.A(FrameData[10]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 _059_ (.A(FrameData[11]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 _060_ (.A(FrameData[12]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 _061_ (.A(FrameData[13]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 _062_ (.A(FrameData[14]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _063_ (.A(FrameData[15]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _064_ (.A(FrameData[16]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _065_ (.A(FrameData[17]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 _066_ (.A(FrameData[18]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _067_ (.A(FrameData[19]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 _068_ (.A(FrameData[20]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _069_ (.A(FrameData[21]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _070_ (.A(FrameData[22]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _071_ (.A(FrameData[23]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _072_ (.A(FrameData[24]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _073_ (.A(FrameData[25]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _074_ (.A(FrameData[26]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(FrameData[27]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _076_ (.A(FrameData[28]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _077_ (.A(FrameData[29]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _078_ (.A(FrameData[30]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(FrameData[31]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 _080_ (.A(FrameStrobe[0]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 _081_ (.A(FrameStrobe[1]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 _082_ (.A(FrameStrobe[2]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 _083_ (.A(FrameStrobe[3]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 _084_ (.A(FrameStrobe[4]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 _085_ (.A(FrameStrobe[5]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 _086_ (.A(FrameStrobe[6]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 _087_ (.A(FrameStrobe[7]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 _088_ (.A(FrameStrobe[8]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(FrameStrobe[9]),
    .X(net100));
 sky130_fd_sc_hd__buf_1 _090_ (.A(FrameStrobe[10]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 _091_ (.A(FrameStrobe[11]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 _092_ (.A(FrameStrobe[12]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _093_ (.A(FrameStrobe[13]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 _094_ (.A(FrameStrobe[14]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 _095_ (.A(FrameStrobe[15]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 _096_ (.A(FrameStrobe[16]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 _097_ (.A(FrameStrobe[17]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 _098_ (.A(FrameStrobe[18]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 _099_ (.A(FrameStrobe[19]),
    .X(net91));
 sky130_fd_sc_hd__buf_2 _100_ (.A(UserCLK),
    .X(net101));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_223 ();
 sky130_fd_sc_hd__buf_2 output1 (.A(net1),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(UserCLKo));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(FrameData[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameStrobe[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(FrameStrobe[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(FrameStrobe[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(FrameStrobe[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameStrobe[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(W2END[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(WW4END[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(FrameStrobe[17]));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_71 ();
endmodule
