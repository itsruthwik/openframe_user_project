magic
tech sky130A
magscale 1 2
timestamp 1746697978
<< viali >>
rect 1869 8585 1903 8619
rect 4077 8585 4111 8619
rect 6469 8585 6503 8619
rect 8309 8585 8343 8619
rect 10425 8585 10459 8619
rect 12541 8585 12575 8619
rect 14657 8585 14691 8619
rect 16773 8585 16807 8619
rect 18889 8585 18923 8619
rect 21005 8585 21039 8619
rect 23121 8585 23155 8619
rect 25237 8585 25271 8619
rect 27353 8585 27387 8619
rect 29653 8585 29687 8619
rect 31585 8585 31619 8619
rect 33701 8585 33735 8619
rect 35817 8585 35851 8619
rect 37933 8585 37967 8619
rect 40141 8585 40175 8619
rect 42625 8585 42659 8619
rect 43269 8585 43303 8619
rect 44005 8585 44039 8619
rect 44373 8585 44407 8619
rect 2053 8449 2087 8483
rect 4261 8449 4295 8483
rect 6653 8449 6687 8483
rect 8493 8449 8527 8483
rect 10609 8449 10643 8483
rect 12725 8449 12759 8483
rect 14841 8449 14875 8483
rect 16957 8449 16991 8483
rect 19073 8449 19107 8483
rect 21189 8449 21223 8483
rect 23305 8449 23339 8483
rect 25421 8449 25455 8483
rect 27537 8449 27571 8483
rect 29837 8449 29871 8483
rect 31769 8449 31803 8483
rect 33885 8449 33919 8483
rect 36001 8449 36035 8483
rect 38117 8449 38151 8483
rect 39957 8449 39991 8483
rect 42441 8449 42475 8483
rect 43085 8449 43119 8483
rect 43453 8449 43487 8483
rect 43821 8449 43855 8483
rect 44189 8449 44223 8483
rect 43637 8313 43671 8347
rect 6193 8041 6227 8075
rect 9965 8041 9999 8075
rect 11989 8041 12023 8075
rect 36553 8041 36587 8075
rect 38117 8041 38151 8075
rect 39865 8041 39899 8075
rect 40877 8041 40911 8075
rect 41613 8041 41647 8075
rect 41981 8041 42015 8075
rect 42717 8041 42751 8075
rect 43729 8041 43763 8075
rect 42257 7973 42291 8007
rect 42993 7973 43027 8007
rect 43361 7973 43395 8007
rect 2697 7905 2731 7939
rect 3065 7905 3099 7939
rect 3433 7905 3467 7939
rect 3249 7837 3283 7871
rect 9873 7837 9907 7871
rect 10149 7837 10183 7871
rect 12173 7837 12207 7871
rect 12265 7837 12299 7871
rect 14289 7837 14323 7871
rect 23581 7837 23615 7871
rect 32597 7837 32631 7871
rect 34897 7837 34931 7871
rect 36001 7837 36035 7871
rect 36737 7837 36771 7871
rect 38301 7837 38335 7871
rect 39497 7837 39531 7871
rect 40049 7837 40083 7871
rect 40693 7837 40727 7871
rect 41337 7837 41371 7871
rect 41705 7837 41739 7871
rect 41797 7837 41831 7871
rect 42073 7837 42107 7871
rect 42533 7837 42567 7871
rect 42809 7837 42843 7871
rect 43177 7837 43211 7871
rect 43545 7837 43579 7871
rect 43913 7837 43947 7871
rect 44281 7837 44315 7871
rect 2513 7769 2547 7803
rect 2881 7769 2915 7803
rect 6101 7769 6135 7803
rect 35449 7769 35483 7803
rect 35633 7769 35667 7803
rect 12449 7701 12483 7735
rect 14105 7701 14139 7735
rect 23765 7701 23799 7735
rect 32413 7701 32447 7735
rect 34713 7701 34747 7735
rect 35817 7701 35851 7735
rect 39313 7701 39347 7735
rect 41521 7701 41555 7735
rect 42349 7701 42383 7735
rect 44097 7701 44131 7735
rect 44465 7701 44499 7735
rect 26341 7497 26375 7531
rect 44097 7497 44131 7531
rect 35449 7429 35483 7463
rect 12081 7361 12115 7395
rect 14381 7361 14415 7395
rect 26157 7361 26191 7395
rect 28733 7361 28767 7395
rect 28825 7361 28859 7395
rect 35633 7361 35667 7395
rect 41429 7361 41463 7395
rect 43821 7361 43855 7395
rect 43913 7361 43947 7395
rect 44281 7361 44315 7395
rect 12265 7225 12299 7259
rect 14565 7157 14599 7191
rect 28641 7157 28675 7191
rect 29009 7157 29043 7191
rect 41245 7157 41279 7191
rect 43637 7157 43671 7191
rect 44465 7157 44499 7191
rect 2789 6817 2823 6851
rect 2605 6749 2639 6783
rect 31585 6749 31619 6783
rect 31677 6749 31711 6783
rect 41429 6749 41463 6783
rect 43913 6749 43947 6783
rect 44281 6749 44315 6783
rect 5973 6681 6007 6715
rect 6193 6681 6227 6715
rect 31493 6613 31527 6647
rect 31861 6613 31895 6647
rect 41245 6613 41279 6647
rect 44097 6613 44131 6647
rect 44465 6613 44499 6647
rect 36921 6409 36955 6443
rect 38209 6409 38243 6443
rect 40693 6409 40727 6443
rect 43085 6409 43119 6443
rect 44465 6409 44499 6443
rect 4353 6273 4387 6307
rect 5089 6273 5123 6307
rect 18153 6273 18187 6307
rect 22845 6273 22879 6307
rect 23029 6273 23063 6307
rect 25789 6273 25823 6307
rect 37105 6273 37139 6307
rect 37473 6273 37507 6307
rect 38393 6273 38427 6307
rect 39589 6273 39623 6307
rect 40877 6273 40911 6307
rect 42809 6273 42843 6307
rect 42901 6273 42935 6307
rect 43913 6273 43947 6307
rect 44281 6273 44315 6307
rect 4537 6137 4571 6171
rect 23213 6137 23247 6171
rect 37289 6137 37323 6171
rect 39405 6137 39439 6171
rect 44097 6137 44131 6171
rect 5181 6069 5215 6103
rect 18337 6069 18371 6103
rect 25973 6069 26007 6103
rect 27169 5797 27203 5831
rect 44465 5797 44499 5831
rect 2237 5729 2271 5763
rect 43177 5729 43211 5763
rect 2053 5661 2087 5695
rect 16313 5661 16347 5695
rect 16773 5661 16807 5695
rect 22385 5661 22419 5695
rect 26985 5661 27019 5695
rect 31585 5661 31619 5695
rect 31677 5661 31711 5695
rect 43269 5661 43303 5695
rect 43361 5661 43395 5695
rect 43913 5661 43947 5695
rect 44281 5661 44315 5695
rect 16497 5525 16531 5559
rect 16589 5525 16623 5559
rect 22569 5525 22603 5559
rect 31493 5525 31527 5559
rect 31861 5525 31895 5559
rect 43545 5525 43579 5559
rect 44097 5525 44131 5559
rect 43269 5321 43303 5355
rect 44465 5321 44499 5355
rect 3065 5253 3099 5287
rect 16037 5185 16071 5219
rect 20453 5185 20487 5219
rect 31493 5185 31527 5219
rect 42441 5185 42475 5219
rect 42717 5185 42751 5219
rect 42993 5185 43027 5219
rect 43085 5185 43119 5219
rect 43913 5185 43947 5219
rect 44281 5185 44315 5219
rect 3249 5117 3283 5151
rect 42901 5049 42935 5083
rect 44097 5049 44131 5083
rect 16221 4981 16255 5015
rect 20637 4981 20671 5015
rect 31677 4981 31711 5015
rect 42625 4981 42659 5015
rect 43821 4777 43855 4811
rect 42809 4709 42843 4743
rect 44465 4709 44499 4743
rect 23213 4641 23247 4675
rect 42441 4641 42475 4675
rect 2145 4573 2179 4607
rect 6285 4573 6319 4607
rect 6653 4573 6687 4607
rect 7113 4573 7147 4607
rect 10885 4573 10919 4607
rect 11897 4573 11931 4607
rect 12817 4573 12851 4607
rect 14105 4573 14139 4607
rect 16405 4573 16439 4607
rect 23305 4573 23339 4607
rect 23397 4573 23431 4607
rect 39313 4573 39347 4607
rect 41153 4573 41187 4607
rect 41429 4573 41463 4607
rect 42533 4573 42567 4607
rect 42625 4573 42659 4607
rect 43637 4573 43671 4607
rect 43913 4573 43947 4607
rect 44281 4573 44315 4607
rect 2329 4505 2363 4539
rect 6469 4437 6503 4471
rect 6837 4437 6871 4471
rect 7297 4437 7331 4471
rect 11069 4437 11103 4471
rect 12081 4437 12115 4471
rect 13001 4437 13035 4471
rect 14289 4437 14323 4471
rect 16589 4437 16623 4471
rect 23581 4437 23615 4471
rect 39129 4437 39163 4471
rect 41061 4437 41095 4471
rect 41245 4437 41279 4471
rect 44097 4437 44131 4471
rect 43361 4233 43395 4267
rect 4997 4097 5031 4131
rect 7665 4097 7699 4131
rect 9873 4097 9907 4131
rect 27077 4097 27111 4131
rect 38577 4097 38611 4131
rect 43085 4097 43119 4131
rect 43177 4097 43211 4131
rect 43913 4097 43947 4131
rect 44281 4097 44315 4131
rect 42993 3961 43027 3995
rect 44097 3961 44131 3995
rect 44465 3961 44499 3995
rect 5181 3893 5215 3927
rect 7849 3893 7883 3927
rect 10057 3893 10091 3927
rect 27261 3893 27295 3927
rect 38393 3893 38427 3927
rect 17141 3689 17175 3723
rect 34897 3689 34931 3723
rect 43085 3689 43119 3723
rect 42809 3621 42843 3655
rect 44465 3621 44499 3655
rect 16589 3485 16623 3519
rect 16957 3485 16991 3519
rect 18705 3485 18739 3519
rect 19625 3485 19659 3519
rect 27721 3485 27755 3519
rect 27813 3485 27847 3519
rect 28365 3485 28399 3519
rect 28457 3485 28491 3519
rect 28917 3485 28951 3519
rect 29009 3485 29043 3519
rect 29561 3485 29595 3519
rect 34713 3485 34747 3519
rect 35541 3485 35575 3519
rect 42809 3485 42843 3519
rect 42901 3485 42935 3519
rect 43913 3485 43947 3519
rect 44281 3485 44315 3519
rect 16773 3349 16807 3383
rect 18889 3349 18923 3383
rect 19809 3349 19843 3383
rect 27629 3349 27663 3383
rect 27997 3349 28031 3383
rect 28273 3349 28307 3383
rect 28641 3349 28675 3383
rect 28917 3349 28951 3383
rect 29193 3349 29227 3383
rect 29745 3349 29779 3383
rect 34989 3349 35023 3383
rect 35725 3349 35759 3383
rect 44097 3349 44131 3383
rect 2329 3145 2363 3179
rect 3433 3145 3467 3179
rect 5181 3145 5215 3179
rect 41521 3145 41555 3179
rect 41889 3145 41923 3179
rect 42257 3145 42291 3179
rect 42625 3145 42659 3179
rect 43453 3145 43487 3179
rect 2973 3077 3007 3111
rect 41797 3077 41831 3111
rect 2237 3009 2271 3043
rect 2605 3009 2639 3043
rect 3341 3009 3375 3043
rect 4997 3009 5031 3043
rect 5273 3009 5307 3043
rect 17417 3009 17451 3043
rect 19349 3009 19383 3043
rect 19993 3009 20027 3043
rect 28825 3009 28859 3043
rect 30297 3009 30331 3043
rect 30389 3009 30423 3043
rect 30665 3009 30699 3043
rect 31125 3009 31159 3043
rect 31493 3009 31527 3043
rect 33701 3009 33735 3043
rect 36277 3009 36311 3043
rect 41705 3009 41739 3043
rect 42073 3009 42107 3043
rect 42441 3009 42475 3043
rect 42717 3009 42751 3043
rect 43177 3009 43211 3043
rect 43269 3009 43303 3043
rect 43913 3009 43947 3043
rect 44281 3009 44315 3043
rect 41613 2941 41647 2975
rect 41981 2941 42015 2975
rect 3157 2873 3191 2907
rect 5457 2873 5491 2907
rect 30205 2873 30239 2907
rect 30849 2873 30883 2907
rect 42901 2873 42935 2907
rect 43729 2873 43763 2907
rect 2697 2805 2731 2839
rect 17601 2805 17635 2839
rect 19533 2805 19567 2839
rect 20177 2805 20211 2839
rect 28641 2805 28675 2839
rect 30573 2805 30607 2839
rect 31309 2805 31343 2839
rect 31677 2805 31711 2839
rect 33885 2805 33919 2839
rect 36461 2805 36495 2839
rect 42993 2805 43027 2839
rect 43545 2805 43579 2839
rect 44097 2805 44131 2839
rect 44465 2805 44499 2839
rect 30849 2601 30883 2635
rect 36737 2601 36771 2635
rect 38577 2601 38611 2635
rect 42533 2601 42567 2635
rect 44465 2601 44499 2635
rect 23213 2533 23247 2567
rect 25329 2533 25363 2567
rect 27537 2533 27571 2567
rect 28641 2533 28675 2567
rect 29745 2533 29779 2567
rect 31217 2533 31251 2567
rect 32689 2533 32723 2567
rect 33793 2533 33827 2567
rect 35173 2533 35207 2567
rect 36277 2533 36311 2567
rect 37841 2533 37875 2567
rect 38853 2533 38887 2567
rect 43729 2533 43763 2567
rect 19533 2397 19567 2431
rect 19889 2397 19923 2431
rect 20269 2397 20303 2431
rect 20637 2397 20671 2431
rect 21005 2397 21039 2431
rect 21373 2397 21407 2431
rect 21925 2397 21959 2431
rect 22293 2397 22327 2431
rect 22661 2397 22695 2431
rect 23029 2397 23063 2431
rect 23397 2397 23431 2431
rect 23765 2397 23799 2431
rect 24409 2397 24443 2431
rect 24777 2397 24811 2431
rect 25145 2397 25179 2431
rect 25513 2397 25547 2431
rect 25881 2397 25915 2431
rect 26249 2397 26283 2431
rect 26985 2397 27019 2431
rect 27353 2397 27387 2431
rect 27721 2397 27755 2431
rect 28089 2397 28123 2431
rect 28457 2397 28491 2431
rect 28825 2397 28859 2431
rect 29561 2397 29595 2431
rect 29929 2397 29963 2431
rect 30297 2397 30331 2431
rect 30665 2397 30699 2431
rect 31033 2397 31067 2431
rect 31401 2397 31435 2431
rect 32137 2397 32171 2431
rect 32505 2397 32539 2431
rect 32873 2397 32907 2431
rect 33241 2397 33275 2431
rect 33609 2397 33643 2431
rect 33977 2397 34011 2431
rect 34713 2397 34747 2431
rect 35357 2397 35391 2431
rect 35449 2397 35483 2431
rect 35817 2397 35851 2431
rect 36461 2397 36495 2431
rect 36553 2397 36587 2431
rect 37289 2397 37323 2431
rect 37657 2397 37691 2431
rect 38301 2397 38335 2431
rect 38393 2397 38427 2431
rect 39037 2397 39071 2431
rect 42717 2397 42751 2431
rect 42809 2397 42843 2431
rect 43177 2397 43211 2431
rect 43545 2397 43579 2431
rect 43913 2397 43947 2431
rect 44281 2397 44315 2431
rect 2605 2329 2639 2363
rect 2789 2329 2823 2363
rect 19717 2261 19751 2295
rect 20085 2261 20119 2295
rect 20453 2261 20487 2295
rect 20821 2261 20855 2295
rect 21189 2261 21223 2295
rect 21557 2261 21591 2295
rect 22109 2261 22143 2295
rect 22477 2261 22511 2295
rect 22845 2261 22879 2295
rect 23581 2261 23615 2295
rect 23949 2261 23983 2295
rect 24593 2261 24627 2295
rect 24961 2261 24995 2295
rect 25697 2261 25731 2295
rect 26065 2261 26099 2295
rect 26433 2261 26467 2295
rect 27169 2261 27203 2295
rect 27905 2261 27939 2295
rect 28273 2261 28307 2295
rect 29009 2261 29043 2295
rect 30113 2261 30147 2295
rect 30481 2261 30515 2295
rect 31585 2261 31619 2295
rect 32321 2261 32355 2295
rect 33057 2261 33091 2295
rect 33425 2261 33459 2295
rect 34161 2261 34195 2295
rect 34897 2261 34931 2295
rect 35633 2261 35667 2295
rect 36001 2261 36035 2295
rect 37473 2261 37507 2295
rect 38117 2261 38151 2295
rect 42993 2261 43027 2295
rect 43361 2261 43395 2295
rect 44097 2261 44131 2295
<< metal1 >>
rect 23290 9324 23296 9376
rect 23348 9364 23354 9376
rect 37458 9364 37464 9376
rect 23348 9336 37464 9364
rect 23348 9324 23354 9336
rect 37458 9324 37464 9336
rect 37516 9324 37522 9376
rect 1302 9256 1308 9308
rect 1360 9296 1366 9308
rect 42518 9296 42524 9308
rect 1360 9268 42524 9296
rect 1360 9256 1366 9268
rect 42518 9256 42524 9268
rect 42576 9256 42582 9308
rect 6638 9188 6644 9240
rect 6696 9228 6702 9240
rect 34422 9228 34428 9240
rect 6696 9200 34428 9228
rect 6696 9188 6702 9200
rect 34422 9188 34428 9200
rect 34480 9188 34486 9240
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 35434 9160 35440 9172
rect 6604 9132 35440 9160
rect 6604 9120 6610 9132
rect 35434 9120 35440 9132
rect 35492 9120 35498 9172
rect 12406 9064 19334 9092
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 12406 9024 12434 9064
rect 6788 8996 12434 9024
rect 6788 8984 6794 8996
rect 19306 8956 19334 9064
rect 23198 9052 23204 9104
rect 23256 9092 23262 9104
rect 37642 9092 37648 9104
rect 23256 9064 37648 9092
rect 23256 9052 23262 9064
rect 37642 9052 37648 9064
rect 37700 9052 37706 9104
rect 25406 8984 25412 9036
rect 25464 9024 25470 9036
rect 34330 9024 34336 9036
rect 25464 8996 34336 9024
rect 25464 8984 25470 8996
rect 34330 8984 34336 8996
rect 34388 8984 34394 9036
rect 25130 8956 25136 8968
rect 19306 8928 25136 8956
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 25314 8916 25320 8968
rect 25372 8956 25378 8968
rect 44634 8956 44640 8968
rect 25372 8928 44640 8956
rect 25372 8916 25378 8928
rect 44634 8916 44640 8928
rect 44692 8916 44698 8968
rect 19058 8848 19064 8900
rect 19116 8888 19122 8900
rect 25406 8888 25412 8900
rect 19116 8860 25412 8888
rect 19116 8848 19122 8860
rect 25406 8848 25412 8860
rect 25464 8848 25470 8900
rect 32858 8888 32864 8900
rect 25516 8860 32864 8888
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 25516 8820 25544 8860
rect 32858 8848 32864 8860
rect 32916 8848 32922 8900
rect 17000 8792 25544 8820
rect 17000 8780 17006 8792
rect 29822 8780 29828 8832
rect 29880 8820 29886 8832
rect 38562 8820 38568 8832
rect 29880 8792 38568 8820
rect 29880 8780 29886 8792
rect 38562 8780 38568 8792
rect 38620 8780 38626 8832
rect 1104 8730 44896 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 44896 8730
rect 1104 8656 44896 8678
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 1857 8619 1915 8625
rect 1857 8616 1869 8619
rect 1820 8588 1869 8616
rect 1820 8576 1826 8588
rect 1857 8585 1869 8588
rect 1903 8585 1915 8619
rect 1857 8579 1915 8585
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 3936 8588 4077 8616
rect 3936 8576 3942 8588
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 6052 8588 6469 8616
rect 6052 8576 6058 8588
rect 6457 8585 6469 8588
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 8297 8619 8355 8625
rect 8297 8616 8309 8619
rect 8168 8588 8309 8616
rect 8168 8576 8174 8588
rect 8297 8585 8309 8588
rect 8343 8585 8355 8619
rect 8297 8579 8355 8585
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 10284 8588 10425 8616
rect 10284 8576 10290 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 10413 8579 10471 8585
rect 12342 8576 12348 8628
rect 12400 8616 12406 8628
rect 12529 8619 12587 8625
rect 12529 8616 12541 8619
rect 12400 8588 12541 8616
rect 12400 8576 12406 8588
rect 12529 8585 12541 8588
rect 12575 8585 12587 8619
rect 12529 8579 12587 8585
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 14645 8619 14703 8625
rect 14645 8616 14657 8619
rect 14516 8588 14657 8616
rect 14516 8576 14522 8588
rect 14645 8585 14657 8588
rect 14691 8585 14703 8619
rect 14645 8579 14703 8585
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 16761 8619 16819 8625
rect 16761 8616 16773 8619
rect 16632 8588 16773 8616
rect 16632 8576 16638 8588
rect 16761 8585 16773 8588
rect 16807 8585 16819 8619
rect 16761 8579 16819 8585
rect 16942 8576 16948 8628
rect 17000 8576 17006 8628
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 18877 8619 18935 8625
rect 18877 8616 18889 8619
rect 18748 8588 18889 8616
rect 18748 8576 18754 8588
rect 18877 8585 18889 8588
rect 18923 8585 18935 8619
rect 18877 8579 18935 8585
rect 19058 8576 19064 8628
rect 19116 8576 19122 8628
rect 20806 8576 20812 8628
rect 20864 8616 20870 8628
rect 20993 8619 21051 8625
rect 20993 8616 21005 8619
rect 20864 8588 21005 8616
rect 20864 8576 20870 8588
rect 20993 8585 21005 8588
rect 21039 8585 21051 8619
rect 20993 8579 21051 8585
rect 22922 8576 22928 8628
rect 22980 8616 22986 8628
rect 23109 8619 23167 8625
rect 23109 8616 23121 8619
rect 22980 8588 23121 8616
rect 22980 8576 22986 8588
rect 23109 8585 23121 8588
rect 23155 8585 23167 8619
rect 23109 8579 23167 8585
rect 25038 8576 25044 8628
rect 25096 8616 25102 8628
rect 25225 8619 25283 8625
rect 25225 8616 25237 8619
rect 25096 8588 25237 8616
rect 25096 8576 25102 8588
rect 25225 8585 25237 8588
rect 25271 8585 25283 8619
rect 25225 8579 25283 8585
rect 27338 8576 27344 8628
rect 27396 8576 27402 8628
rect 29270 8576 29276 8628
rect 29328 8616 29334 8628
rect 29641 8619 29699 8625
rect 29641 8616 29653 8619
rect 29328 8588 29653 8616
rect 29328 8576 29334 8588
rect 29641 8585 29653 8588
rect 29687 8585 29699 8619
rect 29641 8579 29699 8585
rect 31386 8576 31392 8628
rect 31444 8616 31450 8628
rect 31573 8619 31631 8625
rect 31573 8616 31585 8619
rect 31444 8588 31585 8616
rect 31444 8576 31450 8588
rect 31573 8585 31585 8588
rect 31619 8585 31631 8619
rect 31573 8579 31631 8585
rect 33502 8576 33508 8628
rect 33560 8616 33566 8628
rect 33689 8619 33747 8625
rect 33689 8616 33701 8619
rect 33560 8588 33701 8616
rect 33560 8576 33566 8588
rect 33689 8585 33701 8588
rect 33735 8585 33747 8619
rect 33689 8579 33747 8585
rect 35618 8576 35624 8628
rect 35676 8616 35682 8628
rect 35805 8619 35863 8625
rect 35805 8616 35817 8619
rect 35676 8588 35817 8616
rect 35676 8576 35682 8588
rect 35805 8585 35817 8588
rect 35851 8585 35863 8619
rect 35805 8579 35863 8585
rect 37734 8576 37740 8628
rect 37792 8616 37798 8628
rect 37921 8619 37979 8625
rect 37921 8616 37933 8619
rect 37792 8588 37933 8616
rect 37792 8576 37798 8588
rect 37921 8585 37933 8588
rect 37967 8585 37979 8619
rect 37921 8579 37979 8585
rect 39850 8576 39856 8628
rect 39908 8616 39914 8628
rect 40129 8619 40187 8625
rect 40129 8616 40141 8619
rect 39908 8588 40141 8616
rect 39908 8576 39914 8588
rect 40129 8585 40141 8588
rect 40175 8585 40187 8619
rect 40129 8579 40187 8585
rect 41966 8576 41972 8628
rect 42024 8616 42030 8628
rect 42613 8619 42671 8625
rect 42613 8616 42625 8619
rect 42024 8588 42625 8616
rect 42024 8576 42030 8588
rect 42613 8585 42625 8588
rect 42659 8585 42671 8619
rect 42613 8579 42671 8585
rect 43254 8576 43260 8628
rect 43312 8576 43318 8628
rect 43993 8619 44051 8625
rect 43993 8585 44005 8619
rect 44039 8585 44051 8619
rect 43993 8579 44051 8585
rect 6546 8508 6552 8560
rect 6604 8508 6610 8560
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8480 4307 8483
rect 6564 8480 6592 8508
rect 4295 8452 6592 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 2056 8412 2084 8443
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 9950 8480 9956 8492
rect 8527 8452 9956 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 11974 8480 11980 8492
rect 10643 8452 11980 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8480 12771 8483
rect 13814 8480 13820 8492
rect 12759 8452 13820 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8480 14887 8483
rect 16850 8480 16856 8492
rect 14875 8452 16856 8480
rect 14875 8449 14887 8452
rect 14829 8443 14887 8449
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 16960 8489 16988 8576
rect 19076 8489 19104 8576
rect 44008 8548 44036 8579
rect 44082 8576 44088 8628
rect 44140 8616 44146 8628
rect 44361 8619 44419 8625
rect 44361 8616 44373 8619
rect 44140 8588 44373 8616
rect 44140 8576 44146 8588
rect 44361 8585 44373 8588
rect 44407 8585 44419 8619
rect 44361 8579 44419 8585
rect 44910 8548 44916 8560
rect 24228 8520 25636 8548
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8480 21235 8483
rect 23198 8480 23204 8492
rect 21223 8452 23204 8480
rect 21223 8449 21235 8452
rect 21177 8443 21235 8449
rect 23198 8440 23204 8452
rect 23256 8440 23262 8492
rect 23290 8440 23296 8492
rect 23348 8440 23354 8492
rect 24228 8412 24256 8520
rect 25409 8483 25467 8489
rect 25409 8449 25421 8483
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 2056 8384 24256 8412
rect 25424 8344 25452 8443
rect 25608 8412 25636 8520
rect 27540 8520 39896 8548
rect 44008 8520 44916 8548
rect 27540 8489 27568 8520
rect 39868 8492 39896 8520
rect 44910 8508 44916 8520
rect 44968 8508 44974 8560
rect 27525 8483 27583 8489
rect 27525 8449 27537 8483
rect 27571 8449 27583 8483
rect 27525 8443 27583 8449
rect 29822 8440 29828 8492
rect 29880 8440 29886 8492
rect 31757 8483 31815 8489
rect 31757 8449 31769 8483
rect 31803 8480 31815 8483
rect 32398 8480 32404 8492
rect 31803 8452 32404 8480
rect 31803 8449 31815 8452
rect 31757 8443 31815 8449
rect 32398 8440 32404 8452
rect 32456 8440 32462 8492
rect 33873 8483 33931 8489
rect 33873 8449 33885 8483
rect 33919 8480 33931 8483
rect 34698 8480 34704 8492
rect 33919 8452 34704 8480
rect 33919 8449 33931 8452
rect 33873 8443 33931 8449
rect 34698 8440 34704 8452
rect 34756 8440 34762 8492
rect 35802 8440 35808 8492
rect 35860 8480 35866 8492
rect 35989 8483 36047 8489
rect 35989 8480 36001 8483
rect 35860 8452 36001 8480
rect 35860 8440 35866 8452
rect 35989 8449 36001 8452
rect 36035 8449 36047 8483
rect 35989 8443 36047 8449
rect 38105 8483 38163 8489
rect 38105 8449 38117 8483
rect 38151 8480 38163 8483
rect 38286 8480 38292 8492
rect 38151 8452 38292 8480
rect 38151 8449 38163 8452
rect 38105 8443 38163 8449
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 39850 8440 39856 8492
rect 39908 8440 39914 8492
rect 39942 8440 39948 8492
rect 40000 8440 40006 8492
rect 40862 8440 40868 8492
rect 40920 8480 40926 8492
rect 42429 8483 42487 8489
rect 42429 8480 42441 8483
rect 40920 8452 42441 8480
rect 40920 8440 40926 8452
rect 42429 8449 42441 8452
rect 42475 8449 42487 8483
rect 42429 8443 42487 8449
rect 42794 8440 42800 8492
rect 42852 8480 42858 8492
rect 43073 8483 43131 8489
rect 43073 8480 43085 8483
rect 42852 8452 43085 8480
rect 42852 8440 42858 8452
rect 43073 8449 43085 8452
rect 43119 8449 43131 8483
rect 43073 8443 43131 8449
rect 43438 8440 43444 8492
rect 43496 8440 43502 8492
rect 43806 8440 43812 8492
rect 43864 8440 43870 8492
rect 44177 8483 44235 8489
rect 44177 8449 44189 8483
rect 44223 8449 44235 8483
rect 44177 8443 44235 8449
rect 36538 8412 36544 8424
rect 25608 8384 36544 8412
rect 36538 8372 36544 8384
rect 36596 8372 36602 8424
rect 43530 8372 43536 8424
rect 43588 8412 43594 8424
rect 44192 8412 44220 8443
rect 43588 8384 44220 8412
rect 43588 8372 43594 8384
rect 40586 8344 40592 8356
rect 25424 8316 40592 8344
rect 40586 8304 40592 8316
rect 40644 8304 40650 8356
rect 43625 8347 43683 8353
rect 43625 8313 43637 8347
rect 43671 8344 43683 8347
rect 44726 8344 44732 8356
rect 43671 8316 44732 8344
rect 43671 8313 43683 8316
rect 43625 8307 43683 8313
rect 44726 8304 44732 8316
rect 44784 8304 44790 8356
rect 39758 8236 39764 8288
rect 39816 8276 39822 8288
rect 43070 8276 43076 8288
rect 39816 8248 43076 8276
rect 39816 8236 39822 8248
rect 43070 8236 43076 8248
rect 43128 8236 43134 8288
rect 1104 8186 44896 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 43950 8186
rect 44002 8134 44014 8186
rect 44066 8134 44078 8186
rect 44130 8134 44142 8186
rect 44194 8134 44206 8186
rect 44258 8134 44896 8186
rect 1104 8112 44896 8134
rect 6181 8075 6239 8081
rect 6181 8041 6193 8075
rect 6227 8072 6239 8075
rect 6730 8072 6736 8084
rect 6227 8044 6736 8072
rect 6227 8041 6239 8044
rect 6181 8035 6239 8041
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 9950 8032 9956 8084
rect 10008 8032 10014 8084
rect 11974 8032 11980 8084
rect 12032 8032 12038 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 36446 8072 36452 8084
rect 12124 8044 36452 8072
rect 12124 8032 12130 8044
rect 36446 8032 36452 8044
rect 36504 8032 36510 8084
rect 36538 8032 36544 8084
rect 36596 8032 36602 8084
rect 38105 8075 38163 8081
rect 38105 8041 38117 8075
rect 38151 8072 38163 8075
rect 38286 8072 38292 8084
rect 38151 8044 38292 8072
rect 38151 8041 38163 8044
rect 38105 8035 38163 8041
rect 38286 8032 38292 8044
rect 38344 8032 38350 8084
rect 39853 8075 39911 8081
rect 39853 8041 39865 8075
rect 39899 8072 39911 8075
rect 39942 8072 39948 8084
rect 39899 8044 39948 8072
rect 39899 8041 39911 8044
rect 39853 8035 39911 8041
rect 39942 8032 39948 8044
rect 40000 8032 40006 8084
rect 40862 8032 40868 8084
rect 40920 8032 40926 8084
rect 41598 8032 41604 8084
rect 41656 8032 41662 8084
rect 41969 8075 42027 8081
rect 41969 8041 41981 8075
rect 42015 8072 42027 8075
rect 42705 8075 42763 8081
rect 42015 8044 42564 8072
rect 42015 8041 42027 8044
rect 41969 8035 42027 8041
rect 1026 7964 1032 8016
rect 1084 8004 1090 8016
rect 42245 8007 42303 8013
rect 1084 7976 41368 8004
rect 1084 7964 1090 7976
rect 2682 7896 2688 7948
rect 2740 7896 2746 7948
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7936 3111 7939
rect 3421 7939 3479 7945
rect 3099 7908 3372 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 1360 7840 3249 7868
rect 1360 7828 1366 7840
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 3344 7868 3372 7908
rect 3421 7905 3433 7939
rect 3467 7936 3479 7939
rect 39758 7936 39764 7948
rect 3467 7908 39764 7936
rect 3467 7905 3479 7908
rect 3421 7899 3479 7905
rect 39758 7896 39764 7908
rect 39816 7896 39822 7948
rect 9861 7871 9919 7877
rect 3344 7840 7696 7868
rect 3237 7831 3295 7837
rect 750 7760 756 7812
rect 808 7800 814 7812
rect 2501 7803 2559 7809
rect 2501 7800 2513 7803
rect 808 7772 2513 7800
rect 808 7760 814 7772
rect 2501 7769 2513 7772
rect 2547 7769 2559 7803
rect 2501 7763 2559 7769
rect 2866 7760 2872 7812
rect 2924 7760 2930 7812
rect 3694 7760 3700 7812
rect 3752 7800 3758 7812
rect 6089 7803 6147 7809
rect 6089 7800 6101 7803
rect 3752 7772 6101 7800
rect 3752 7760 3758 7772
rect 6089 7769 6101 7772
rect 6135 7769 6147 7803
rect 7668 7800 7696 7840
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 10134 7868 10140 7880
rect 9907 7840 10140 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 12158 7828 12164 7880
rect 12216 7828 12222 7880
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 12066 7800 12072 7812
rect 7668 7772 12072 7800
rect 6089 7763 6147 7769
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 3602 7692 3608 7744
rect 3660 7732 3666 7744
rect 12268 7732 12296 7831
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 23566 7828 23572 7880
rect 23624 7828 23630 7880
rect 32585 7871 32643 7877
rect 32585 7837 32597 7871
rect 32631 7868 32643 7871
rect 34790 7868 34796 7880
rect 32631 7840 34796 7868
rect 32631 7837 32643 7840
rect 32585 7831 32643 7837
rect 34790 7828 34796 7840
rect 34848 7828 34854 7880
rect 34882 7828 34888 7880
rect 34940 7828 34946 7880
rect 35986 7828 35992 7880
rect 36044 7828 36050 7880
rect 36725 7871 36783 7877
rect 36725 7837 36737 7871
rect 36771 7837 36783 7871
rect 36725 7831 36783 7837
rect 38289 7871 38347 7877
rect 38289 7837 38301 7871
rect 38335 7868 38347 7871
rect 38335 7840 39436 7868
rect 38335 7837 38347 7840
rect 38289 7831 38347 7837
rect 21910 7800 21916 7812
rect 12452 7772 21916 7800
rect 12452 7741 12480 7772
rect 21910 7760 21916 7772
rect 21968 7760 21974 7812
rect 34422 7760 34428 7812
rect 34480 7800 34486 7812
rect 35437 7803 35495 7809
rect 35437 7800 35449 7803
rect 34480 7772 35449 7800
rect 34480 7760 34486 7772
rect 35437 7769 35449 7772
rect 35483 7769 35495 7803
rect 35437 7763 35495 7769
rect 35621 7803 35679 7809
rect 35621 7769 35633 7803
rect 35667 7800 35679 7803
rect 36630 7800 36636 7812
rect 35667 7772 36636 7800
rect 35667 7769 35679 7772
rect 35621 7763 35679 7769
rect 36630 7760 36636 7772
rect 36688 7760 36694 7812
rect 36740 7800 36768 7831
rect 38378 7800 38384 7812
rect 36740 7772 38384 7800
rect 38378 7760 38384 7772
rect 38436 7760 38442 7812
rect 39408 7800 39436 7840
rect 39482 7828 39488 7880
rect 39540 7828 39546 7880
rect 40034 7828 40040 7880
rect 40092 7828 40098 7880
rect 40678 7828 40684 7880
rect 40736 7828 40742 7880
rect 41340 7877 41368 7976
rect 42245 7973 42257 8007
rect 42291 7973 42303 8007
rect 42536 8004 42564 8044
rect 42705 8041 42717 8075
rect 42751 8072 42763 8075
rect 43438 8072 43444 8084
rect 42751 8044 43444 8072
rect 42751 8041 42763 8044
rect 42705 8035 42763 8041
rect 43438 8032 43444 8044
rect 43496 8032 43502 8084
rect 43714 8032 43720 8084
rect 43772 8032 43778 8084
rect 42794 8004 42800 8016
rect 42536 7976 42800 8004
rect 42245 7967 42303 7973
rect 42260 7936 42288 7967
rect 42794 7964 42800 7976
rect 42852 7964 42858 8016
rect 42981 8007 43039 8013
rect 42981 7973 42993 8007
rect 43027 7973 43039 8007
rect 42981 7967 43039 7973
rect 42260 7908 42840 7936
rect 41325 7871 41383 7877
rect 41325 7837 41337 7871
rect 41371 7837 41383 7871
rect 41325 7831 41383 7837
rect 41693 7871 41751 7877
rect 41693 7837 41705 7871
rect 41739 7868 41751 7871
rect 41785 7871 41843 7877
rect 41785 7868 41797 7871
rect 41739 7840 41797 7868
rect 41739 7837 41751 7840
rect 41693 7831 41751 7837
rect 41785 7837 41797 7840
rect 41831 7837 41843 7871
rect 41785 7831 41843 7837
rect 42058 7828 42064 7880
rect 42116 7828 42122 7880
rect 42518 7828 42524 7880
rect 42576 7828 42582 7880
rect 42812 7877 42840 7908
rect 42996 7880 43024 7967
rect 43346 7964 43352 8016
rect 43404 7964 43410 8016
rect 43070 7896 43076 7948
rect 43128 7936 43134 7948
rect 43128 7908 43944 7936
rect 43128 7896 43134 7908
rect 42797 7871 42855 7877
rect 42797 7837 42809 7871
rect 42843 7837 42855 7871
rect 42797 7831 42855 7837
rect 42978 7828 42984 7880
rect 43036 7828 43042 7880
rect 43162 7828 43168 7880
rect 43220 7828 43226 7880
rect 43916 7877 43944 7908
rect 43533 7871 43591 7877
rect 43533 7837 43545 7871
rect 43579 7837 43591 7871
rect 43533 7831 43591 7837
rect 43901 7871 43959 7877
rect 43901 7837 43913 7871
rect 43947 7837 43959 7871
rect 43901 7831 43959 7837
rect 44269 7871 44327 7877
rect 44269 7837 44281 7871
rect 44315 7868 44327 7871
rect 44542 7868 44548 7880
rect 44315 7840 44548 7868
rect 44315 7837 44327 7840
rect 44269 7831 44327 7837
rect 39666 7800 39672 7812
rect 39408 7772 39672 7800
rect 39666 7760 39672 7772
rect 39724 7760 39730 7812
rect 41524 7772 42472 7800
rect 3660 7704 12296 7732
rect 12437 7735 12495 7741
rect 3660 7692 3666 7704
rect 12437 7701 12449 7735
rect 12483 7701 12495 7735
rect 12437 7695 12495 7701
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13872 7704 14105 7732
rect 13872 7692 13878 7704
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 23753 7735 23811 7741
rect 23753 7701 23765 7735
rect 23799 7732 23811 7735
rect 27890 7732 27896 7744
rect 23799 7704 27896 7732
rect 23799 7701 23811 7704
rect 23753 7695 23811 7701
rect 27890 7692 27896 7704
rect 27948 7692 27954 7744
rect 32398 7692 32404 7744
rect 32456 7692 32462 7744
rect 34698 7692 34704 7744
rect 34756 7692 34762 7744
rect 35802 7692 35808 7744
rect 35860 7692 35866 7744
rect 37550 7692 37556 7744
rect 37608 7732 37614 7744
rect 41524 7741 41552 7772
rect 39301 7735 39359 7741
rect 39301 7732 39313 7735
rect 37608 7704 39313 7732
rect 37608 7692 37614 7704
rect 39301 7701 39313 7704
rect 39347 7701 39359 7735
rect 39301 7695 39359 7701
rect 41509 7735 41567 7741
rect 41509 7701 41521 7735
rect 41555 7701 41567 7735
rect 41509 7695 41567 7701
rect 42058 7692 42064 7744
rect 42116 7732 42122 7744
rect 42337 7735 42395 7741
rect 42337 7732 42349 7735
rect 42116 7704 42349 7732
rect 42116 7692 42122 7704
rect 42337 7701 42349 7704
rect 42383 7701 42395 7735
rect 42444 7732 42472 7772
rect 43548 7732 43576 7831
rect 44542 7828 44548 7840
rect 44600 7828 44606 7880
rect 42444 7704 43576 7732
rect 44085 7735 44143 7741
rect 42337 7695 42395 7701
rect 44085 7701 44097 7735
rect 44131 7732 44143 7735
rect 44266 7732 44272 7744
rect 44131 7704 44272 7732
rect 44131 7701 44143 7704
rect 44085 7695 44143 7701
rect 44266 7692 44272 7704
rect 44324 7692 44330 7744
rect 44450 7692 44456 7744
rect 44508 7692 44514 7744
rect 1104 7642 44896 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 44896 7642
rect 1104 7568 44896 7590
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 26329 7531 26387 7537
rect 14332 7500 26096 7528
rect 14332 7488 14338 7500
rect 12618 7420 12624 7472
rect 12676 7460 12682 7472
rect 23566 7460 23572 7472
rect 12676 7432 23572 7460
rect 12676 7420 12682 7432
rect 23566 7420 23572 7432
rect 23624 7420 23630 7472
rect 26068 7460 26096 7500
rect 26329 7497 26341 7531
rect 26375 7528 26387 7531
rect 33962 7528 33968 7540
rect 26375 7500 33968 7528
rect 26375 7497 26387 7500
rect 26329 7491 26387 7497
rect 33962 7488 33968 7500
rect 34020 7488 34026 7540
rect 34882 7488 34888 7540
rect 34940 7528 34946 7540
rect 37274 7528 37280 7540
rect 34940 7500 37280 7528
rect 34940 7488 34946 7500
rect 37274 7488 37280 7500
rect 37332 7488 37338 7540
rect 40678 7488 40684 7540
rect 40736 7528 40742 7540
rect 42702 7528 42708 7540
rect 40736 7500 42708 7528
rect 40736 7488 40742 7500
rect 42702 7488 42708 7500
rect 42760 7488 42766 7540
rect 43622 7488 43628 7540
rect 43680 7528 43686 7540
rect 44085 7531 44143 7537
rect 44085 7528 44097 7531
rect 43680 7500 44097 7528
rect 43680 7488 43686 7500
rect 44085 7497 44097 7500
rect 44131 7497 44143 7531
rect 44085 7491 44143 7497
rect 33778 7460 33784 7472
rect 26068 7432 33784 7460
rect 33778 7420 33784 7432
rect 33836 7420 33842 7472
rect 35434 7420 35440 7472
rect 35492 7420 35498 7472
rect 36630 7420 36636 7472
rect 36688 7460 36694 7472
rect 39390 7460 39396 7472
rect 36688 7432 39396 7460
rect 36688 7420 36694 7432
rect 39390 7420 39396 7432
rect 39448 7420 39454 7472
rect 39500 7432 43944 7460
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 2746 7364 12081 7392
rect 2746 7336 2774 7364
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 14369 7395 14427 7401
rect 14369 7392 14381 7395
rect 12069 7355 12127 7361
rect 12406 7364 14381 7392
rect 2682 7284 2688 7336
rect 2740 7296 2774 7336
rect 2740 7284 2746 7296
rect 3786 7284 3792 7336
rect 3844 7324 3850 7336
rect 12406 7324 12434 7364
rect 14369 7361 14381 7364
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 18230 7352 18236 7404
rect 18288 7392 18294 7404
rect 26145 7395 26203 7401
rect 26145 7392 26157 7395
rect 18288 7364 26157 7392
rect 18288 7352 18294 7364
rect 26145 7361 26157 7364
rect 26191 7361 26203 7395
rect 26145 7355 26203 7361
rect 28721 7395 28779 7401
rect 28721 7361 28733 7395
rect 28767 7392 28779 7395
rect 28813 7395 28871 7401
rect 28813 7392 28825 7395
rect 28767 7364 28825 7392
rect 28767 7361 28779 7364
rect 28721 7355 28779 7361
rect 28813 7361 28825 7364
rect 28859 7361 28871 7395
rect 28813 7355 28871 7361
rect 35621 7395 35679 7401
rect 35621 7361 35633 7395
rect 35667 7392 35679 7395
rect 38746 7392 38752 7404
rect 35667 7364 38752 7392
rect 35667 7361 35679 7364
rect 35621 7355 35679 7361
rect 38746 7352 38752 7364
rect 38804 7352 38810 7404
rect 3844 7296 12434 7324
rect 3844 7284 3850 7296
rect 36446 7284 36452 7336
rect 36504 7324 36510 7336
rect 39500 7324 39528 7432
rect 41417 7395 41475 7401
rect 41417 7361 41429 7395
rect 41463 7392 41475 7395
rect 43070 7392 43076 7404
rect 41463 7364 43076 7392
rect 41463 7361 41475 7364
rect 41417 7355 41475 7361
rect 43070 7352 43076 7364
rect 43128 7352 43134 7404
rect 43916 7401 43944 7432
rect 43809 7395 43867 7401
rect 43809 7361 43821 7395
rect 43855 7361 43867 7395
rect 43809 7355 43867 7361
rect 43901 7395 43959 7401
rect 43901 7361 43913 7395
rect 43947 7361 43959 7395
rect 43901 7355 43959 7361
rect 44269 7395 44327 7401
rect 44269 7361 44281 7395
rect 44315 7392 44327 7395
rect 44358 7392 44364 7404
rect 44315 7364 44364 7392
rect 44315 7361 44327 7364
rect 44269 7355 44327 7361
rect 36504 7296 39528 7324
rect 36504 7284 36510 7296
rect 12253 7259 12311 7265
rect 12253 7225 12265 7259
rect 12299 7256 12311 7259
rect 19702 7256 19708 7268
rect 12299 7228 19708 7256
rect 12299 7225 12311 7228
rect 12253 7219 12311 7225
rect 19702 7216 19708 7228
rect 19760 7216 19766 7268
rect 21726 7216 21732 7268
rect 21784 7256 21790 7268
rect 43824 7256 43852 7355
rect 44358 7352 44364 7364
rect 44416 7352 44422 7404
rect 21784 7228 43852 7256
rect 21784 7216 21790 7228
rect 14553 7191 14611 7197
rect 14553 7157 14565 7191
rect 14599 7188 14611 7191
rect 20530 7188 20536 7200
rect 14599 7160 20536 7188
rect 14599 7157 14611 7160
rect 14553 7151 14611 7157
rect 20530 7148 20536 7160
rect 20588 7148 20594 7200
rect 28166 7148 28172 7200
rect 28224 7188 28230 7200
rect 28629 7191 28687 7197
rect 28629 7188 28641 7191
rect 28224 7160 28641 7188
rect 28224 7148 28230 7160
rect 28629 7157 28641 7160
rect 28675 7157 28687 7191
rect 28629 7151 28687 7157
rect 28997 7191 29055 7197
rect 28997 7157 29009 7191
rect 29043 7188 29055 7191
rect 33686 7188 33692 7200
rect 29043 7160 33692 7188
rect 29043 7157 29055 7160
rect 28997 7151 29055 7157
rect 33686 7148 33692 7160
rect 33744 7148 33750 7200
rect 38562 7148 38568 7200
rect 38620 7188 38626 7200
rect 41233 7191 41291 7197
rect 41233 7188 41245 7191
rect 38620 7160 41245 7188
rect 38620 7148 38626 7160
rect 41233 7157 41245 7160
rect 41279 7157 41291 7191
rect 41233 7151 41291 7157
rect 42978 7148 42984 7200
rect 43036 7188 43042 7200
rect 43625 7191 43683 7197
rect 43625 7188 43637 7191
rect 43036 7160 43637 7188
rect 43036 7148 43042 7160
rect 43625 7157 43637 7160
rect 43671 7157 43683 7191
rect 43625 7151 43683 7157
rect 44450 7148 44456 7200
rect 44508 7148 44514 7200
rect 1104 7098 44896 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 43950 7098
rect 44002 7046 44014 7098
rect 44066 7046 44078 7098
rect 44130 7046 44142 7098
rect 44194 7046 44206 7098
rect 44258 7046 44896 7098
rect 1104 7024 44896 7046
rect 40034 6944 40040 6996
rect 40092 6984 40098 6996
rect 44910 6984 44916 6996
rect 40092 6956 44916 6984
rect 40092 6944 40098 6956
rect 44910 6944 44916 6956
rect 44968 6944 44974 6996
rect 1210 6808 1216 6860
rect 1268 6848 1274 6860
rect 2777 6851 2835 6857
rect 1268 6820 2728 6848
rect 1268 6808 1274 6820
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 1360 6752 2605 6780
rect 1360 6740 1366 6752
rect 2593 6749 2605 6752
rect 2639 6749 2651 6783
rect 2700 6780 2728 6820
rect 2777 6817 2789 6851
rect 2823 6848 2835 6851
rect 2823 6820 44312 6848
rect 2823 6817 2835 6820
rect 2777 6811 2835 6817
rect 17310 6780 17316 6792
rect 2700 6752 17316 6780
rect 2593 6743 2651 6749
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 31573 6783 31631 6789
rect 31573 6749 31585 6783
rect 31619 6780 31631 6783
rect 31665 6783 31723 6789
rect 31665 6780 31677 6783
rect 31619 6752 31677 6780
rect 31619 6749 31631 6752
rect 31573 6743 31631 6749
rect 31665 6749 31677 6752
rect 31711 6749 31723 6783
rect 31665 6743 31723 6749
rect 41417 6783 41475 6789
rect 41417 6749 41429 6783
rect 41463 6749 41475 6783
rect 41417 6743 41475 6749
rect 5534 6672 5540 6724
rect 5592 6712 5598 6724
rect 5961 6715 6019 6721
rect 5961 6712 5973 6715
rect 5592 6684 5973 6712
rect 5592 6672 5598 6684
rect 5961 6681 5973 6684
rect 6007 6681 6019 6715
rect 5961 6675 6019 6681
rect 6178 6672 6184 6724
rect 6236 6672 6242 6724
rect 41432 6712 41460 6743
rect 41506 6740 41512 6792
rect 41564 6780 41570 6792
rect 44284 6789 44312 6820
rect 43901 6783 43959 6789
rect 43901 6780 43913 6783
rect 41564 6752 43913 6780
rect 41564 6740 41570 6752
rect 43901 6749 43913 6752
rect 43947 6749 43959 6783
rect 43901 6743 43959 6749
rect 44269 6783 44327 6789
rect 44269 6749 44281 6783
rect 44315 6749 44327 6783
rect 44269 6743 44327 6749
rect 42886 6712 42892 6724
rect 41432 6684 42892 6712
rect 42886 6672 42892 6684
rect 42944 6672 42950 6724
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 18138 6644 18144 6656
rect 4212 6616 18144 6644
rect 4212 6604 4218 6616
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 28810 6604 28816 6656
rect 28868 6644 28874 6656
rect 31481 6647 31539 6653
rect 31481 6644 31493 6647
rect 28868 6616 31493 6644
rect 28868 6604 28874 6616
rect 31481 6613 31493 6616
rect 31527 6613 31539 6647
rect 31481 6607 31539 6613
rect 31849 6647 31907 6653
rect 31849 6613 31861 6647
rect 31895 6644 31907 6647
rect 33502 6644 33508 6656
rect 31895 6616 33508 6644
rect 31895 6613 31907 6616
rect 31849 6607 31907 6613
rect 33502 6604 33508 6616
rect 33560 6604 33566 6656
rect 39850 6604 39856 6656
rect 39908 6644 39914 6656
rect 41233 6647 41291 6653
rect 41233 6644 41245 6647
rect 39908 6616 41245 6644
rect 39908 6604 39914 6616
rect 41233 6613 41245 6616
rect 41279 6613 41291 6647
rect 41233 6607 41291 6613
rect 44082 6604 44088 6656
rect 44140 6604 44146 6656
rect 44450 6604 44456 6656
rect 44508 6604 44514 6656
rect 1104 6554 44896 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 44896 6554
rect 1104 6480 44896 6502
rect 6178 6400 6184 6452
rect 6236 6440 6242 6452
rect 36814 6440 36820 6452
rect 6236 6412 36820 6440
rect 6236 6400 6242 6412
rect 36814 6400 36820 6412
rect 36872 6400 36878 6452
rect 36909 6443 36967 6449
rect 36909 6409 36921 6443
rect 36955 6409 36967 6443
rect 36909 6403 36967 6409
rect 1118 6332 1124 6384
rect 1176 6372 1182 6384
rect 17954 6372 17960 6384
rect 1176 6344 17960 6372
rect 1176 6332 1182 6344
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 18506 6332 18512 6384
rect 18564 6372 18570 6384
rect 26970 6372 26976 6384
rect 18564 6344 26976 6372
rect 18564 6332 18570 6344
rect 26970 6332 26976 6344
rect 27028 6332 27034 6384
rect 4338 6264 4344 6316
rect 4396 6264 4402 6316
rect 5074 6264 5080 6316
rect 5132 6264 5138 6316
rect 18138 6264 18144 6316
rect 18196 6264 18202 6316
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 22833 6307 22891 6313
rect 22833 6304 22845 6307
rect 20496 6276 22845 6304
rect 20496 6264 20502 6276
rect 22833 6273 22845 6276
rect 22879 6304 22891 6307
rect 23017 6307 23075 6313
rect 23017 6304 23029 6307
rect 22879 6276 23029 6304
rect 22879 6273 22891 6276
rect 22833 6267 22891 6273
rect 23017 6273 23029 6276
rect 23063 6273 23075 6307
rect 23017 6267 23075 6273
rect 25777 6307 25835 6313
rect 25777 6273 25789 6307
rect 25823 6273 25835 6307
rect 25777 6267 25835 6273
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 25792 6236 25820 6267
rect 32858 6264 32864 6316
rect 32916 6304 32922 6316
rect 36924 6304 36952 6403
rect 37734 6400 37740 6452
rect 37792 6440 37798 6452
rect 38197 6443 38255 6449
rect 38197 6440 38209 6443
rect 37792 6412 38209 6440
rect 37792 6400 37798 6412
rect 38197 6409 38209 6412
rect 38243 6409 38255 6443
rect 38197 6403 38255 6409
rect 40678 6400 40684 6452
rect 40736 6400 40742 6452
rect 43073 6443 43131 6449
rect 43073 6409 43085 6443
rect 43119 6440 43131 6443
rect 43806 6440 43812 6452
rect 43119 6412 43812 6440
rect 43119 6409 43131 6412
rect 43073 6403 43131 6409
rect 43806 6400 43812 6412
rect 43864 6400 43870 6452
rect 44450 6400 44456 6452
rect 44508 6400 44514 6452
rect 41598 6372 41604 6384
rect 38396 6344 41604 6372
rect 38396 6313 38424 6344
rect 41598 6332 41604 6344
rect 41656 6332 41662 6384
rect 32916 6276 36952 6304
rect 37093 6307 37151 6313
rect 32916 6264 32922 6276
rect 37093 6273 37105 6307
rect 37139 6304 37151 6307
rect 37461 6307 37519 6313
rect 37139 6276 37412 6304
rect 37139 6273 37151 6276
rect 37093 6267 37151 6273
rect 12308 6208 25820 6236
rect 12308 6196 12314 6208
rect 4522 6128 4528 6180
rect 4580 6128 4586 6180
rect 12158 6128 12164 6180
rect 12216 6168 12222 6180
rect 23106 6168 23112 6180
rect 12216 6140 23112 6168
rect 12216 6128 12222 6140
rect 23106 6128 23112 6140
rect 23164 6128 23170 6180
rect 23201 6171 23259 6177
rect 23201 6137 23213 6171
rect 23247 6168 23259 6171
rect 27338 6168 27344 6180
rect 23247 6140 27344 6168
rect 23247 6137 23259 6140
rect 23201 6131 23259 6137
rect 27338 6128 27344 6140
rect 27396 6128 27402 6180
rect 37277 6171 37335 6177
rect 37277 6168 37289 6171
rect 36556 6140 37289 6168
rect 5166 6060 5172 6112
rect 5224 6060 5230 6112
rect 18325 6103 18383 6109
rect 18325 6069 18337 6103
rect 18371 6100 18383 6103
rect 20622 6100 20628 6112
rect 18371 6072 20628 6100
rect 18371 6069 18383 6072
rect 18325 6063 18383 6069
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 25961 6103 26019 6109
rect 25961 6069 25973 6103
rect 26007 6100 26019 6103
rect 26786 6100 26792 6112
rect 26007 6072 26792 6100
rect 26007 6069 26019 6072
rect 25961 6063 26019 6069
rect 26786 6060 26792 6072
rect 26844 6060 26850 6112
rect 34330 6060 34336 6112
rect 34388 6100 34394 6112
rect 36556 6100 36584 6140
rect 37277 6137 37289 6140
rect 37323 6137 37335 6171
rect 37277 6131 37335 6137
rect 34388 6072 36584 6100
rect 37384 6100 37412 6276
rect 37461 6273 37473 6307
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 38381 6307 38439 6313
rect 38381 6273 38393 6307
rect 38427 6273 38439 6307
rect 38381 6267 38439 6273
rect 39577 6307 39635 6313
rect 39577 6273 39589 6307
rect 39623 6273 39635 6307
rect 39577 6267 39635 6273
rect 40865 6307 40923 6313
rect 40865 6273 40877 6307
rect 40911 6304 40923 6307
rect 42334 6304 42340 6316
rect 40911 6276 42340 6304
rect 40911 6273 40923 6276
rect 40865 6267 40923 6273
rect 37476 6236 37504 6267
rect 39592 6236 39620 6267
rect 42334 6264 42340 6276
rect 42392 6264 42398 6316
rect 42794 6264 42800 6316
rect 42852 6304 42858 6316
rect 42889 6307 42947 6313
rect 42889 6304 42901 6307
rect 42852 6276 42901 6304
rect 42852 6264 42858 6276
rect 42889 6273 42901 6276
rect 42935 6273 42947 6307
rect 43901 6307 43959 6313
rect 43901 6304 43913 6307
rect 42889 6267 42947 6273
rect 42996 6276 43913 6304
rect 42058 6236 42064 6248
rect 37476 6208 39528 6236
rect 39592 6208 42064 6236
rect 37458 6128 37464 6180
rect 37516 6168 37522 6180
rect 39393 6171 39451 6177
rect 39393 6168 39405 6171
rect 37516 6140 39405 6168
rect 37516 6128 37522 6140
rect 39393 6137 39405 6140
rect 39439 6137 39451 6171
rect 39500 6168 39528 6208
rect 42058 6196 42064 6208
rect 42116 6196 42122 6248
rect 41322 6168 41328 6180
rect 39500 6140 41328 6168
rect 39393 6131 39451 6137
rect 41322 6128 41328 6140
rect 41380 6128 41386 6180
rect 40954 6100 40960 6112
rect 37384 6072 40960 6100
rect 34388 6060 34394 6072
rect 40954 6060 40960 6072
rect 41012 6060 41018 6112
rect 41046 6060 41052 6112
rect 41104 6100 41110 6112
rect 42996 6100 43024 6276
rect 43901 6273 43913 6276
rect 43947 6273 43959 6307
rect 43901 6267 43959 6273
rect 44269 6307 44327 6313
rect 44269 6273 44281 6307
rect 44315 6273 44327 6307
rect 44269 6267 44327 6273
rect 43254 6196 43260 6248
rect 43312 6236 43318 6248
rect 44284 6236 44312 6267
rect 43312 6208 44312 6236
rect 43312 6196 43318 6208
rect 44082 6128 44088 6180
rect 44140 6128 44146 6180
rect 41104 6072 43024 6100
rect 41104 6060 41110 6072
rect 1104 6010 44896 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 43950 6010
rect 44002 5958 44014 6010
rect 44066 5958 44078 6010
rect 44130 5958 44142 6010
rect 44194 5958 44206 6010
rect 44258 5958 44896 6010
rect 1104 5936 44896 5958
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 37182 5896 37188 5908
rect 5224 5868 37188 5896
rect 5224 5856 5230 5868
rect 37182 5856 37188 5868
rect 37240 5856 37246 5908
rect 39666 5856 39672 5908
rect 39724 5896 39730 5908
rect 44634 5896 44640 5908
rect 39724 5868 44640 5896
rect 39724 5856 39730 5868
rect 44634 5856 44640 5868
rect 44692 5856 44698 5908
rect 6086 5788 6092 5840
rect 6144 5828 6150 5840
rect 16482 5828 16488 5840
rect 6144 5800 16488 5828
rect 6144 5788 6150 5800
rect 16482 5788 16488 5800
rect 16540 5788 16546 5840
rect 16666 5788 16672 5840
rect 16724 5828 16730 5840
rect 27157 5831 27215 5837
rect 16724 5800 22416 5828
rect 16724 5788 16730 5800
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 2271 5732 2774 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 1026 5652 1032 5704
rect 1084 5692 1090 5704
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 1084 5664 2053 5692
rect 1084 5652 1090 5664
rect 2041 5661 2053 5664
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2746 5624 2774 5732
rect 16684 5732 22094 5760
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 16301 5695 16359 5701
rect 16301 5692 16313 5695
rect 7156 5664 16313 5692
rect 7156 5652 7162 5664
rect 16301 5661 16313 5664
rect 16347 5661 16359 5695
rect 16684 5692 16712 5732
rect 16301 5655 16359 5661
rect 16408 5664 16712 5692
rect 16761 5695 16819 5701
rect 16408 5624 16436 5664
rect 16761 5661 16773 5695
rect 16807 5692 16819 5695
rect 16807 5664 21680 5692
rect 16807 5661 16819 5664
rect 16761 5655 16819 5661
rect 16850 5624 16856 5636
rect 2746 5596 16436 5624
rect 16592 5596 16856 5624
rect 16482 5516 16488 5568
rect 16540 5516 16546 5568
rect 16592 5565 16620 5596
rect 16850 5584 16856 5596
rect 16908 5584 16914 5636
rect 16577 5559 16635 5565
rect 16577 5525 16589 5559
rect 16623 5525 16635 5559
rect 16577 5519 16635 5525
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 21450 5556 21456 5568
rect 16724 5528 21456 5556
rect 16724 5516 16730 5528
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 21652 5556 21680 5664
rect 22066 5624 22094 5732
rect 22388 5701 22416 5800
rect 27157 5797 27169 5831
rect 27203 5828 27215 5831
rect 32766 5828 32772 5840
rect 27203 5800 32772 5828
rect 27203 5797 27215 5800
rect 27157 5791 27215 5797
rect 32766 5788 32772 5800
rect 32824 5788 32830 5840
rect 36814 5788 36820 5840
rect 36872 5828 36878 5840
rect 36872 5800 43300 5828
rect 36872 5788 36878 5800
rect 23106 5720 23112 5772
rect 23164 5760 23170 5772
rect 31110 5760 31116 5772
rect 23164 5732 31116 5760
rect 23164 5720 23170 5732
rect 31110 5720 31116 5732
rect 31168 5720 31174 5772
rect 41506 5760 41512 5772
rect 35866 5732 41512 5760
rect 22373 5695 22431 5701
rect 22373 5661 22385 5695
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 26970 5652 26976 5704
rect 27028 5652 27034 5704
rect 31573 5695 31631 5701
rect 31573 5661 31585 5695
rect 31619 5692 31631 5695
rect 31665 5695 31723 5701
rect 31665 5692 31677 5695
rect 31619 5664 31677 5692
rect 31619 5661 31631 5664
rect 31573 5655 31631 5661
rect 31665 5661 31677 5664
rect 31711 5661 31723 5695
rect 31665 5655 31723 5661
rect 35866 5624 35894 5732
rect 41506 5720 41512 5732
rect 41564 5720 41570 5772
rect 43162 5720 43168 5772
rect 43220 5720 43226 5772
rect 43272 5760 43300 5800
rect 44450 5788 44456 5840
rect 44508 5788 44514 5840
rect 44818 5760 44824 5772
rect 43272 5732 44824 5760
rect 44818 5720 44824 5732
rect 44876 5720 44882 5772
rect 43257 5695 43315 5701
rect 43257 5661 43269 5695
rect 43303 5692 43315 5695
rect 43349 5695 43407 5701
rect 43349 5692 43361 5695
rect 43303 5664 43361 5692
rect 43303 5661 43315 5664
rect 43257 5655 43315 5661
rect 43349 5661 43361 5664
rect 43395 5661 43407 5695
rect 43901 5695 43959 5701
rect 43901 5692 43913 5695
rect 43349 5655 43407 5661
rect 43456 5664 43913 5692
rect 22066 5596 35894 5624
rect 41414 5584 41420 5636
rect 41472 5624 41478 5636
rect 43456 5624 43484 5664
rect 43901 5661 43913 5664
rect 43947 5661 43959 5695
rect 43901 5655 43959 5661
rect 44269 5695 44327 5701
rect 44269 5661 44281 5695
rect 44315 5661 44327 5695
rect 44269 5655 44327 5661
rect 44284 5624 44312 5655
rect 41472 5596 43484 5624
rect 43548 5596 44312 5624
rect 41472 5584 41478 5596
rect 22370 5556 22376 5568
rect 21652 5528 22376 5556
rect 22370 5516 22376 5528
rect 22428 5516 22434 5568
rect 22557 5559 22615 5565
rect 22557 5525 22569 5559
rect 22603 5556 22615 5559
rect 25130 5556 25136 5568
rect 22603 5528 25136 5556
rect 22603 5525 22615 5528
rect 22557 5519 22615 5525
rect 25130 5516 25136 5528
rect 25188 5516 25194 5568
rect 31478 5516 31484 5568
rect 31536 5516 31542 5568
rect 31849 5559 31907 5565
rect 31849 5525 31861 5559
rect 31895 5556 31907 5559
rect 34422 5556 34428 5568
rect 31895 5528 34428 5556
rect 31895 5525 31907 5528
rect 31849 5519 31907 5525
rect 34422 5516 34428 5528
rect 34480 5516 34486 5568
rect 43548 5565 43576 5596
rect 43533 5559 43591 5565
rect 43533 5525 43545 5559
rect 43579 5525 43591 5559
rect 43533 5519 43591 5525
rect 44085 5559 44143 5565
rect 44085 5525 44097 5559
rect 44131 5556 44143 5559
rect 45186 5556 45192 5568
rect 44131 5528 45192 5556
rect 44131 5525 44143 5528
rect 44085 5519 44143 5525
rect 45186 5516 45192 5528
rect 45244 5516 45250 5568
rect 1104 5466 44896 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 44896 5466
rect 1104 5392 44896 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 17218 5352 17224 5364
rect 4120 5324 17224 5352
rect 4120 5312 4126 5324
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 17310 5312 17316 5364
rect 17368 5352 17374 5364
rect 17368 5324 31754 5352
rect 17368 5312 17374 5324
rect 1302 5244 1308 5296
rect 1360 5284 1366 5296
rect 3053 5287 3111 5293
rect 3053 5284 3065 5287
rect 1360 5256 3065 5284
rect 1360 5244 1366 5256
rect 3053 5253 3065 5256
rect 3099 5253 3111 5287
rect 3053 5247 3111 5253
rect 4522 5244 4528 5296
rect 4580 5284 4586 5296
rect 31726 5284 31754 5324
rect 37182 5312 37188 5364
rect 37240 5352 37246 5364
rect 37240 5324 42564 5352
rect 37240 5312 37246 5324
rect 42536 5284 42564 5324
rect 43254 5312 43260 5364
rect 43312 5312 43318 5364
rect 44450 5312 44456 5364
rect 44508 5312 44514 5364
rect 4580 5256 16252 5284
rect 4580 5244 4586 5256
rect 6362 5176 6368 5228
rect 6420 5216 6426 5228
rect 15930 5216 15936 5228
rect 6420 5188 15936 5216
rect 6420 5176 6426 5188
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16022 5176 16028 5228
rect 16080 5176 16086 5228
rect 16224 5216 16252 5256
rect 19306 5256 31616 5284
rect 31726 5256 42472 5284
rect 42536 5256 43944 5284
rect 19306 5216 19334 5256
rect 16224 5188 19334 5216
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5185 20499 5219
rect 31481 5219 31539 5225
rect 31481 5216 31493 5219
rect 20441 5179 20499 5185
rect 22066 5188 31493 5216
rect 3234 5108 3240 5160
rect 3292 5108 3298 5160
rect 16114 5108 16120 5160
rect 16172 5148 16178 5160
rect 19518 5148 19524 5160
rect 16172 5120 19524 5148
rect 16172 5108 16178 5120
rect 19518 5108 19524 5120
rect 19576 5108 19582 5160
rect 16298 5040 16304 5092
rect 16356 5080 16362 5092
rect 20456 5080 20484 5179
rect 22066 5148 22094 5188
rect 31481 5185 31493 5188
rect 31527 5185 31539 5219
rect 31481 5179 31539 5185
rect 16356 5052 20484 5080
rect 20548 5120 22094 5148
rect 31588 5148 31616 5256
rect 42444 5225 42472 5256
rect 43916 5225 43944 5256
rect 42429 5219 42487 5225
rect 42429 5185 42441 5219
rect 42475 5216 42487 5219
rect 42705 5219 42763 5225
rect 42705 5216 42717 5219
rect 42475 5188 42717 5216
rect 42475 5185 42487 5188
rect 42429 5179 42487 5185
rect 42705 5185 42717 5188
rect 42751 5185 42763 5219
rect 42705 5179 42763 5185
rect 42981 5219 43039 5225
rect 42981 5185 42993 5219
rect 43027 5216 43039 5219
rect 43073 5219 43131 5225
rect 43073 5216 43085 5219
rect 43027 5188 43085 5216
rect 43027 5185 43039 5188
rect 42981 5179 43039 5185
rect 43073 5185 43085 5188
rect 43119 5185 43131 5219
rect 43073 5179 43131 5185
rect 43901 5219 43959 5225
rect 43901 5185 43913 5219
rect 43947 5185 43959 5219
rect 43901 5179 43959 5185
rect 44269 5219 44327 5225
rect 44269 5185 44281 5219
rect 44315 5185 44327 5219
rect 44269 5179 44327 5185
rect 44284 5148 44312 5179
rect 31588 5120 44312 5148
rect 16356 5040 16362 5052
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 16114 5012 16120 5024
rect 6512 4984 16120 5012
rect 6512 4972 6518 4984
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 16206 4972 16212 5024
rect 16264 4972 16270 5024
rect 16666 4972 16672 5024
rect 16724 5012 16730 5024
rect 20548 5012 20576 5120
rect 22462 5040 22468 5092
rect 22520 5080 22526 5092
rect 42889 5083 42947 5089
rect 42889 5080 42901 5083
rect 22520 5052 42901 5080
rect 22520 5040 22526 5052
rect 42889 5049 42901 5052
rect 42935 5049 42947 5083
rect 42889 5043 42947 5049
rect 44082 5040 44088 5092
rect 44140 5040 44146 5092
rect 16724 4984 20576 5012
rect 20625 5015 20683 5021
rect 16724 4972 16730 4984
rect 20625 4981 20637 5015
rect 20671 5012 20683 5015
rect 23382 5012 23388 5024
rect 20671 4984 23388 5012
rect 20671 4981 20683 4984
rect 20625 4975 20683 4981
rect 23382 4972 23388 4984
rect 23440 4972 23446 5024
rect 31665 5015 31723 5021
rect 31665 4981 31677 5015
rect 31711 5012 31723 5015
rect 33870 5012 33876 5024
rect 31711 4984 33876 5012
rect 31711 4981 31723 4984
rect 31665 4975 31723 4981
rect 33870 4972 33876 4984
rect 33928 4972 33934 5024
rect 42613 5015 42671 5021
rect 42613 4981 42625 5015
rect 42659 5012 42671 5015
rect 44542 5012 44548 5024
rect 42659 4984 44548 5012
rect 42659 4981 42671 4984
rect 42613 4975 42671 4981
rect 44542 4972 44548 4984
rect 44600 4972 44606 5024
rect 1104 4922 44896 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 43950 4922
rect 44002 4870 44014 4922
rect 44066 4870 44078 4922
rect 44130 4870 44142 4922
rect 44194 4870 44206 4922
rect 44258 4870 44896 4922
rect 1104 4848 44896 4870
rect 4522 4768 4528 4820
rect 4580 4808 4586 4820
rect 11882 4808 11888 4820
rect 4580 4780 11888 4808
rect 4580 4768 4586 4780
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 11992 4780 12434 4808
rect 3418 4700 3424 4752
rect 3476 4740 3482 4752
rect 11992 4740 12020 4780
rect 3476 4712 12020 4740
rect 12406 4740 12434 4780
rect 16206 4768 16212 4820
rect 16264 4808 16270 4820
rect 30282 4808 30288 4820
rect 16264 4780 30288 4808
rect 16264 4768 16270 4780
rect 30282 4768 30288 4780
rect 30340 4768 30346 4820
rect 43530 4768 43536 4820
rect 43588 4808 43594 4820
rect 43809 4811 43867 4817
rect 43809 4808 43821 4811
rect 43588 4780 43821 4808
rect 43588 4768 43594 4780
rect 43809 4777 43821 4780
rect 43855 4777 43867 4811
rect 43809 4771 43867 4777
rect 22278 4740 22284 4752
rect 12406 4712 22284 4740
rect 3476 4700 3482 4712
rect 22278 4700 22284 4712
rect 22336 4700 22342 4752
rect 42797 4743 42855 4749
rect 42797 4709 42809 4743
rect 42843 4740 42855 4743
rect 44358 4740 44364 4752
rect 42843 4712 44364 4740
rect 42843 4709 42855 4712
rect 42797 4703 42855 4709
rect 44358 4700 44364 4712
rect 44416 4700 44422 4752
rect 44450 4700 44456 4752
rect 44508 4700 44514 4752
rect 474 4632 480 4684
rect 532 4672 538 4684
rect 532 4644 7144 4672
rect 532 4632 538 4644
rect 658 4564 664 4616
rect 716 4604 722 4616
rect 7116 4613 7144 4644
rect 7742 4632 7748 4684
rect 7800 4672 7806 4684
rect 7800 4644 12020 4672
rect 7800 4632 7806 4644
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 716 4576 2145 4604
rect 716 4564 722 4576
rect 2133 4573 2145 4576
rect 2179 4573 2191 4607
rect 6273 4607 6331 4613
rect 6273 4604 6285 4607
rect 2133 4567 2191 4573
rect 2240 4576 6285 4604
rect 842 4496 848 4548
rect 900 4536 906 4548
rect 2240 4536 2268 4576
rect 6273 4573 6285 4576
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 900 4508 2268 4536
rect 900 4496 906 4508
rect 2314 4496 2320 4548
rect 2372 4496 2378 4548
rect 4890 4496 4896 4548
rect 4948 4536 4954 4548
rect 6656 4536 6684 4567
rect 10870 4564 10876 4616
rect 10928 4564 10934 4616
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4573 11943 4607
rect 11992 4604 12020 4644
rect 12066 4632 12072 4684
rect 12124 4672 12130 4684
rect 23201 4675 23259 4681
rect 23201 4672 23213 4675
rect 12124 4644 23213 4672
rect 12124 4632 12130 4644
rect 23201 4641 23213 4644
rect 23247 4641 23259 4675
rect 23201 4635 23259 4641
rect 42426 4632 42432 4684
rect 42484 4632 42490 4684
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 11992 4576 12817 4604
rect 11885 4567 11943 4573
rect 12805 4573 12817 4576
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 4948 4508 6684 4536
rect 4948 4496 4954 4508
rect 7466 4496 7472 4548
rect 7524 4536 7530 4548
rect 11900 4536 11928 4567
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13872 4576 14105 4604
rect 13872 4564 13878 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 16390 4564 16396 4616
rect 16448 4564 16454 4616
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 23293 4607 23351 4613
rect 17276 4576 22094 4604
rect 17276 4564 17282 4576
rect 15930 4536 15936 4548
rect 7524 4508 11928 4536
rect 13004 4508 15936 4536
rect 7524 4496 7530 4508
rect 6454 4428 6460 4480
rect 6512 4428 6518 4480
rect 6825 4471 6883 4477
rect 6825 4437 6837 4471
rect 6871 4468 6883 4471
rect 7190 4468 7196 4480
rect 6871 4440 7196 4468
rect 6871 4437 6883 4440
rect 6825 4431 6883 4437
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 7282 4428 7288 4480
rect 7340 4428 7346 4480
rect 11054 4428 11060 4480
rect 11112 4428 11118 4480
rect 12066 4428 12072 4480
rect 12124 4428 12130 4480
rect 13004 4477 13032 4508
rect 15930 4496 15936 4508
rect 15988 4496 15994 4548
rect 17586 4536 17592 4548
rect 16500 4508 17592 4536
rect 12989 4471 13047 4477
rect 12989 4437 13001 4471
rect 13035 4437 13047 4471
rect 12989 4431 13047 4437
rect 14277 4471 14335 4477
rect 14277 4437 14289 4471
rect 14323 4468 14335 4471
rect 16500 4468 16528 4508
rect 17586 4496 17592 4508
rect 17644 4496 17650 4548
rect 22066 4536 22094 4576
rect 23293 4573 23305 4607
rect 23339 4604 23351 4607
rect 23385 4607 23443 4613
rect 23385 4604 23397 4607
rect 23339 4576 23397 4604
rect 23339 4573 23351 4576
rect 23293 4567 23351 4573
rect 23385 4573 23397 4576
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 38654 4564 38660 4616
rect 38712 4604 38718 4616
rect 39301 4607 39359 4613
rect 39301 4604 39313 4607
rect 38712 4576 39313 4604
rect 38712 4564 38718 4576
rect 39301 4573 39313 4576
rect 39347 4573 39359 4607
rect 39301 4567 39359 4573
rect 41141 4607 41199 4613
rect 41141 4573 41153 4607
rect 41187 4604 41199 4607
rect 41417 4607 41475 4613
rect 41417 4604 41429 4607
rect 41187 4576 41429 4604
rect 41187 4573 41199 4576
rect 41141 4567 41199 4573
rect 41417 4573 41429 4576
rect 41463 4573 41475 4607
rect 41417 4567 41475 4573
rect 42521 4607 42579 4613
rect 42521 4573 42533 4607
rect 42567 4604 42579 4607
rect 42613 4607 42671 4613
rect 42613 4604 42625 4607
rect 42567 4576 42625 4604
rect 42567 4573 42579 4576
rect 42521 4567 42579 4573
rect 42613 4573 42625 4576
rect 42659 4573 42671 4607
rect 42613 4567 42671 4573
rect 43625 4607 43683 4613
rect 43625 4573 43637 4607
rect 43671 4573 43683 4607
rect 43625 4567 43683 4573
rect 25590 4536 25596 4548
rect 22066 4508 25596 4536
rect 25590 4496 25596 4508
rect 25648 4496 25654 4548
rect 43640 4536 43668 4567
rect 43898 4564 43904 4616
rect 43956 4564 43962 4616
rect 44269 4607 44327 4613
rect 44269 4573 44281 4607
rect 44315 4604 44327 4607
rect 44818 4604 44824 4616
rect 44315 4576 44824 4604
rect 44315 4573 44327 4576
rect 44269 4567 44327 4573
rect 44818 4564 44824 4576
rect 44876 4564 44882 4616
rect 45738 4536 45744 4548
rect 43640 4508 45744 4536
rect 45738 4496 45744 4508
rect 45796 4496 45802 4548
rect 14323 4440 16528 4468
rect 16577 4471 16635 4477
rect 14323 4437 14335 4440
rect 14277 4431 14335 4437
rect 16577 4437 16589 4471
rect 16623 4468 16635 4471
rect 17678 4468 17684 4480
rect 16623 4440 17684 4468
rect 16623 4437 16635 4440
rect 16577 4431 16635 4437
rect 17678 4428 17684 4440
rect 17736 4428 17742 4480
rect 23569 4471 23627 4477
rect 23569 4437 23581 4471
rect 23615 4468 23627 4471
rect 24946 4468 24952 4480
rect 23615 4440 24952 4468
rect 23615 4437 23627 4440
rect 23569 4431 23627 4437
rect 24946 4428 24952 4440
rect 25004 4428 25010 4480
rect 38838 4428 38844 4480
rect 38896 4468 38902 4480
rect 39117 4471 39175 4477
rect 39117 4468 39129 4471
rect 38896 4440 39129 4468
rect 38896 4428 38902 4440
rect 39117 4437 39129 4440
rect 39163 4437 39175 4471
rect 39117 4431 39175 4437
rect 41046 4428 41052 4480
rect 41104 4428 41110 4480
rect 41230 4428 41236 4480
rect 41288 4428 41294 4480
rect 44082 4428 44088 4480
rect 44140 4428 44146 4480
rect 1104 4378 44896 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 44896 4378
rect 1104 4304 44896 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 10870 4264 10876 4276
rect 2464 4236 10876 4264
rect 2464 4224 2470 4236
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 43349 4267 43407 4273
rect 43349 4233 43361 4267
rect 43395 4264 43407 4267
rect 43898 4264 43904 4276
rect 43395 4236 43904 4264
rect 43395 4233 43407 4236
rect 43349 4227 43407 4233
rect 43898 4224 43904 4236
rect 43956 4224 43962 4276
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 16390 4196 16396 4208
rect 9732 4168 16396 4196
rect 9732 4156 9738 4168
rect 16390 4156 16396 4168
rect 16448 4156 16454 4208
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 1912 4100 4997 4128
rect 1912 4088 1918 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 5316 4100 7665 4128
rect 5316 4088 5322 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 5626 4020 5632 4072
rect 5684 4060 5690 4072
rect 9876 4060 9904 4091
rect 20898 4088 20904 4140
rect 20956 4128 20962 4140
rect 27065 4131 27123 4137
rect 27065 4128 27077 4131
rect 20956 4100 27077 4128
rect 20956 4088 20962 4100
rect 27065 4097 27077 4100
rect 27111 4097 27123 4131
rect 27065 4091 27123 4097
rect 38562 4088 38568 4140
rect 38620 4088 38626 4140
rect 43073 4131 43131 4137
rect 43073 4097 43085 4131
rect 43119 4128 43131 4131
rect 43165 4131 43223 4137
rect 43165 4128 43177 4131
rect 43119 4100 43177 4128
rect 43119 4097 43131 4100
rect 43073 4091 43131 4097
rect 43165 4097 43177 4100
rect 43211 4097 43223 4131
rect 43165 4091 43223 4097
rect 43438 4088 43444 4140
rect 43496 4128 43502 4140
rect 43901 4131 43959 4137
rect 43901 4128 43913 4131
rect 43496 4100 43913 4128
rect 43496 4088 43502 4100
rect 43901 4097 43913 4100
rect 43947 4097 43959 4131
rect 43901 4091 43959 4097
rect 44269 4131 44327 4137
rect 44269 4097 44281 4131
rect 44315 4097 44327 4131
rect 44269 4091 44327 4097
rect 5684 4032 9904 4060
rect 5684 4020 5690 4032
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 19610 4060 19616 4072
rect 10008 4032 19616 4060
rect 10008 4020 10014 4032
rect 19610 4020 19616 4032
rect 19668 4020 19674 4072
rect 22370 4020 22376 4072
rect 22428 4060 22434 4072
rect 35066 4060 35072 4072
rect 22428 4032 35072 4060
rect 22428 4020 22434 4032
rect 35066 4020 35072 4032
rect 35124 4020 35130 4072
rect 43254 4020 43260 4072
rect 43312 4060 43318 4072
rect 44284 4060 44312 4091
rect 43312 4032 44312 4060
rect 43312 4020 43318 4032
rect 750 3952 756 4004
rect 808 3992 814 4004
rect 42981 3995 43039 4001
rect 42981 3992 42993 3995
rect 808 3964 42993 3992
rect 808 3952 814 3964
rect 42981 3961 42993 3964
rect 43027 3961 43039 3995
rect 42981 3955 43039 3961
rect 44082 3952 44088 4004
rect 44140 3952 44146 4004
rect 44450 3952 44456 4004
rect 44508 3952 44514 4004
rect 5169 3927 5227 3933
rect 5169 3893 5181 3927
rect 5215 3924 5227 3927
rect 6178 3924 6184 3936
rect 5215 3896 6184 3924
rect 5215 3893 5227 3896
rect 5169 3887 5227 3893
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 7834 3884 7840 3936
rect 7892 3884 7898 3936
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 14642 3924 14648 3936
rect 10091 3896 14648 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 27249 3927 27307 3933
rect 27249 3893 27261 3927
rect 27295 3924 27307 3927
rect 27430 3924 27436 3936
rect 27295 3896 27436 3924
rect 27295 3893 27307 3896
rect 27249 3887 27307 3893
rect 27430 3884 27436 3896
rect 27488 3884 27494 3936
rect 38381 3927 38439 3933
rect 38381 3893 38393 3927
rect 38427 3924 38439 3927
rect 38470 3924 38476 3936
rect 38427 3896 38476 3924
rect 38427 3893 38439 3896
rect 38381 3887 38439 3893
rect 38470 3884 38476 3896
rect 38528 3884 38534 3936
rect 1104 3834 44896 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 43950 3834
rect 44002 3782 44014 3834
rect 44066 3782 44078 3834
rect 44130 3782 44142 3834
rect 44194 3782 44206 3834
rect 44258 3782 44896 3834
rect 1104 3760 44896 3782
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 14366 3720 14372 3732
rect 7892 3692 14372 3720
rect 7892 3680 7898 3692
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 17129 3723 17187 3729
rect 17129 3689 17141 3723
rect 17175 3720 17187 3723
rect 34514 3720 34520 3732
rect 17175 3692 34520 3720
rect 17175 3689 17187 3692
rect 17129 3683 17187 3689
rect 34514 3680 34520 3692
rect 34572 3680 34578 3732
rect 34885 3723 34943 3729
rect 34885 3689 34897 3723
rect 34931 3720 34943 3723
rect 36538 3720 36544 3732
rect 34931 3692 36544 3720
rect 34931 3689 34943 3692
rect 34885 3683 34943 3689
rect 36538 3680 36544 3692
rect 36596 3680 36602 3732
rect 43073 3723 43131 3729
rect 43073 3689 43085 3723
rect 43119 3720 43131 3723
rect 43254 3720 43260 3732
rect 43119 3692 43260 3720
rect 43119 3689 43131 3692
rect 43073 3683 43131 3689
rect 43254 3680 43260 3692
rect 43312 3680 43318 3732
rect 1302 3612 1308 3664
rect 1360 3652 1366 3664
rect 42797 3655 42855 3661
rect 42797 3652 42809 3655
rect 1360 3624 42809 3652
rect 1360 3612 1366 3624
rect 42797 3621 42809 3624
rect 42843 3621 42855 3655
rect 42797 3615 42855 3621
rect 44450 3612 44456 3664
rect 44508 3612 44514 3664
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 43346 3584 43352 3596
rect 2372 3556 43352 3584
rect 2372 3544 2378 3556
rect 43346 3544 43352 3556
rect 43404 3544 43410 3596
rect 6730 3476 6736 3528
rect 6788 3516 6794 3528
rect 9950 3516 9956 3528
rect 6788 3488 9956 3516
rect 6788 3476 6794 3488
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 16574 3476 16580 3528
rect 16632 3476 16638 3528
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 14458 3408 14464 3460
rect 14516 3448 14522 3460
rect 16960 3448 16988 3479
rect 18690 3476 18696 3528
rect 18748 3476 18754 3528
rect 19610 3476 19616 3528
rect 19668 3476 19674 3528
rect 27709 3519 27767 3525
rect 27709 3485 27721 3519
rect 27755 3516 27767 3519
rect 27801 3519 27859 3525
rect 27801 3516 27813 3519
rect 27755 3488 27813 3516
rect 27755 3485 27767 3488
rect 27709 3479 27767 3485
rect 27801 3485 27813 3488
rect 27847 3485 27859 3519
rect 27801 3479 27859 3485
rect 28353 3519 28411 3525
rect 28353 3485 28365 3519
rect 28399 3516 28411 3519
rect 28445 3519 28503 3525
rect 28445 3516 28457 3519
rect 28399 3488 28457 3516
rect 28399 3485 28411 3488
rect 28353 3479 28411 3485
rect 28445 3485 28457 3488
rect 28491 3485 28503 3519
rect 28445 3479 28503 3485
rect 28905 3519 28963 3525
rect 28905 3485 28917 3519
rect 28951 3516 28963 3519
rect 28997 3519 29055 3525
rect 28997 3516 29009 3519
rect 28951 3488 29009 3516
rect 28951 3485 28963 3488
rect 28905 3479 28963 3485
rect 28997 3485 29009 3488
rect 29043 3485 29055 3519
rect 28997 3479 29055 3485
rect 29086 3476 29092 3528
rect 29144 3516 29150 3528
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 29144 3488 29561 3516
rect 29144 3476 29150 3488
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 34606 3476 34612 3528
rect 34664 3516 34670 3528
rect 34701 3519 34759 3525
rect 34701 3516 34713 3519
rect 34664 3488 34713 3516
rect 34664 3476 34670 3488
rect 34701 3485 34713 3488
rect 34747 3485 34759 3519
rect 35529 3519 35587 3525
rect 35529 3516 35541 3519
rect 34701 3479 34759 3485
rect 34808 3488 35541 3516
rect 28718 3448 28724 3460
rect 14516 3420 16988 3448
rect 28000 3420 28724 3448
rect 14516 3408 14522 3420
rect 106 3340 112 3392
rect 164 3380 170 3392
rect 4982 3380 4988 3392
rect 164 3352 4988 3380
rect 164 3340 170 3352
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 16761 3383 16819 3389
rect 16761 3349 16773 3383
rect 16807 3380 16819 3383
rect 17034 3380 17040 3392
rect 16807 3352 17040 3380
rect 16807 3349 16819 3352
rect 16761 3343 16819 3349
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 18874 3340 18880 3392
rect 18932 3340 18938 3392
rect 19797 3383 19855 3389
rect 19797 3349 19809 3383
rect 19843 3380 19855 3383
rect 24394 3380 24400 3392
rect 19843 3352 24400 3380
rect 19843 3349 19855 3352
rect 19797 3343 19855 3349
rect 24394 3340 24400 3352
rect 24452 3340 24458 3392
rect 27614 3340 27620 3392
rect 27672 3340 27678 3392
rect 28000 3389 28028 3420
rect 28718 3408 28724 3420
rect 28776 3408 28782 3460
rect 27985 3383 28043 3389
rect 27985 3349 27997 3383
rect 28031 3349 28043 3383
rect 27985 3343 28043 3349
rect 28258 3340 28264 3392
rect 28316 3340 28322 3392
rect 28626 3340 28632 3392
rect 28684 3340 28690 3392
rect 28902 3340 28908 3392
rect 28960 3340 28966 3392
rect 29181 3383 29239 3389
rect 29181 3349 29193 3383
rect 29227 3380 29239 3383
rect 29546 3380 29552 3392
rect 29227 3352 29552 3380
rect 29227 3349 29239 3352
rect 29181 3343 29239 3349
rect 29546 3340 29552 3352
rect 29604 3340 29610 3392
rect 29733 3383 29791 3389
rect 29733 3349 29745 3383
rect 29779 3380 29791 3383
rect 29914 3380 29920 3392
rect 29779 3352 29920 3380
rect 29779 3349 29791 3352
rect 29733 3343 29791 3349
rect 29914 3340 29920 3352
rect 29972 3340 29978 3392
rect 33410 3340 33416 3392
rect 33468 3380 33474 3392
rect 34808 3380 34836 3488
rect 35529 3485 35541 3488
rect 35575 3485 35587 3519
rect 35529 3479 35587 3485
rect 42797 3519 42855 3525
rect 42797 3485 42809 3519
rect 42843 3516 42855 3519
rect 42889 3519 42947 3525
rect 42889 3516 42901 3519
rect 42843 3488 42901 3516
rect 42843 3485 42855 3488
rect 42797 3479 42855 3485
rect 42889 3485 42901 3488
rect 42935 3485 42947 3519
rect 42889 3479 42947 3485
rect 43901 3519 43959 3525
rect 43901 3485 43913 3519
rect 43947 3485 43959 3519
rect 43901 3479 43959 3485
rect 44269 3519 44327 3525
rect 44269 3485 44281 3519
rect 44315 3516 44327 3519
rect 44726 3516 44732 3528
rect 44315 3488 44732 3516
rect 44315 3485 44327 3488
rect 44269 3479 44327 3485
rect 35066 3408 35072 3460
rect 35124 3448 35130 3460
rect 40586 3448 40592 3460
rect 35124 3420 40592 3448
rect 35124 3408 35130 3420
rect 40586 3408 40592 3420
rect 40644 3408 40650 3460
rect 42242 3408 42248 3460
rect 42300 3448 42306 3460
rect 43916 3448 43944 3479
rect 44726 3476 44732 3488
rect 44784 3476 44790 3528
rect 42300 3420 43944 3448
rect 42300 3408 42306 3420
rect 33468 3352 34836 3380
rect 33468 3340 33474 3352
rect 34882 3340 34888 3392
rect 34940 3380 34946 3392
rect 34977 3383 35035 3389
rect 34977 3380 34989 3383
rect 34940 3352 34989 3380
rect 34940 3340 34946 3352
rect 34977 3349 34989 3352
rect 35023 3349 35035 3383
rect 34977 3343 35035 3349
rect 35713 3383 35771 3389
rect 35713 3349 35725 3383
rect 35759 3380 35771 3383
rect 36262 3380 36268 3392
rect 35759 3352 36268 3380
rect 35759 3349 35771 3352
rect 35713 3343 35771 3349
rect 36262 3340 36268 3352
rect 36320 3340 36326 3392
rect 44082 3340 44088 3392
rect 44140 3340 44146 3392
rect 1104 3290 44896 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 44896 3290
rect 1104 3216 44896 3238
rect 2314 3136 2320 3188
rect 2372 3136 2378 3188
rect 3418 3136 3424 3188
rect 3476 3136 3482 3188
rect 5169 3179 5227 3185
rect 5169 3145 5181 3179
rect 5215 3176 5227 3179
rect 5215 3148 12434 3176
rect 5215 3145 5227 3148
rect 5169 3139 5227 3145
rect 1210 3068 1216 3120
rect 1268 3108 1274 3120
rect 2961 3111 3019 3117
rect 2961 3108 2973 3111
rect 1268 3080 2973 3108
rect 1268 3068 1274 3080
rect 2961 3077 2973 3080
rect 3007 3077 3019 3111
rect 2961 3071 3019 3077
rect 3694 3068 3700 3120
rect 3752 3108 3758 3120
rect 12406 3108 12434 3148
rect 14826 3136 14832 3188
rect 14884 3176 14890 3188
rect 18690 3176 18696 3188
rect 14884 3148 18696 3176
rect 14884 3136 14890 3148
rect 18690 3136 18696 3148
rect 18748 3136 18754 3188
rect 18874 3136 18880 3188
rect 18932 3176 18938 3188
rect 36630 3176 36636 3188
rect 18932 3148 36636 3176
rect 18932 3136 18938 3148
rect 36630 3136 36636 3148
rect 36688 3136 36694 3188
rect 41506 3136 41512 3188
rect 41564 3136 41570 3188
rect 41874 3136 41880 3188
rect 41932 3136 41938 3188
rect 42242 3136 42248 3188
rect 42300 3136 42306 3188
rect 42613 3179 42671 3185
rect 42613 3145 42625 3179
rect 42659 3145 42671 3179
rect 42613 3139 42671 3145
rect 15194 3108 15200 3120
rect 3752 3080 6040 3108
rect 12406 3080 15200 3108
rect 3752 3068 3758 3080
rect 1118 3000 1124 3052
rect 1176 3040 1182 3052
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 1176 3012 2237 3040
rect 1176 3000 1182 3012
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2590 3000 2596 3052
rect 2648 3000 2654 3052
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 2746 3012 3341 3040
rect 382 2932 388 2984
rect 440 2972 446 2984
rect 2746 2972 2774 3012
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 4982 3000 4988 3052
rect 5040 3000 5046 3052
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 6012 3040 6040 3080
rect 15194 3068 15200 3080
rect 15252 3068 15258 3120
rect 15378 3068 15384 3120
rect 15436 3108 15442 3120
rect 15436 3080 20024 3108
rect 15436 3068 15442 3080
rect 19996 3049 20024 3080
rect 25774 3068 25780 3120
rect 25832 3108 25838 3120
rect 28902 3108 28908 3120
rect 25832 3080 28908 3108
rect 25832 3068 25838 3080
rect 28902 3068 28908 3080
rect 28960 3068 28966 3120
rect 41785 3111 41843 3117
rect 41785 3077 41797 3111
rect 41831 3108 41843 3111
rect 42628 3108 42656 3139
rect 43438 3136 43444 3188
rect 43496 3136 43502 3188
rect 44634 3108 44640 3120
rect 41831 3080 42472 3108
rect 42628 3080 44640 3108
rect 41831 3077 41843 3080
rect 41785 3071 41843 3077
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 6012 3012 17417 3040
rect 5261 3003 5319 3009
rect 17405 3009 17417 3012
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3009 19395 3043
rect 19337 3003 19395 3009
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 5276 2972 5304 3003
rect 19352 2972 19380 3003
rect 28626 3000 28632 3052
rect 28684 3040 28690 3052
rect 28813 3043 28871 3049
rect 28813 3040 28825 3043
rect 28684 3012 28825 3040
rect 28684 3000 28690 3012
rect 28813 3009 28825 3012
rect 28859 3009 28871 3043
rect 28813 3003 28871 3009
rect 30285 3043 30343 3049
rect 30285 3009 30297 3043
rect 30331 3040 30343 3043
rect 30377 3043 30435 3049
rect 30377 3040 30389 3043
rect 30331 3012 30389 3040
rect 30331 3009 30343 3012
rect 30285 3003 30343 3009
rect 30377 3009 30389 3012
rect 30423 3009 30435 3043
rect 30377 3003 30435 3009
rect 30653 3043 30711 3049
rect 30653 3009 30665 3043
rect 30699 3009 30711 3043
rect 31113 3043 31171 3049
rect 31113 3040 31125 3043
rect 30653 3003 30711 3009
rect 30852 3012 31125 3040
rect 440 2944 2774 2972
rect 3068 2944 5304 2972
rect 5460 2944 19380 2972
rect 440 2932 446 2944
rect 1026 2864 1032 2916
rect 1084 2904 1090 2916
rect 3068 2904 3096 2944
rect 5460 2913 5488 2944
rect 25038 2932 25044 2984
rect 25096 2972 25102 2984
rect 30668 2972 30696 3003
rect 25096 2944 30696 2972
rect 25096 2932 25102 2944
rect 1084 2876 3096 2904
rect 3145 2907 3203 2913
rect 1084 2864 1090 2876
rect 3145 2873 3157 2907
rect 3191 2904 3203 2907
rect 5445 2907 5503 2913
rect 3191 2876 5396 2904
rect 3191 2873 3203 2876
rect 3145 2867 3203 2873
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2836 2743 2839
rect 4062 2836 4068 2848
rect 2731 2808 4068 2836
rect 2731 2805 2743 2808
rect 2685 2799 2743 2805
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 5368 2836 5396 2876
rect 5445 2873 5457 2907
rect 5491 2873 5503 2907
rect 23198 2904 23204 2916
rect 5445 2867 5503 2873
rect 12406 2876 23204 2904
rect 12406 2836 12434 2876
rect 23198 2864 23204 2876
rect 23256 2864 23262 2916
rect 25222 2864 25228 2916
rect 25280 2904 25286 2916
rect 30852 2913 30880 3012
rect 31113 3009 31125 3012
rect 31159 3009 31171 3043
rect 31113 3003 31171 3009
rect 31478 3000 31484 3052
rect 31536 3000 31542 3052
rect 33686 3000 33692 3052
rect 33744 3000 33750 3052
rect 36262 3000 36268 3052
rect 36320 3000 36326 3052
rect 41690 3000 41696 3052
rect 41748 3000 41754 3052
rect 42444 3049 42472 3080
rect 44634 3068 44640 3080
rect 44692 3068 44698 3120
rect 42061 3043 42119 3049
rect 42061 3040 42073 3043
rect 41800 3012 42073 3040
rect 41601 2975 41659 2981
rect 41601 2941 41613 2975
rect 41647 2972 41659 2975
rect 41800 2972 41828 3012
rect 42061 3009 42073 3012
rect 42107 3009 42119 3043
rect 42061 3003 42119 3009
rect 42429 3043 42487 3049
rect 42429 3009 42441 3043
rect 42475 3009 42487 3043
rect 42429 3003 42487 3009
rect 42705 3043 42763 3049
rect 42705 3009 42717 3043
rect 42751 3009 42763 3043
rect 42705 3003 42763 3009
rect 41647 2944 41828 2972
rect 41969 2975 42027 2981
rect 41647 2941 41659 2944
rect 41601 2935 41659 2941
rect 41969 2941 41981 2975
rect 42015 2972 42027 2975
rect 42720 2972 42748 3003
rect 43162 3000 43168 3052
rect 43220 3000 43226 3052
rect 43254 3000 43260 3052
rect 43312 3000 43318 3052
rect 43346 3000 43352 3052
rect 43404 3040 43410 3052
rect 43901 3043 43959 3049
rect 43901 3040 43913 3043
rect 43404 3012 43913 3040
rect 43404 3000 43410 3012
rect 43901 3009 43913 3012
rect 43947 3009 43959 3043
rect 43901 3003 43959 3009
rect 44269 3043 44327 3049
rect 44269 3009 44281 3043
rect 44315 3009 44327 3043
rect 44269 3003 44327 3009
rect 44284 2972 44312 3003
rect 42015 2944 42748 2972
rect 42904 2944 44312 2972
rect 42015 2941 42027 2944
rect 41969 2935 42027 2941
rect 42904 2913 42932 2944
rect 30193 2907 30251 2913
rect 30193 2904 30205 2907
rect 25280 2876 30205 2904
rect 25280 2864 25286 2876
rect 30193 2873 30205 2876
rect 30239 2873 30251 2907
rect 30193 2867 30251 2873
rect 30837 2907 30895 2913
rect 30837 2873 30849 2907
rect 30883 2873 30895 2907
rect 30837 2867 30895 2873
rect 42889 2907 42947 2913
rect 42889 2873 42901 2907
rect 42935 2873 42947 2907
rect 42889 2867 42947 2873
rect 43162 2864 43168 2916
rect 43220 2904 43226 2916
rect 43717 2907 43775 2913
rect 43717 2904 43729 2907
rect 43220 2876 43729 2904
rect 43220 2864 43226 2876
rect 43717 2873 43729 2876
rect 43763 2873 43775 2907
rect 43717 2867 43775 2873
rect 5368 2808 12434 2836
rect 17589 2839 17647 2845
rect 17589 2805 17601 2839
rect 17635 2836 17647 2839
rect 19150 2836 19156 2848
rect 17635 2808 19156 2836
rect 17635 2805 17647 2808
rect 17589 2799 17647 2805
rect 19150 2796 19156 2808
rect 19208 2796 19214 2848
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 19521 2839 19579 2845
rect 19521 2836 19533 2839
rect 19300 2808 19533 2836
rect 19300 2796 19306 2808
rect 19521 2805 19533 2808
rect 19567 2805 19579 2839
rect 19521 2799 19579 2805
rect 20165 2839 20223 2845
rect 20165 2805 20177 2839
rect 20211 2836 20223 2839
rect 23382 2836 23388 2848
rect 20211 2808 23388 2836
rect 20211 2805 20223 2808
rect 20165 2799 20223 2805
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 28442 2796 28448 2848
rect 28500 2836 28506 2848
rect 28629 2839 28687 2845
rect 28629 2836 28641 2839
rect 28500 2808 28641 2836
rect 28500 2796 28506 2808
rect 28629 2805 28641 2808
rect 28675 2805 28687 2839
rect 28629 2799 28687 2805
rect 30558 2796 30564 2848
rect 30616 2796 30622 2848
rect 31018 2796 31024 2848
rect 31076 2836 31082 2848
rect 31297 2839 31355 2845
rect 31297 2836 31309 2839
rect 31076 2808 31309 2836
rect 31076 2796 31082 2808
rect 31297 2805 31309 2808
rect 31343 2805 31355 2839
rect 31297 2799 31355 2805
rect 31665 2839 31723 2845
rect 31665 2805 31677 2839
rect 31711 2836 31723 2839
rect 32950 2836 32956 2848
rect 31711 2808 32956 2836
rect 31711 2805 31723 2808
rect 31665 2799 31723 2805
rect 32950 2796 32956 2808
rect 33008 2796 33014 2848
rect 33594 2796 33600 2848
rect 33652 2836 33658 2848
rect 33873 2839 33931 2845
rect 33873 2836 33885 2839
rect 33652 2808 33885 2836
rect 33652 2796 33658 2808
rect 33873 2805 33885 2808
rect 33919 2805 33931 2839
rect 33873 2799 33931 2805
rect 36170 2796 36176 2848
rect 36228 2836 36234 2848
rect 36449 2839 36507 2845
rect 36449 2836 36461 2839
rect 36228 2808 36461 2836
rect 36228 2796 36234 2808
rect 36449 2805 36461 2808
rect 36495 2805 36507 2839
rect 36449 2799 36507 2805
rect 42978 2796 42984 2848
rect 43036 2796 43042 2848
rect 43254 2796 43260 2848
rect 43312 2836 43318 2848
rect 43533 2839 43591 2845
rect 43533 2836 43545 2839
rect 43312 2808 43545 2836
rect 43312 2796 43318 2808
rect 43533 2805 43545 2808
rect 43579 2805 43591 2839
rect 43533 2799 43591 2805
rect 44085 2839 44143 2845
rect 44085 2805 44097 2839
rect 44131 2836 44143 2839
rect 44358 2836 44364 2848
rect 44131 2808 44364 2836
rect 44131 2805 44143 2808
rect 44085 2799 44143 2805
rect 44358 2796 44364 2808
rect 44416 2796 44422 2848
rect 44450 2796 44456 2848
rect 44508 2796 44514 2848
rect 1104 2746 44896 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 43950 2746
rect 44002 2694 44014 2746
rect 44066 2694 44078 2746
rect 44130 2694 44142 2746
rect 44194 2694 44206 2746
rect 44258 2694 44896 2746
rect 1104 2672 44896 2694
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11112 2604 22692 2632
rect 11112 2592 11118 2604
rect 10042 2524 10048 2576
rect 10100 2564 10106 2576
rect 16574 2564 16580 2576
rect 10100 2536 16580 2564
rect 10100 2524 10106 2536
rect 16574 2524 16580 2536
rect 16632 2524 16638 2576
rect 19150 2524 19156 2576
rect 19208 2564 19214 2576
rect 19208 2536 21404 2564
rect 19208 2524 19214 2536
rect 7282 2456 7288 2508
rect 7340 2496 7346 2508
rect 7340 2468 19840 2496
rect 7340 2456 7346 2468
rect 19518 2388 19524 2440
rect 19576 2388 19582 2440
rect 19812 2428 19840 2468
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 20036 2468 20392 2496
rect 20036 2456 20042 2468
rect 19877 2431 19935 2437
rect 19877 2428 19889 2431
rect 19812 2400 19889 2428
rect 19877 2397 19889 2400
rect 19923 2397 19935 2431
rect 20257 2431 20315 2437
rect 20257 2428 20269 2431
rect 19877 2391 19935 2397
rect 19996 2400 20269 2428
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 2593 2363 2651 2369
rect 2593 2360 2605 2363
rect 1360 2332 2605 2360
rect 1360 2320 1366 2332
rect 2593 2329 2605 2332
rect 2639 2329 2651 2363
rect 2593 2323 2651 2329
rect 2777 2363 2835 2369
rect 2777 2329 2789 2363
rect 2823 2360 2835 2363
rect 2823 2332 6914 2360
rect 2823 2329 2835 2332
rect 2777 2323 2835 2329
rect 6886 2292 6914 2332
rect 8202 2320 8208 2372
rect 8260 2360 8266 2372
rect 13814 2360 13820 2372
rect 8260 2332 13820 2360
rect 8260 2320 8266 2332
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 15194 2320 15200 2372
rect 15252 2360 15258 2372
rect 19996 2360 20024 2400
rect 20257 2397 20269 2400
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 15252 2332 20024 2360
rect 20364 2360 20392 2468
rect 20530 2456 20536 2508
rect 20588 2496 20594 2508
rect 20588 2468 21036 2496
rect 20588 2456 20594 2468
rect 20622 2388 20628 2440
rect 20680 2388 20686 2440
rect 21008 2437 21036 2468
rect 21376 2437 21404 2536
rect 21450 2524 21456 2576
rect 21508 2564 21514 2576
rect 21508 2536 22600 2564
rect 21508 2524 21514 2536
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 21361 2431 21419 2437
rect 21361 2397 21373 2431
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 21910 2388 21916 2440
rect 21968 2388 21974 2440
rect 22281 2431 22339 2437
rect 22281 2428 22293 2431
rect 22066 2400 22293 2428
rect 22066 2360 22094 2400
rect 22281 2397 22293 2400
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 20364 2332 22094 2360
rect 22572 2360 22600 2536
rect 22664 2437 22692 2604
rect 26786 2592 26792 2644
rect 26844 2632 26850 2644
rect 28074 2632 28080 2644
rect 26844 2604 28080 2632
rect 26844 2592 26850 2604
rect 28074 2592 28080 2604
rect 28132 2592 28138 2644
rect 30006 2592 30012 2644
rect 30064 2632 30070 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 30064 2604 30849 2632
rect 30064 2592 30070 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 33502 2592 33508 2644
rect 33560 2632 33566 2644
rect 33560 2604 35572 2632
rect 33560 2592 33566 2604
rect 22922 2524 22928 2576
rect 22980 2564 22986 2576
rect 23201 2567 23259 2573
rect 23201 2564 23213 2567
rect 22980 2536 23213 2564
rect 22980 2524 22986 2536
rect 23201 2533 23213 2536
rect 23247 2533 23259 2567
rect 23201 2527 23259 2533
rect 24762 2524 24768 2576
rect 24820 2564 24826 2576
rect 25317 2567 25375 2573
rect 25317 2564 25329 2567
rect 24820 2536 25329 2564
rect 24820 2524 24826 2536
rect 25317 2533 25329 2536
rect 25363 2533 25375 2567
rect 25317 2527 25375 2533
rect 26602 2524 26608 2576
rect 26660 2564 26666 2576
rect 27525 2567 27583 2573
rect 27525 2564 27537 2567
rect 26660 2536 27537 2564
rect 26660 2524 26666 2536
rect 27525 2533 27537 2536
rect 27571 2533 27583 2567
rect 27525 2527 27583 2533
rect 27706 2524 27712 2576
rect 27764 2564 27770 2576
rect 28629 2567 28687 2573
rect 28629 2564 28641 2567
rect 27764 2536 28641 2564
rect 27764 2524 27770 2536
rect 28629 2533 28641 2536
rect 28675 2533 28687 2567
rect 28629 2527 28687 2533
rect 28810 2524 28816 2576
rect 28868 2564 28874 2576
rect 29733 2567 29791 2573
rect 29733 2564 29745 2567
rect 28868 2536 29745 2564
rect 28868 2524 28874 2536
rect 29733 2533 29745 2536
rect 29779 2533 29791 2567
rect 29733 2527 29791 2533
rect 30282 2524 30288 2576
rect 30340 2564 30346 2576
rect 31205 2567 31263 2573
rect 31205 2564 31217 2567
rect 30340 2536 31217 2564
rect 30340 2524 30346 2536
rect 31205 2533 31217 2536
rect 31251 2533 31263 2567
rect 31205 2527 31263 2533
rect 31754 2524 31760 2576
rect 31812 2564 31818 2576
rect 32677 2567 32735 2573
rect 32677 2564 32689 2567
rect 31812 2536 32689 2564
rect 31812 2524 31818 2536
rect 32677 2533 32689 2536
rect 32723 2533 32735 2567
rect 32677 2527 32735 2533
rect 32766 2524 32772 2576
rect 32824 2564 32830 2576
rect 33781 2567 33839 2573
rect 33781 2564 33793 2567
rect 32824 2536 33793 2564
rect 32824 2524 32830 2536
rect 33781 2533 33793 2536
rect 33827 2533 33839 2567
rect 33781 2527 33839 2533
rect 34330 2524 34336 2576
rect 34388 2564 34394 2576
rect 35161 2567 35219 2573
rect 35161 2564 35173 2567
rect 34388 2536 35173 2564
rect 34388 2524 34394 2536
rect 35161 2533 35173 2536
rect 35207 2533 35219 2567
rect 35161 2527 35219 2533
rect 22756 2468 23520 2496
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 22756 2360 22784 2468
rect 23014 2388 23020 2440
rect 23072 2388 23078 2440
rect 23382 2388 23388 2440
rect 23440 2388 23446 2440
rect 23492 2428 23520 2468
rect 23566 2456 23572 2508
rect 23624 2496 23630 2508
rect 23624 2468 24808 2496
rect 23624 2456 23630 2468
rect 23753 2431 23811 2437
rect 23753 2428 23765 2431
rect 23492 2400 23765 2428
rect 23753 2397 23765 2400
rect 23799 2397 23811 2431
rect 23753 2391 23811 2397
rect 24394 2388 24400 2440
rect 24452 2388 24458 2440
rect 24780 2437 24808 2468
rect 24946 2456 24952 2508
rect 25004 2496 25010 2508
rect 25004 2468 27016 2496
rect 25004 2456 25010 2468
rect 24765 2431 24823 2437
rect 24765 2397 24777 2431
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 25130 2388 25136 2440
rect 25188 2388 25194 2440
rect 25498 2388 25504 2440
rect 25556 2388 25562 2440
rect 25866 2388 25872 2440
rect 25924 2388 25930 2440
rect 26988 2437 27016 2468
rect 27430 2456 27436 2508
rect 27488 2496 27494 2508
rect 27488 2468 28488 2496
rect 27488 2456 27494 2468
rect 26237 2431 26295 2437
rect 26237 2397 26249 2431
rect 26283 2397 26295 2431
rect 26237 2391 26295 2397
rect 26973 2431 27031 2437
rect 26973 2397 26985 2431
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 22572 2332 22784 2360
rect 15252 2320 15258 2332
rect 24118 2320 24124 2372
rect 24176 2360 24182 2372
rect 26252 2360 26280 2391
rect 27338 2388 27344 2440
rect 27396 2388 27402 2440
rect 27709 2431 27767 2437
rect 27709 2397 27721 2431
rect 27755 2428 27767 2431
rect 27890 2428 27896 2440
rect 27755 2400 27896 2428
rect 27755 2397 27767 2400
rect 27709 2391 27767 2397
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 28074 2388 28080 2440
rect 28132 2388 28138 2440
rect 28460 2437 28488 2468
rect 28534 2456 28540 2508
rect 28592 2496 28598 2508
rect 28592 2468 30052 2496
rect 28592 2456 28598 2468
rect 28445 2431 28503 2437
rect 28445 2397 28457 2431
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 28718 2388 28724 2440
rect 28776 2428 28782 2440
rect 28813 2431 28871 2437
rect 28813 2428 28825 2431
rect 28776 2400 28825 2428
rect 28776 2388 28782 2400
rect 28813 2397 28825 2400
rect 28859 2397 28871 2431
rect 28813 2391 28871 2397
rect 29546 2388 29552 2440
rect 29604 2388 29610 2440
rect 29914 2388 29920 2440
rect 29972 2388 29978 2440
rect 30024 2428 30052 2468
rect 30190 2456 30196 2508
rect 30248 2496 30254 2508
rect 30248 2468 31064 2496
rect 30248 2456 30254 2468
rect 30285 2431 30343 2437
rect 30285 2428 30297 2431
rect 30024 2400 30297 2428
rect 30285 2397 30297 2400
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 30650 2388 30656 2440
rect 30708 2388 30714 2440
rect 31036 2437 31064 2468
rect 32692 2468 33640 2496
rect 32692 2440 32720 2468
rect 31021 2431 31079 2437
rect 31021 2397 31033 2431
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 31389 2431 31447 2437
rect 31389 2397 31401 2431
rect 31435 2397 31447 2431
rect 31389 2391 31447 2397
rect 24176 2332 26280 2360
rect 24176 2320 24182 2332
rect 27430 2320 27436 2372
rect 27488 2360 27494 2372
rect 27488 2332 28304 2360
rect 27488 2320 27494 2332
rect 16574 2292 16580 2304
rect 6886 2264 16580 2292
rect 16574 2252 16580 2264
rect 16632 2252 16638 2304
rect 19610 2252 19616 2304
rect 19668 2292 19674 2304
rect 19705 2295 19763 2301
rect 19705 2292 19717 2295
rect 19668 2264 19717 2292
rect 19668 2252 19674 2264
rect 19705 2261 19717 2264
rect 19751 2261 19763 2295
rect 19705 2255 19763 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 20036 2264 20085 2292
rect 20036 2252 20042 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 20346 2252 20352 2304
rect 20404 2292 20410 2304
rect 20441 2295 20499 2301
rect 20441 2292 20453 2295
rect 20404 2264 20453 2292
rect 20404 2252 20410 2264
rect 20441 2261 20453 2264
rect 20487 2261 20499 2295
rect 20441 2255 20499 2261
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 20809 2295 20867 2301
rect 20809 2292 20821 2295
rect 20772 2264 20821 2292
rect 20772 2252 20778 2264
rect 20809 2261 20821 2264
rect 20855 2261 20867 2295
rect 20809 2255 20867 2261
rect 21177 2295 21235 2301
rect 21177 2261 21189 2295
rect 21223 2292 21235 2295
rect 21358 2292 21364 2304
rect 21223 2264 21364 2292
rect 21223 2261 21235 2264
rect 21177 2255 21235 2261
rect 21358 2252 21364 2264
rect 21416 2252 21422 2304
rect 21450 2252 21456 2304
rect 21508 2292 21514 2304
rect 21545 2295 21603 2301
rect 21545 2292 21557 2295
rect 21508 2264 21557 2292
rect 21508 2252 21514 2264
rect 21545 2261 21557 2264
rect 21591 2261 21603 2295
rect 21545 2255 21603 2261
rect 21818 2252 21824 2304
rect 21876 2292 21882 2304
rect 22097 2295 22155 2301
rect 22097 2292 22109 2295
rect 21876 2264 22109 2292
rect 21876 2252 21882 2264
rect 22097 2261 22109 2264
rect 22143 2261 22155 2295
rect 22097 2255 22155 2261
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 22465 2295 22523 2301
rect 22465 2292 22477 2295
rect 22244 2264 22477 2292
rect 22244 2252 22250 2264
rect 22465 2261 22477 2264
rect 22511 2261 22523 2295
rect 22465 2255 22523 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 22833 2255 22891 2261
rect 23290 2252 23296 2304
rect 23348 2292 23354 2304
rect 23569 2295 23627 2301
rect 23569 2292 23581 2295
rect 23348 2264 23581 2292
rect 23348 2252 23354 2264
rect 23569 2261 23581 2264
rect 23615 2261 23627 2295
rect 23569 2255 23627 2261
rect 23658 2252 23664 2304
rect 23716 2292 23722 2304
rect 23937 2295 23995 2301
rect 23937 2292 23949 2295
rect 23716 2264 23949 2292
rect 23716 2252 23722 2264
rect 23937 2261 23949 2264
rect 23983 2261 23995 2295
rect 23937 2255 23995 2261
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24084 2264 24593 2292
rect 24084 2252 24090 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 24670 2252 24676 2304
rect 24728 2292 24734 2304
rect 24949 2295 25007 2301
rect 24949 2292 24961 2295
rect 24728 2264 24961 2292
rect 24728 2252 24734 2264
rect 24949 2261 24961 2264
rect 24995 2261 25007 2295
rect 24949 2255 25007 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25685 2295 25743 2301
rect 25685 2292 25697 2295
rect 25188 2264 25697 2292
rect 25188 2252 25194 2264
rect 25685 2261 25697 2264
rect 25731 2261 25743 2295
rect 25685 2255 25743 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 26142 2252 26148 2304
rect 26200 2292 26206 2304
rect 26421 2295 26479 2301
rect 26421 2292 26433 2295
rect 26200 2264 26433 2292
rect 26200 2252 26206 2264
rect 26421 2261 26433 2264
rect 26467 2261 26479 2295
rect 26421 2255 26479 2261
rect 26510 2252 26516 2304
rect 26568 2292 26574 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26568 2264 27169 2292
rect 26568 2252 26574 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 27338 2252 27344 2304
rect 27396 2292 27402 2304
rect 28276 2301 28304 2332
rect 29638 2320 29644 2372
rect 29696 2360 29702 2372
rect 29696 2332 30512 2360
rect 29696 2320 29702 2332
rect 27893 2295 27951 2301
rect 27893 2292 27905 2295
rect 27396 2264 27905 2292
rect 27396 2252 27402 2264
rect 27893 2261 27905 2264
rect 27939 2261 27951 2295
rect 27893 2255 27951 2261
rect 28261 2295 28319 2301
rect 28261 2261 28273 2295
rect 28307 2261 28319 2295
rect 28261 2255 28319 2261
rect 28350 2252 28356 2304
rect 28408 2292 28414 2304
rect 28997 2295 29055 2301
rect 28997 2292 29009 2295
rect 28408 2264 29009 2292
rect 28408 2252 28414 2264
rect 28997 2261 29009 2264
rect 29043 2261 29055 2295
rect 28997 2255 29055 2261
rect 29178 2252 29184 2304
rect 29236 2292 29242 2304
rect 30484 2301 30512 2332
rect 30558 2320 30564 2372
rect 30616 2360 30622 2372
rect 31404 2360 31432 2391
rect 32122 2388 32128 2440
rect 32180 2388 32186 2440
rect 32490 2388 32496 2440
rect 32548 2388 32554 2440
rect 32674 2388 32680 2440
rect 32732 2388 32738 2440
rect 32858 2388 32864 2440
rect 32916 2388 32922 2440
rect 32950 2388 32956 2440
rect 33008 2428 33014 2440
rect 33612 2437 33640 2468
rect 33870 2456 33876 2508
rect 33928 2496 33934 2508
rect 33928 2468 35480 2496
rect 33928 2456 33934 2468
rect 33229 2431 33287 2437
rect 33229 2428 33241 2431
rect 33008 2400 33241 2428
rect 33008 2388 33014 2400
rect 33229 2397 33241 2400
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 33597 2431 33655 2437
rect 33597 2397 33609 2431
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 33962 2388 33968 2440
rect 34020 2388 34026 2440
rect 34422 2388 34428 2440
rect 34480 2428 34486 2440
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 34480 2400 34713 2428
rect 34480 2388 34486 2400
rect 34701 2397 34713 2400
rect 34747 2397 34759 2431
rect 34701 2391 34759 2397
rect 35342 2388 35348 2440
rect 35400 2388 35406 2440
rect 35452 2437 35480 2468
rect 35437 2431 35495 2437
rect 35437 2397 35449 2431
rect 35483 2397 35495 2431
rect 35544 2428 35572 2604
rect 35802 2592 35808 2644
rect 35860 2632 35866 2644
rect 36725 2635 36783 2641
rect 36725 2632 36737 2635
rect 35860 2604 36737 2632
rect 35860 2592 35866 2604
rect 36725 2601 36737 2604
rect 36771 2601 36783 2635
rect 36725 2595 36783 2601
rect 37642 2592 37648 2644
rect 37700 2632 37706 2644
rect 38565 2635 38623 2641
rect 38565 2632 38577 2635
rect 37700 2604 38577 2632
rect 37700 2592 37706 2604
rect 38565 2601 38577 2604
rect 38611 2601 38623 2635
rect 38565 2595 38623 2601
rect 42521 2635 42579 2641
rect 42521 2601 42533 2635
rect 42567 2632 42579 2635
rect 44174 2632 44180 2644
rect 42567 2604 44180 2632
rect 42567 2601 42579 2604
rect 42521 2595 42579 2601
rect 44174 2592 44180 2604
rect 44232 2592 44238 2644
rect 44453 2635 44511 2641
rect 44453 2601 44465 2635
rect 44499 2632 44511 2635
rect 44542 2632 44548 2644
rect 44499 2604 44548 2632
rect 44499 2601 44511 2604
rect 44453 2595 44511 2601
rect 44542 2592 44548 2604
rect 44600 2592 44606 2644
rect 35710 2524 35716 2576
rect 35768 2564 35774 2576
rect 36265 2567 36323 2573
rect 36265 2564 36277 2567
rect 35768 2536 36277 2564
rect 35768 2524 35774 2536
rect 36265 2533 36277 2536
rect 36311 2533 36323 2567
rect 36265 2527 36323 2533
rect 36906 2524 36912 2576
rect 36964 2564 36970 2576
rect 37829 2567 37887 2573
rect 37829 2564 37841 2567
rect 36964 2536 37841 2564
rect 36964 2524 36970 2536
rect 37829 2533 37841 2536
rect 37875 2533 37887 2567
rect 37829 2527 37887 2533
rect 38010 2524 38016 2576
rect 38068 2564 38074 2576
rect 38841 2567 38899 2573
rect 38841 2564 38853 2567
rect 38068 2536 38853 2564
rect 38068 2524 38074 2536
rect 38841 2533 38853 2536
rect 38887 2533 38899 2567
rect 38841 2527 38899 2533
rect 43717 2567 43775 2573
rect 43717 2533 43729 2567
rect 43763 2564 43775 2567
rect 44818 2564 44824 2576
rect 43763 2536 44824 2564
rect 43763 2533 43775 2536
rect 43717 2527 43775 2533
rect 44818 2524 44824 2536
rect 44876 2524 44882 2576
rect 35618 2456 35624 2508
rect 35676 2496 35682 2508
rect 37550 2496 37556 2508
rect 35676 2468 36124 2496
rect 35676 2456 35682 2468
rect 35805 2431 35863 2437
rect 35805 2428 35817 2431
rect 35544 2400 35817 2428
rect 35437 2391 35495 2397
rect 35805 2397 35817 2400
rect 35851 2397 35863 2431
rect 35805 2391 35863 2397
rect 30616 2332 31432 2360
rect 30616 2320 30622 2332
rect 32582 2320 32588 2372
rect 32640 2360 32646 2372
rect 32640 2332 33456 2360
rect 32640 2320 32646 2332
rect 30101 2295 30159 2301
rect 30101 2292 30113 2295
rect 29236 2264 30113 2292
rect 29236 2252 29242 2264
rect 30101 2261 30113 2264
rect 30147 2261 30159 2295
rect 30101 2255 30159 2261
rect 30469 2295 30527 2301
rect 30469 2261 30481 2295
rect 30515 2261 30527 2295
rect 30469 2255 30527 2261
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 31573 2295 31631 2301
rect 31573 2292 31585 2295
rect 30984 2264 31585 2292
rect 30984 2252 30990 2264
rect 31573 2261 31585 2264
rect 31619 2261 31631 2295
rect 31573 2255 31631 2261
rect 31662 2252 31668 2304
rect 31720 2292 31726 2304
rect 32309 2295 32367 2301
rect 32309 2292 32321 2295
rect 31720 2264 32321 2292
rect 31720 2252 31726 2264
rect 32309 2261 32321 2264
rect 32355 2261 32367 2295
rect 32309 2255 32367 2261
rect 32398 2252 32404 2304
rect 32456 2292 32462 2304
rect 33428 2301 33456 2332
rect 35066 2320 35072 2372
rect 35124 2360 35130 2372
rect 36096 2360 36124 2468
rect 36464 2468 37556 2496
rect 36464 2437 36492 2468
rect 37550 2456 37556 2468
rect 37608 2456 37614 2508
rect 42978 2496 42984 2508
rect 42720 2468 42984 2496
rect 36449 2431 36507 2437
rect 36449 2397 36461 2431
rect 36495 2397 36507 2431
rect 36449 2391 36507 2397
rect 36538 2388 36544 2440
rect 36596 2388 36602 2440
rect 36630 2388 36636 2440
rect 36688 2428 36694 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36688 2400 37289 2428
rect 36688 2388 36694 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37645 2431 37703 2437
rect 37645 2397 37657 2431
rect 37691 2397 37703 2431
rect 37645 2391 37703 2397
rect 38289 2431 38347 2437
rect 38289 2397 38301 2431
rect 38335 2397 38347 2431
rect 38289 2391 38347 2397
rect 38381 2431 38439 2437
rect 38381 2397 38393 2431
rect 38427 2428 38439 2431
rect 38470 2428 38476 2440
rect 38427 2400 38476 2428
rect 38427 2397 38439 2400
rect 38381 2391 38439 2397
rect 37660 2360 37688 2391
rect 35124 2332 36032 2360
rect 36096 2332 37688 2360
rect 38304 2360 38332 2391
rect 38470 2388 38476 2400
rect 38528 2388 38534 2440
rect 39025 2431 39083 2437
rect 39025 2397 39037 2431
rect 39071 2428 39083 2431
rect 41230 2428 41236 2440
rect 39071 2400 41236 2428
rect 39071 2397 39083 2400
rect 39025 2391 39083 2397
rect 41230 2388 41236 2400
rect 41288 2388 41294 2440
rect 42720 2437 42748 2468
rect 42978 2456 42984 2468
rect 43036 2456 43042 2508
rect 42705 2431 42763 2437
rect 42705 2397 42717 2431
rect 42751 2397 42763 2431
rect 42705 2391 42763 2397
rect 42797 2431 42855 2437
rect 42797 2397 42809 2431
rect 42843 2397 42855 2431
rect 42797 2391 42855 2397
rect 43165 2431 43223 2437
rect 43165 2397 43177 2431
rect 43211 2397 43223 2431
rect 43165 2391 43223 2397
rect 38838 2360 38844 2372
rect 38304 2332 38844 2360
rect 35124 2320 35130 2332
rect 33045 2295 33103 2301
rect 33045 2292 33057 2295
rect 32456 2264 33057 2292
rect 32456 2252 32462 2264
rect 33045 2261 33057 2264
rect 33091 2261 33103 2295
rect 33045 2255 33103 2261
rect 33413 2295 33471 2301
rect 33413 2261 33425 2295
rect 33459 2261 33471 2295
rect 33413 2255 33471 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 34149 2295 34207 2301
rect 34149 2292 34161 2295
rect 33560 2264 34161 2292
rect 33560 2252 33566 2264
rect 34149 2261 34161 2264
rect 34195 2261 34207 2295
rect 34149 2255 34207 2261
rect 34238 2252 34244 2304
rect 34296 2292 34302 2304
rect 34885 2295 34943 2301
rect 34885 2292 34897 2295
rect 34296 2264 34897 2292
rect 34296 2252 34302 2264
rect 34885 2261 34897 2264
rect 34931 2261 34943 2295
rect 34885 2255 34943 2261
rect 34974 2252 34980 2304
rect 35032 2292 35038 2304
rect 36004 2301 36032 2332
rect 38838 2320 38844 2332
rect 38896 2320 38902 2372
rect 41506 2320 41512 2372
rect 41564 2360 41570 2372
rect 42812 2360 42840 2391
rect 43180 2360 43208 2391
rect 43254 2388 43260 2440
rect 43312 2428 43318 2440
rect 43533 2431 43591 2437
rect 43533 2428 43545 2431
rect 43312 2400 43545 2428
rect 43312 2388 43318 2400
rect 43533 2397 43545 2400
rect 43579 2397 43591 2431
rect 43533 2391 43591 2397
rect 43622 2388 43628 2440
rect 43680 2428 43686 2440
rect 43901 2431 43959 2437
rect 43901 2428 43913 2431
rect 43680 2400 43913 2428
rect 43680 2388 43686 2400
rect 43901 2397 43913 2400
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 44269 2431 44327 2437
rect 44269 2397 44281 2431
rect 44315 2428 44327 2431
rect 44634 2428 44640 2440
rect 44315 2400 44640 2428
rect 44315 2397 44327 2400
rect 44269 2391 44327 2397
rect 44634 2388 44640 2400
rect 44692 2388 44698 2440
rect 41564 2332 42840 2360
rect 42904 2332 43208 2360
rect 41564 2320 41570 2332
rect 35621 2295 35679 2301
rect 35621 2292 35633 2295
rect 35032 2264 35633 2292
rect 35032 2252 35038 2264
rect 35621 2261 35633 2264
rect 35667 2261 35679 2295
rect 35621 2255 35679 2261
rect 35989 2295 36047 2301
rect 35989 2261 36001 2295
rect 36035 2261 36047 2295
rect 35989 2255 36047 2261
rect 36814 2252 36820 2304
rect 36872 2292 36878 2304
rect 37461 2295 37519 2301
rect 37461 2292 37473 2295
rect 36872 2264 37473 2292
rect 36872 2252 36878 2264
rect 37461 2261 37473 2264
rect 37507 2261 37519 2295
rect 37461 2255 37519 2261
rect 37550 2252 37556 2304
rect 37608 2292 37614 2304
rect 38105 2295 38163 2301
rect 38105 2292 38117 2295
rect 37608 2264 38117 2292
rect 37608 2252 37614 2264
rect 38105 2261 38117 2264
rect 38151 2261 38163 2295
rect 38105 2255 38163 2261
rect 38194 2252 38200 2304
rect 38252 2292 38258 2304
rect 42904 2292 42932 2332
rect 38252 2264 42932 2292
rect 38252 2252 38258 2264
rect 42978 2252 42984 2304
rect 43036 2252 43042 2304
rect 43346 2252 43352 2304
rect 43404 2252 43410 2304
rect 44082 2252 44088 2304
rect 44140 2252 44146 2304
rect 1104 2202 44896 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 44896 2202
rect 1104 2128 44896 2150
rect 15194 2048 15200 2100
rect 15252 2088 15258 2100
rect 22830 2088 22836 2100
rect 15252 2060 22836 2088
rect 15252 2048 15258 2060
rect 22830 2048 22836 2060
rect 22888 2048 22894 2100
rect 34514 2048 34520 2100
rect 34572 2088 34578 2100
rect 35618 2088 35624 2100
rect 34572 2060 35624 2088
rect 34572 2048 34578 2060
rect 35618 2048 35624 2060
rect 35676 2048 35682 2100
rect 40218 2088 40224 2100
rect 38626 2060 40224 2088
rect 17034 1980 17040 2032
rect 17092 2020 17098 2032
rect 28534 2020 28540 2032
rect 17092 1992 28540 2020
rect 17092 1980 17098 1992
rect 28534 1980 28540 1992
rect 28592 1980 28598 2032
rect 33778 1980 33784 2032
rect 33836 2020 33842 2032
rect 38626 2020 38654 2060
rect 40218 2048 40224 2060
rect 40276 2048 40282 2100
rect 33836 1992 38654 2020
rect 33836 1980 33842 1992
rect 6178 1912 6184 1964
rect 6236 1952 6242 1964
rect 23014 1952 23020 1964
rect 6236 1924 23020 1952
rect 6236 1912 6242 1924
rect 23014 1912 23020 1924
rect 23072 1912 23078 1964
rect 23198 1912 23204 1964
rect 23256 1952 23262 1964
rect 38194 1952 38200 1964
rect 23256 1924 38200 1952
rect 23256 1912 23262 1924
rect 38194 1912 38200 1924
rect 38252 1912 38258 1964
rect 9306 1844 9312 1896
rect 9364 1884 9370 1896
rect 16022 1884 16028 1896
rect 9364 1856 16028 1884
rect 9364 1844 9370 1856
rect 16022 1844 16028 1856
rect 16080 1844 16086 1896
rect 25498 1884 25504 1896
rect 16132 1856 25504 1884
rect 14642 1776 14648 1828
rect 14700 1816 14706 1828
rect 16132 1816 16160 1856
rect 25498 1844 25504 1856
rect 25556 1844 25562 1896
rect 25590 1844 25596 1896
rect 25648 1884 25654 1896
rect 25648 1856 38654 1884
rect 25648 1844 25654 1856
rect 25866 1816 25872 1828
rect 14700 1788 16160 1816
rect 16224 1788 25872 1816
rect 14700 1776 14706 1788
rect 14366 1708 14372 1760
rect 14424 1748 14430 1760
rect 16224 1748 16252 1788
rect 25866 1776 25872 1788
rect 25924 1776 25930 1828
rect 32122 1816 32128 1828
rect 26896 1788 32128 1816
rect 14424 1720 16252 1748
rect 14424 1708 14430 1720
rect 17586 1708 17592 1760
rect 17644 1748 17650 1760
rect 26896 1748 26924 1788
rect 32122 1776 32128 1788
rect 32180 1776 32186 1828
rect 38626 1816 38654 1856
rect 43254 1816 43260 1828
rect 38626 1788 43260 1816
rect 43254 1776 43260 1788
rect 43312 1776 43318 1828
rect 33410 1748 33416 1760
rect 17644 1720 26924 1748
rect 26988 1720 33416 1748
rect 17644 1708 17650 1720
rect 22830 1640 22836 1692
rect 22888 1680 22894 1692
rect 26988 1680 27016 1720
rect 33410 1708 33416 1720
rect 33468 1708 33474 1760
rect 41506 1680 41512 1692
rect 22888 1652 27016 1680
rect 31726 1652 41512 1680
rect 22888 1640 22894 1652
rect 22278 1572 22284 1624
rect 22336 1612 22342 1624
rect 31726 1612 31754 1652
rect 41506 1640 41512 1652
rect 41564 1640 41570 1692
rect 22336 1584 31754 1612
rect 22336 1572 22342 1584
rect 35342 1572 35348 1624
rect 35400 1612 35406 1624
rect 42886 1612 42892 1624
rect 35400 1584 42892 1612
rect 35400 1572 35406 1584
rect 42886 1572 42892 1584
rect 42944 1572 42950 1624
rect 17678 1504 17684 1556
rect 17736 1544 17742 1556
rect 30650 1544 30656 1556
rect 17736 1516 30656 1544
rect 17736 1504 17742 1516
rect 30650 1504 30656 1516
rect 30708 1504 30714 1556
rect 17034 1232 17040 1284
rect 17092 1272 17098 1284
rect 21726 1272 21732 1284
rect 17092 1244 21732 1272
rect 17092 1232 17098 1244
rect 21726 1232 21732 1244
rect 21784 1232 21790 1284
rect 35986 1232 35992 1284
rect 36044 1272 36050 1284
rect 44266 1272 44272 1284
rect 36044 1244 44272 1272
rect 36044 1232 36050 1244
rect 44266 1232 44272 1244
rect 44324 1232 44330 1284
rect 12986 1096 12992 1148
rect 13044 1136 13050 1148
rect 20438 1136 20444 1148
rect 13044 1108 20444 1136
rect 13044 1096 13050 1108
rect 20438 1096 20444 1108
rect 20496 1096 20502 1148
rect 42702 416 42708 468
rect 42760 456 42766 468
rect 45370 456 45376 468
rect 42760 428 45376 456
rect 42760 416 42766 428
rect 45370 416 45376 428
rect 45428 416 45434 468
rect 16298 348 16304 400
rect 16356 388 16362 400
rect 28902 388 28908 400
rect 16356 360 28908 388
rect 16356 348 16362 360
rect 28902 348 28908 360
rect 28960 348 28966 400
rect 15930 280 15936 332
rect 15988 320 15994 332
rect 39482 320 39488 332
rect 15988 292 39488 320
rect 15988 280 15994 292
rect 39482 280 39488 292
rect 39540 280 39546 332
rect 8938 212 8944 264
rect 8996 252 9002 264
rect 25222 252 25228 264
rect 8996 224 25228 252
rect 8996 212 9002 224
rect 25222 212 25228 224
rect 25280 212 25286 264
rect 31110 212 31116 264
rect 31168 252 31174 264
rect 39850 252 39856 264
rect 31168 224 39856 252
rect 31168 212 31174 224
rect 39850 212 39856 224
rect 39908 212 39914 264
rect 13722 144 13728 196
rect 13780 144 13786 196
rect 15562 144 15568 196
rect 15620 184 15626 196
rect 34606 184 34612 196
rect 15620 156 34612 184
rect 15620 144 15626 156
rect 34606 144 34612 156
rect 34664 144 34670 196
rect 13740 116 13768 144
rect 38562 116 38568 128
rect 13740 88 38568 116
rect 38562 76 38568 88
rect 38620 76 38626 128
rect 13446 8 13452 60
rect 13504 48 13510 60
rect 41046 48 41052 60
rect 13504 20 41052 48
rect 13504 8 13510 20
rect 41046 8 41052 20
rect 41104 8 41110 60
<< via1 >>
rect 23296 9324 23348 9376
rect 37464 9324 37516 9376
rect 1308 9256 1360 9308
rect 42524 9256 42576 9308
rect 6644 9188 6696 9240
rect 34428 9188 34480 9240
rect 6552 9120 6604 9172
rect 35440 9120 35492 9172
rect 6736 8984 6788 9036
rect 23204 9052 23256 9104
rect 37648 9052 37700 9104
rect 25412 8984 25464 9036
rect 34336 8984 34388 9036
rect 25136 8916 25188 8968
rect 25320 8916 25372 8968
rect 44640 8916 44692 8968
rect 19064 8848 19116 8900
rect 25412 8848 25464 8900
rect 16948 8780 17000 8832
rect 32864 8848 32916 8900
rect 29828 8780 29880 8832
rect 38568 8780 38620 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 1768 8576 1820 8628
rect 3884 8576 3936 8628
rect 6000 8576 6052 8628
rect 8116 8576 8168 8628
rect 10232 8576 10284 8628
rect 12348 8576 12400 8628
rect 14464 8576 14516 8628
rect 16580 8576 16632 8628
rect 16948 8576 17000 8628
rect 18696 8576 18748 8628
rect 19064 8576 19116 8628
rect 20812 8576 20864 8628
rect 22928 8576 22980 8628
rect 25044 8576 25096 8628
rect 27344 8619 27396 8628
rect 27344 8585 27353 8619
rect 27353 8585 27387 8619
rect 27387 8585 27396 8619
rect 27344 8576 27396 8585
rect 29276 8576 29328 8628
rect 31392 8576 31444 8628
rect 33508 8576 33560 8628
rect 35624 8576 35676 8628
rect 37740 8576 37792 8628
rect 39856 8576 39908 8628
rect 41972 8576 42024 8628
rect 43260 8619 43312 8628
rect 43260 8585 43269 8619
rect 43269 8585 43303 8619
rect 43303 8585 43312 8619
rect 43260 8576 43312 8585
rect 6552 8508 6604 8560
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 9956 8440 10008 8492
rect 11980 8440 12032 8492
rect 13820 8440 13872 8492
rect 16856 8440 16908 8492
rect 44088 8576 44140 8628
rect 23204 8440 23256 8492
rect 23296 8483 23348 8492
rect 23296 8449 23305 8483
rect 23305 8449 23339 8483
rect 23339 8449 23348 8483
rect 23296 8440 23348 8449
rect 44916 8508 44968 8560
rect 29828 8483 29880 8492
rect 29828 8449 29837 8483
rect 29837 8449 29871 8483
rect 29871 8449 29880 8483
rect 29828 8440 29880 8449
rect 32404 8440 32456 8492
rect 34704 8440 34756 8492
rect 35808 8440 35860 8492
rect 38292 8440 38344 8492
rect 39856 8440 39908 8492
rect 39948 8483 40000 8492
rect 39948 8449 39957 8483
rect 39957 8449 39991 8483
rect 39991 8449 40000 8483
rect 39948 8440 40000 8449
rect 40868 8440 40920 8492
rect 42800 8440 42852 8492
rect 43444 8483 43496 8492
rect 43444 8449 43453 8483
rect 43453 8449 43487 8483
rect 43487 8449 43496 8483
rect 43444 8440 43496 8449
rect 43812 8483 43864 8492
rect 43812 8449 43821 8483
rect 43821 8449 43855 8483
rect 43855 8449 43864 8483
rect 43812 8440 43864 8449
rect 36544 8372 36596 8424
rect 43536 8372 43588 8424
rect 40592 8304 40644 8356
rect 44732 8304 44784 8356
rect 39764 8236 39816 8288
rect 43076 8236 43128 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 43950 8134 44002 8186
rect 44014 8134 44066 8186
rect 44078 8134 44130 8186
rect 44142 8134 44194 8186
rect 44206 8134 44258 8186
rect 6736 8032 6788 8084
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 11980 8075 12032 8084
rect 11980 8041 11989 8075
rect 11989 8041 12023 8075
rect 12023 8041 12032 8075
rect 11980 8032 12032 8041
rect 12072 8032 12124 8084
rect 36452 8032 36504 8084
rect 36544 8075 36596 8084
rect 36544 8041 36553 8075
rect 36553 8041 36587 8075
rect 36587 8041 36596 8075
rect 36544 8032 36596 8041
rect 38292 8032 38344 8084
rect 39948 8032 40000 8084
rect 40868 8075 40920 8084
rect 40868 8041 40877 8075
rect 40877 8041 40911 8075
rect 40911 8041 40920 8075
rect 40868 8032 40920 8041
rect 41604 8075 41656 8084
rect 41604 8041 41613 8075
rect 41613 8041 41647 8075
rect 41647 8041 41656 8075
rect 41604 8032 41656 8041
rect 1032 7964 1084 8016
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 1308 7828 1360 7880
rect 39764 7896 39816 7948
rect 756 7760 808 7812
rect 2872 7803 2924 7812
rect 2872 7769 2881 7803
rect 2881 7769 2915 7803
rect 2915 7769 2924 7803
rect 2872 7760 2924 7769
rect 3700 7760 3752 7812
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 12072 7760 12124 7812
rect 3608 7692 3660 7744
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 23572 7871 23624 7880
rect 23572 7837 23581 7871
rect 23581 7837 23615 7871
rect 23615 7837 23624 7871
rect 23572 7828 23624 7837
rect 34796 7828 34848 7880
rect 34888 7871 34940 7880
rect 34888 7837 34897 7871
rect 34897 7837 34931 7871
rect 34931 7837 34940 7871
rect 34888 7828 34940 7837
rect 35992 7871 36044 7880
rect 35992 7837 36001 7871
rect 36001 7837 36035 7871
rect 36035 7837 36044 7871
rect 35992 7828 36044 7837
rect 21916 7760 21968 7812
rect 34428 7760 34480 7812
rect 36636 7760 36688 7812
rect 38384 7760 38436 7812
rect 39488 7871 39540 7880
rect 39488 7837 39497 7871
rect 39497 7837 39531 7871
rect 39531 7837 39540 7871
rect 39488 7828 39540 7837
rect 40040 7871 40092 7880
rect 40040 7837 40049 7871
rect 40049 7837 40083 7871
rect 40083 7837 40092 7871
rect 40040 7828 40092 7837
rect 40684 7871 40736 7880
rect 40684 7837 40693 7871
rect 40693 7837 40727 7871
rect 40727 7837 40736 7871
rect 40684 7828 40736 7837
rect 43444 8032 43496 8084
rect 43720 8075 43772 8084
rect 43720 8041 43729 8075
rect 43729 8041 43763 8075
rect 43763 8041 43772 8075
rect 43720 8032 43772 8041
rect 42800 7964 42852 8016
rect 42064 7871 42116 7880
rect 42064 7837 42073 7871
rect 42073 7837 42107 7871
rect 42107 7837 42116 7871
rect 42064 7828 42116 7837
rect 42524 7871 42576 7880
rect 42524 7837 42533 7871
rect 42533 7837 42567 7871
rect 42567 7837 42576 7871
rect 42524 7828 42576 7837
rect 43352 8007 43404 8016
rect 43352 7973 43361 8007
rect 43361 7973 43395 8007
rect 43395 7973 43404 8007
rect 43352 7964 43404 7973
rect 43076 7896 43128 7948
rect 42984 7828 43036 7880
rect 43168 7871 43220 7880
rect 43168 7837 43177 7871
rect 43177 7837 43211 7871
rect 43211 7837 43220 7871
rect 43168 7828 43220 7837
rect 39672 7760 39724 7812
rect 13820 7692 13872 7744
rect 27896 7692 27948 7744
rect 32404 7735 32456 7744
rect 32404 7701 32413 7735
rect 32413 7701 32447 7735
rect 32447 7701 32456 7735
rect 32404 7692 32456 7701
rect 34704 7735 34756 7744
rect 34704 7701 34713 7735
rect 34713 7701 34747 7735
rect 34747 7701 34756 7735
rect 34704 7692 34756 7701
rect 35808 7735 35860 7744
rect 35808 7701 35817 7735
rect 35817 7701 35851 7735
rect 35851 7701 35860 7735
rect 35808 7692 35860 7701
rect 37556 7692 37608 7744
rect 42064 7692 42116 7744
rect 44548 7828 44600 7880
rect 44272 7692 44324 7744
rect 44456 7735 44508 7744
rect 44456 7701 44465 7735
rect 44465 7701 44499 7735
rect 44499 7701 44508 7735
rect 44456 7692 44508 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 14280 7488 14332 7540
rect 12624 7420 12676 7472
rect 23572 7420 23624 7472
rect 33968 7488 34020 7540
rect 34888 7488 34940 7540
rect 37280 7488 37332 7540
rect 40684 7488 40736 7540
rect 42708 7488 42760 7540
rect 43628 7488 43680 7540
rect 33784 7420 33836 7472
rect 35440 7463 35492 7472
rect 35440 7429 35449 7463
rect 35449 7429 35483 7463
rect 35483 7429 35492 7463
rect 35440 7420 35492 7429
rect 36636 7420 36688 7472
rect 39396 7420 39448 7472
rect 2688 7284 2740 7336
rect 3792 7284 3844 7336
rect 18236 7352 18288 7404
rect 38752 7352 38804 7404
rect 36452 7284 36504 7336
rect 43076 7352 43128 7404
rect 19708 7216 19760 7268
rect 21732 7216 21784 7268
rect 44364 7352 44416 7404
rect 20536 7148 20588 7200
rect 28172 7148 28224 7200
rect 33692 7148 33744 7200
rect 38568 7148 38620 7200
rect 42984 7148 43036 7200
rect 44456 7191 44508 7200
rect 44456 7157 44465 7191
rect 44465 7157 44499 7191
rect 44499 7157 44508 7191
rect 44456 7148 44508 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 43950 7046 44002 7098
rect 44014 7046 44066 7098
rect 44078 7046 44130 7098
rect 44142 7046 44194 7098
rect 44206 7046 44258 7098
rect 40040 6944 40092 6996
rect 44916 6944 44968 6996
rect 1216 6808 1268 6860
rect 1308 6740 1360 6792
rect 17316 6740 17368 6792
rect 5540 6672 5592 6724
rect 6184 6715 6236 6724
rect 6184 6681 6193 6715
rect 6193 6681 6227 6715
rect 6227 6681 6236 6715
rect 6184 6672 6236 6681
rect 41512 6740 41564 6792
rect 42892 6672 42944 6724
rect 4160 6604 4212 6656
rect 18144 6604 18196 6656
rect 28816 6604 28868 6656
rect 33508 6604 33560 6656
rect 39856 6604 39908 6656
rect 44088 6647 44140 6656
rect 44088 6613 44097 6647
rect 44097 6613 44131 6647
rect 44131 6613 44140 6647
rect 44088 6604 44140 6613
rect 44456 6647 44508 6656
rect 44456 6613 44465 6647
rect 44465 6613 44499 6647
rect 44499 6613 44508 6647
rect 44456 6604 44508 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 6184 6400 6236 6452
rect 36820 6400 36872 6452
rect 1124 6332 1176 6384
rect 17960 6332 18012 6384
rect 18512 6332 18564 6384
rect 26976 6332 27028 6384
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 5080 6307 5132 6316
rect 5080 6273 5089 6307
rect 5089 6273 5123 6307
rect 5123 6273 5132 6307
rect 5080 6264 5132 6273
rect 18144 6307 18196 6316
rect 18144 6273 18153 6307
rect 18153 6273 18187 6307
rect 18187 6273 18196 6307
rect 18144 6264 18196 6273
rect 20444 6264 20496 6316
rect 12256 6196 12308 6248
rect 32864 6264 32916 6316
rect 37740 6400 37792 6452
rect 40684 6443 40736 6452
rect 40684 6409 40693 6443
rect 40693 6409 40727 6443
rect 40727 6409 40736 6443
rect 40684 6400 40736 6409
rect 43812 6400 43864 6452
rect 44456 6443 44508 6452
rect 44456 6409 44465 6443
rect 44465 6409 44499 6443
rect 44499 6409 44508 6443
rect 44456 6400 44508 6409
rect 41604 6332 41656 6384
rect 4528 6171 4580 6180
rect 4528 6137 4537 6171
rect 4537 6137 4571 6171
rect 4571 6137 4580 6171
rect 4528 6128 4580 6137
rect 12164 6128 12216 6180
rect 23112 6128 23164 6180
rect 27344 6128 27396 6180
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 20628 6060 20680 6112
rect 26792 6060 26844 6112
rect 34336 6060 34388 6112
rect 42340 6264 42392 6316
rect 42800 6307 42852 6316
rect 42800 6273 42809 6307
rect 42809 6273 42843 6307
rect 42843 6273 42852 6307
rect 42800 6264 42852 6273
rect 37464 6128 37516 6180
rect 42064 6196 42116 6248
rect 41328 6128 41380 6180
rect 40960 6060 41012 6112
rect 41052 6060 41104 6112
rect 43260 6196 43312 6248
rect 44088 6171 44140 6180
rect 44088 6137 44097 6171
rect 44097 6137 44131 6171
rect 44131 6137 44140 6171
rect 44088 6128 44140 6137
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 43950 5958 44002 6010
rect 44014 5958 44066 6010
rect 44078 5958 44130 6010
rect 44142 5958 44194 6010
rect 44206 5958 44258 6010
rect 5172 5856 5224 5908
rect 37188 5856 37240 5908
rect 39672 5856 39724 5908
rect 44640 5856 44692 5908
rect 6092 5788 6144 5840
rect 16488 5788 16540 5840
rect 16672 5788 16724 5840
rect 1032 5652 1084 5704
rect 7104 5652 7156 5704
rect 16488 5559 16540 5568
rect 16488 5525 16497 5559
rect 16497 5525 16531 5559
rect 16531 5525 16540 5559
rect 16488 5516 16540 5525
rect 16856 5584 16908 5636
rect 16672 5516 16724 5568
rect 21456 5516 21508 5568
rect 32772 5788 32824 5840
rect 36820 5788 36872 5840
rect 23112 5720 23164 5772
rect 31116 5720 31168 5772
rect 26976 5695 27028 5704
rect 26976 5661 26985 5695
rect 26985 5661 27019 5695
rect 27019 5661 27028 5695
rect 26976 5652 27028 5661
rect 41512 5720 41564 5772
rect 43168 5763 43220 5772
rect 43168 5729 43177 5763
rect 43177 5729 43211 5763
rect 43211 5729 43220 5763
rect 43168 5720 43220 5729
rect 44456 5831 44508 5840
rect 44456 5797 44465 5831
rect 44465 5797 44499 5831
rect 44499 5797 44508 5831
rect 44456 5788 44508 5797
rect 44824 5720 44876 5772
rect 41420 5584 41472 5636
rect 22376 5516 22428 5568
rect 25136 5516 25188 5568
rect 31484 5559 31536 5568
rect 31484 5525 31493 5559
rect 31493 5525 31527 5559
rect 31527 5525 31536 5559
rect 31484 5516 31536 5525
rect 34428 5516 34480 5568
rect 45192 5516 45244 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 4068 5312 4120 5364
rect 17224 5312 17276 5364
rect 17316 5312 17368 5364
rect 1308 5244 1360 5296
rect 4528 5244 4580 5296
rect 37188 5312 37240 5364
rect 43260 5355 43312 5364
rect 43260 5321 43269 5355
rect 43269 5321 43303 5355
rect 43303 5321 43312 5355
rect 43260 5312 43312 5321
rect 44456 5355 44508 5364
rect 44456 5321 44465 5355
rect 44465 5321 44499 5355
rect 44499 5321 44508 5355
rect 44456 5312 44508 5321
rect 6368 5176 6420 5228
rect 15936 5176 15988 5228
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 3240 5151 3292 5160
rect 3240 5117 3249 5151
rect 3249 5117 3283 5151
rect 3283 5117 3292 5151
rect 3240 5108 3292 5117
rect 16120 5108 16172 5160
rect 19524 5108 19576 5160
rect 16304 5040 16356 5092
rect 6460 4972 6512 5024
rect 16120 4972 16172 5024
rect 16212 5015 16264 5024
rect 16212 4981 16221 5015
rect 16221 4981 16255 5015
rect 16255 4981 16264 5015
rect 16212 4972 16264 4981
rect 16672 4972 16724 5024
rect 22468 5040 22520 5092
rect 44088 5083 44140 5092
rect 44088 5049 44097 5083
rect 44097 5049 44131 5083
rect 44131 5049 44140 5083
rect 44088 5040 44140 5049
rect 23388 4972 23440 5024
rect 33876 4972 33928 5024
rect 44548 4972 44600 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 43950 4870 44002 4922
rect 44014 4870 44066 4922
rect 44078 4870 44130 4922
rect 44142 4870 44194 4922
rect 44206 4870 44258 4922
rect 4528 4768 4580 4820
rect 11888 4768 11940 4820
rect 3424 4700 3476 4752
rect 16212 4768 16264 4820
rect 30288 4768 30340 4820
rect 43536 4768 43588 4820
rect 22284 4700 22336 4752
rect 44364 4700 44416 4752
rect 44456 4743 44508 4752
rect 44456 4709 44465 4743
rect 44465 4709 44499 4743
rect 44499 4709 44508 4743
rect 44456 4700 44508 4709
rect 480 4632 532 4684
rect 664 4564 716 4616
rect 7748 4632 7800 4684
rect 848 4496 900 4548
rect 2320 4539 2372 4548
rect 2320 4505 2329 4539
rect 2329 4505 2363 4539
rect 2363 4505 2372 4539
rect 2320 4496 2372 4505
rect 4896 4496 4948 4548
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 12072 4632 12124 4684
rect 42432 4675 42484 4684
rect 42432 4641 42441 4675
rect 42441 4641 42475 4675
rect 42475 4641 42484 4675
rect 42432 4632 42484 4641
rect 7472 4496 7524 4548
rect 13820 4564 13872 4616
rect 16396 4607 16448 4616
rect 16396 4573 16405 4607
rect 16405 4573 16439 4607
rect 16439 4573 16448 4607
rect 16396 4564 16448 4573
rect 17224 4564 17276 4616
rect 6460 4471 6512 4480
rect 6460 4437 6469 4471
rect 6469 4437 6503 4471
rect 6503 4437 6512 4471
rect 6460 4428 6512 4437
rect 7196 4428 7248 4480
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 15936 4496 15988 4548
rect 17592 4496 17644 4548
rect 38660 4564 38712 4616
rect 25596 4496 25648 4548
rect 43904 4607 43956 4616
rect 43904 4573 43913 4607
rect 43913 4573 43947 4607
rect 43947 4573 43956 4607
rect 43904 4564 43956 4573
rect 44824 4564 44876 4616
rect 45744 4496 45796 4548
rect 17684 4428 17736 4480
rect 24952 4428 25004 4480
rect 38844 4428 38896 4480
rect 41052 4471 41104 4480
rect 41052 4437 41061 4471
rect 41061 4437 41095 4471
rect 41095 4437 41104 4471
rect 41052 4428 41104 4437
rect 41236 4471 41288 4480
rect 41236 4437 41245 4471
rect 41245 4437 41279 4471
rect 41279 4437 41288 4471
rect 41236 4428 41288 4437
rect 44088 4471 44140 4480
rect 44088 4437 44097 4471
rect 44097 4437 44131 4471
rect 44131 4437 44140 4471
rect 44088 4428 44140 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 2412 4224 2464 4276
rect 10876 4224 10928 4276
rect 43904 4224 43956 4276
rect 9680 4156 9732 4208
rect 16396 4156 16448 4208
rect 1860 4088 1912 4140
rect 5264 4088 5316 4140
rect 5632 4020 5684 4072
rect 20904 4088 20956 4140
rect 38568 4131 38620 4140
rect 38568 4097 38577 4131
rect 38577 4097 38611 4131
rect 38611 4097 38620 4131
rect 38568 4088 38620 4097
rect 43444 4088 43496 4140
rect 9956 4020 10008 4072
rect 19616 4020 19668 4072
rect 22376 4020 22428 4072
rect 35072 4020 35124 4072
rect 43260 4020 43312 4072
rect 756 3952 808 4004
rect 44088 3995 44140 4004
rect 44088 3961 44097 3995
rect 44097 3961 44131 3995
rect 44131 3961 44140 3995
rect 44088 3952 44140 3961
rect 44456 3995 44508 4004
rect 44456 3961 44465 3995
rect 44465 3961 44499 3995
rect 44499 3961 44508 3995
rect 44456 3952 44508 3961
rect 6184 3884 6236 3936
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 14648 3884 14700 3936
rect 27436 3884 27488 3936
rect 38476 3884 38528 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 43950 3782 44002 3834
rect 44014 3782 44066 3834
rect 44078 3782 44130 3834
rect 44142 3782 44194 3834
rect 44206 3782 44258 3834
rect 7840 3680 7892 3732
rect 14372 3680 14424 3732
rect 34520 3680 34572 3732
rect 36544 3680 36596 3732
rect 43260 3680 43312 3732
rect 1308 3612 1360 3664
rect 44456 3655 44508 3664
rect 44456 3621 44465 3655
rect 44465 3621 44499 3655
rect 44499 3621 44508 3655
rect 44456 3612 44508 3621
rect 2320 3544 2372 3596
rect 43352 3544 43404 3596
rect 6736 3476 6788 3528
rect 9956 3476 10008 3528
rect 16580 3519 16632 3528
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 14464 3408 14516 3460
rect 18696 3519 18748 3528
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 18696 3476 18748 3485
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 29092 3476 29144 3528
rect 34612 3476 34664 3528
rect 112 3340 164 3392
rect 4988 3340 5040 3392
rect 17040 3340 17092 3392
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 18880 3340 18932 3349
rect 24400 3340 24452 3392
rect 27620 3383 27672 3392
rect 27620 3349 27629 3383
rect 27629 3349 27663 3383
rect 27663 3349 27672 3383
rect 27620 3340 27672 3349
rect 28724 3408 28776 3460
rect 28264 3383 28316 3392
rect 28264 3349 28273 3383
rect 28273 3349 28307 3383
rect 28307 3349 28316 3383
rect 28264 3340 28316 3349
rect 28632 3383 28684 3392
rect 28632 3349 28641 3383
rect 28641 3349 28675 3383
rect 28675 3349 28684 3383
rect 28632 3340 28684 3349
rect 28908 3383 28960 3392
rect 28908 3349 28917 3383
rect 28917 3349 28951 3383
rect 28951 3349 28960 3383
rect 28908 3340 28960 3349
rect 29552 3340 29604 3392
rect 29920 3340 29972 3392
rect 33416 3340 33468 3392
rect 35072 3408 35124 3460
rect 40592 3408 40644 3460
rect 42248 3408 42300 3460
rect 44732 3476 44784 3528
rect 34888 3340 34940 3392
rect 36268 3340 36320 3392
rect 44088 3383 44140 3392
rect 44088 3349 44097 3383
rect 44097 3349 44131 3383
rect 44131 3349 44140 3383
rect 44088 3340 44140 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 1216 3068 1268 3120
rect 3700 3068 3752 3120
rect 14832 3136 14884 3188
rect 18696 3136 18748 3188
rect 18880 3136 18932 3188
rect 36636 3136 36688 3188
rect 41512 3179 41564 3188
rect 41512 3145 41521 3179
rect 41521 3145 41555 3179
rect 41555 3145 41564 3179
rect 41512 3136 41564 3145
rect 41880 3179 41932 3188
rect 41880 3145 41889 3179
rect 41889 3145 41923 3179
rect 41923 3145 41932 3179
rect 41880 3136 41932 3145
rect 42248 3179 42300 3188
rect 42248 3145 42257 3179
rect 42257 3145 42291 3179
rect 42291 3145 42300 3179
rect 42248 3136 42300 3145
rect 1124 3000 1176 3052
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 388 2932 440 2984
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 15200 3068 15252 3120
rect 15384 3068 15436 3120
rect 25780 3068 25832 3120
rect 28908 3068 28960 3120
rect 43444 3179 43496 3188
rect 43444 3145 43453 3179
rect 43453 3145 43487 3179
rect 43487 3145 43496 3179
rect 43444 3136 43496 3145
rect 28632 3000 28684 3052
rect 1032 2864 1084 2916
rect 25044 2932 25096 2984
rect 4068 2796 4120 2848
rect 23204 2864 23256 2916
rect 25228 2864 25280 2916
rect 31484 3043 31536 3052
rect 31484 3009 31493 3043
rect 31493 3009 31527 3043
rect 31527 3009 31536 3043
rect 31484 3000 31536 3009
rect 33692 3043 33744 3052
rect 33692 3009 33701 3043
rect 33701 3009 33735 3043
rect 33735 3009 33744 3043
rect 33692 3000 33744 3009
rect 36268 3043 36320 3052
rect 36268 3009 36277 3043
rect 36277 3009 36311 3043
rect 36311 3009 36320 3043
rect 36268 3000 36320 3009
rect 41696 3043 41748 3052
rect 41696 3009 41705 3043
rect 41705 3009 41739 3043
rect 41739 3009 41748 3043
rect 41696 3000 41748 3009
rect 44640 3068 44692 3120
rect 43168 3043 43220 3052
rect 43168 3009 43177 3043
rect 43177 3009 43211 3043
rect 43211 3009 43220 3043
rect 43168 3000 43220 3009
rect 43260 3043 43312 3052
rect 43260 3009 43269 3043
rect 43269 3009 43303 3043
rect 43303 3009 43312 3043
rect 43260 3000 43312 3009
rect 43352 3000 43404 3052
rect 43168 2864 43220 2916
rect 19156 2796 19208 2848
rect 19248 2796 19300 2848
rect 23388 2796 23440 2848
rect 28448 2796 28500 2848
rect 30564 2839 30616 2848
rect 30564 2805 30573 2839
rect 30573 2805 30607 2839
rect 30607 2805 30616 2839
rect 30564 2796 30616 2805
rect 31024 2796 31076 2848
rect 32956 2796 33008 2848
rect 33600 2796 33652 2848
rect 36176 2796 36228 2848
rect 42984 2839 43036 2848
rect 42984 2805 42993 2839
rect 42993 2805 43027 2839
rect 43027 2805 43036 2839
rect 42984 2796 43036 2805
rect 43260 2796 43312 2848
rect 44364 2796 44416 2848
rect 44456 2839 44508 2848
rect 44456 2805 44465 2839
rect 44465 2805 44499 2839
rect 44499 2805 44508 2839
rect 44456 2796 44508 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 43950 2694 44002 2746
rect 44014 2694 44066 2746
rect 44078 2694 44130 2746
rect 44142 2694 44194 2746
rect 44206 2694 44258 2746
rect 11060 2592 11112 2644
rect 10048 2524 10100 2576
rect 16580 2524 16632 2576
rect 19156 2524 19208 2576
rect 7288 2456 7340 2508
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 19984 2456 20036 2508
rect 1308 2320 1360 2372
rect 8208 2320 8260 2372
rect 13820 2320 13872 2372
rect 15200 2320 15252 2372
rect 20536 2456 20588 2508
rect 20628 2431 20680 2440
rect 20628 2397 20637 2431
rect 20637 2397 20671 2431
rect 20671 2397 20680 2431
rect 20628 2388 20680 2397
rect 21456 2524 21508 2576
rect 21916 2431 21968 2440
rect 21916 2397 21925 2431
rect 21925 2397 21959 2431
rect 21959 2397 21968 2431
rect 21916 2388 21968 2397
rect 26792 2592 26844 2644
rect 28080 2592 28132 2644
rect 30012 2592 30064 2644
rect 33508 2592 33560 2644
rect 22928 2524 22980 2576
rect 24768 2524 24820 2576
rect 26608 2524 26660 2576
rect 27712 2524 27764 2576
rect 28816 2524 28868 2576
rect 30288 2524 30340 2576
rect 31760 2524 31812 2576
rect 32772 2524 32824 2576
rect 34336 2524 34388 2576
rect 23020 2431 23072 2440
rect 23020 2397 23029 2431
rect 23029 2397 23063 2431
rect 23063 2397 23072 2431
rect 23020 2388 23072 2397
rect 23388 2431 23440 2440
rect 23388 2397 23397 2431
rect 23397 2397 23431 2431
rect 23431 2397 23440 2431
rect 23388 2388 23440 2397
rect 23572 2456 23624 2508
rect 24400 2431 24452 2440
rect 24400 2397 24409 2431
rect 24409 2397 24443 2431
rect 24443 2397 24452 2431
rect 24400 2388 24452 2397
rect 24952 2456 25004 2508
rect 25136 2431 25188 2440
rect 25136 2397 25145 2431
rect 25145 2397 25179 2431
rect 25179 2397 25188 2431
rect 25136 2388 25188 2397
rect 25504 2431 25556 2440
rect 25504 2397 25513 2431
rect 25513 2397 25547 2431
rect 25547 2397 25556 2431
rect 25504 2388 25556 2397
rect 25872 2431 25924 2440
rect 25872 2397 25881 2431
rect 25881 2397 25915 2431
rect 25915 2397 25924 2431
rect 25872 2388 25924 2397
rect 27436 2456 27488 2508
rect 24124 2320 24176 2372
rect 27344 2431 27396 2440
rect 27344 2397 27353 2431
rect 27353 2397 27387 2431
rect 27387 2397 27396 2431
rect 27344 2388 27396 2397
rect 27896 2388 27948 2440
rect 28080 2431 28132 2440
rect 28080 2397 28089 2431
rect 28089 2397 28123 2431
rect 28123 2397 28132 2431
rect 28080 2388 28132 2397
rect 28540 2456 28592 2508
rect 28724 2388 28776 2440
rect 29552 2431 29604 2440
rect 29552 2397 29561 2431
rect 29561 2397 29595 2431
rect 29595 2397 29604 2431
rect 29552 2388 29604 2397
rect 29920 2431 29972 2440
rect 29920 2397 29929 2431
rect 29929 2397 29963 2431
rect 29963 2397 29972 2431
rect 29920 2388 29972 2397
rect 30196 2456 30248 2508
rect 30656 2431 30708 2440
rect 30656 2397 30665 2431
rect 30665 2397 30699 2431
rect 30699 2397 30708 2431
rect 30656 2388 30708 2397
rect 27436 2320 27488 2372
rect 16580 2252 16632 2304
rect 19616 2252 19668 2304
rect 19984 2252 20036 2304
rect 20352 2252 20404 2304
rect 20720 2252 20772 2304
rect 21364 2252 21416 2304
rect 21456 2252 21508 2304
rect 21824 2252 21876 2304
rect 22192 2252 22244 2304
rect 22560 2252 22612 2304
rect 23296 2252 23348 2304
rect 23664 2252 23716 2304
rect 24032 2252 24084 2304
rect 24676 2252 24728 2304
rect 25136 2252 25188 2304
rect 25780 2252 25832 2304
rect 26148 2252 26200 2304
rect 26516 2252 26568 2304
rect 27344 2252 27396 2304
rect 29644 2320 29696 2372
rect 28356 2252 28408 2304
rect 29184 2252 29236 2304
rect 30564 2320 30616 2372
rect 32128 2431 32180 2440
rect 32128 2397 32137 2431
rect 32137 2397 32171 2431
rect 32171 2397 32180 2431
rect 32128 2388 32180 2397
rect 32496 2431 32548 2440
rect 32496 2397 32505 2431
rect 32505 2397 32539 2431
rect 32539 2397 32548 2431
rect 32496 2388 32548 2397
rect 32680 2388 32732 2440
rect 32864 2431 32916 2440
rect 32864 2397 32873 2431
rect 32873 2397 32907 2431
rect 32907 2397 32916 2431
rect 32864 2388 32916 2397
rect 32956 2388 33008 2440
rect 33876 2456 33928 2508
rect 33968 2431 34020 2440
rect 33968 2397 33977 2431
rect 33977 2397 34011 2431
rect 34011 2397 34020 2431
rect 33968 2388 34020 2397
rect 34428 2388 34480 2440
rect 35348 2431 35400 2440
rect 35348 2397 35357 2431
rect 35357 2397 35391 2431
rect 35391 2397 35400 2431
rect 35348 2388 35400 2397
rect 35808 2592 35860 2644
rect 37648 2592 37700 2644
rect 44180 2592 44232 2644
rect 44548 2592 44600 2644
rect 35716 2524 35768 2576
rect 36912 2524 36964 2576
rect 38016 2524 38068 2576
rect 44824 2524 44876 2576
rect 35624 2456 35676 2508
rect 32588 2320 32640 2372
rect 30932 2252 30984 2304
rect 31668 2252 31720 2304
rect 32404 2252 32456 2304
rect 35072 2320 35124 2372
rect 37556 2456 37608 2508
rect 36544 2431 36596 2440
rect 36544 2397 36553 2431
rect 36553 2397 36587 2431
rect 36587 2397 36596 2431
rect 36544 2388 36596 2397
rect 36636 2388 36688 2440
rect 38476 2388 38528 2440
rect 41236 2388 41288 2440
rect 42984 2456 43036 2508
rect 33508 2252 33560 2304
rect 34244 2252 34296 2304
rect 34980 2252 35032 2304
rect 38844 2320 38896 2372
rect 41512 2320 41564 2372
rect 43260 2388 43312 2440
rect 43628 2388 43680 2440
rect 44640 2388 44692 2440
rect 36820 2252 36872 2304
rect 37556 2252 37608 2304
rect 38200 2252 38252 2304
rect 42984 2295 43036 2304
rect 42984 2261 42993 2295
rect 42993 2261 43027 2295
rect 43027 2261 43036 2295
rect 42984 2252 43036 2261
rect 43352 2295 43404 2304
rect 43352 2261 43361 2295
rect 43361 2261 43395 2295
rect 43395 2261 43404 2295
rect 43352 2252 43404 2261
rect 44088 2295 44140 2304
rect 44088 2261 44097 2295
rect 44097 2261 44131 2295
rect 44131 2261 44140 2295
rect 44088 2252 44140 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 15200 2048 15252 2100
rect 22836 2048 22888 2100
rect 34520 2048 34572 2100
rect 35624 2048 35676 2100
rect 17040 1980 17092 2032
rect 28540 1980 28592 2032
rect 33784 1980 33836 2032
rect 40224 2048 40276 2100
rect 6184 1912 6236 1964
rect 23020 1912 23072 1964
rect 23204 1912 23256 1964
rect 38200 1912 38252 1964
rect 9312 1844 9364 1896
rect 16028 1844 16080 1896
rect 14648 1776 14700 1828
rect 25504 1844 25556 1896
rect 25596 1844 25648 1896
rect 14372 1708 14424 1760
rect 25872 1776 25924 1828
rect 17592 1708 17644 1760
rect 32128 1776 32180 1828
rect 43260 1776 43312 1828
rect 22836 1640 22888 1692
rect 33416 1708 33468 1760
rect 22284 1572 22336 1624
rect 41512 1640 41564 1692
rect 35348 1572 35400 1624
rect 42892 1572 42944 1624
rect 17684 1504 17736 1556
rect 30656 1504 30708 1556
rect 17040 1232 17092 1284
rect 21732 1232 21784 1284
rect 35992 1232 36044 1284
rect 44272 1232 44324 1284
rect 12992 1096 13044 1148
rect 20444 1096 20496 1148
rect 42708 416 42760 468
rect 45376 416 45428 468
rect 16304 348 16356 400
rect 28908 348 28960 400
rect 15936 280 15988 332
rect 39488 280 39540 332
rect 8944 212 8996 264
rect 25228 212 25280 264
rect 31116 212 31168 264
rect 39856 212 39908 264
rect 13728 144 13780 196
rect 15568 144 15620 196
rect 34612 144 34664 196
rect 38568 76 38620 128
rect 13452 8 13504 60
rect 41052 8 41104 60
<< metal2 >>
rect 1766 11096 1822 11152
rect 3882 11096 3938 11152
rect 5998 11096 6054 11152
rect 8114 11096 8170 11152
rect 10230 11096 10286 11152
rect 12346 11096 12402 11152
rect 14462 11096 14518 11152
rect 16578 11096 16634 11152
rect 18694 11096 18750 11152
rect 20810 11096 20866 11152
rect 22926 11096 22982 11152
rect 25042 11096 25098 11152
rect 27158 11098 27214 11152
rect 27264 11110 27384 11138
rect 27264 11098 27292 11110
rect 27158 11096 27292 11098
rect 1214 9616 1270 9625
rect 1214 9551 1270 9560
rect 754 9344 810 9353
rect 754 9279 810 9288
rect 768 7818 796 9279
rect 1030 8800 1086 8809
rect 1030 8735 1086 8744
rect 1044 8022 1072 8735
rect 1032 8016 1084 8022
rect 1032 7958 1084 7964
rect 1228 7857 1256 9551
rect 1308 9308 1360 9314
rect 1308 9250 1360 9256
rect 1320 8265 1348 9250
rect 1780 8634 1808 11096
rect 2870 9072 2926 9081
rect 2870 9007 2926 9016
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2502 7984 2558 7993
rect 2502 7919 2558 7928
rect 2686 7984 2742 7993
rect 2686 7919 2688 7928
rect 1308 7880 1360 7886
rect 1214 7848 1270 7857
rect 756 7812 808 7818
rect 1308 7822 1360 7828
rect 1214 7783 1270 7792
rect 756 7754 808 7760
rect 1214 7712 1270 7721
rect 1214 7647 1270 7656
rect 1122 7168 1178 7177
rect 1122 7103 1178 7112
rect 1030 6624 1086 6633
rect 1030 6559 1086 6568
rect 662 6080 718 6089
rect 662 6015 718 6024
rect 480 4684 532 4690
rect 480 4626 532 4632
rect 112 3392 164 3398
rect 112 3334 164 3340
rect 124 56 152 3334
rect 388 2984 440 2990
rect 388 2926 440 2932
rect 400 1737 428 2926
rect 386 1728 442 1737
rect 386 1663 442 1672
rect 492 56 520 4626
rect 676 4622 704 6015
rect 1044 5710 1072 6559
rect 1136 6390 1164 7103
rect 1228 6866 1256 7647
rect 1320 7449 1348 7822
rect 1306 7440 1362 7449
rect 1306 7375 1362 7384
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1306 6896 1362 6905
rect 1216 6860 1268 6866
rect 1306 6831 1362 6840
rect 1216 6802 1268 6808
rect 1320 6798 1348 6831
rect 1308 6792 1360 6798
rect 2516 6769 2544 7919
rect 2740 7919 2742 7928
rect 2688 7890 2740 7896
rect 2884 7818 2912 9007
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3896 8634 3924 11096
rect 6012 8634 6040 11096
rect 6644 9240 6696 9246
rect 6644 9182 6696 9188
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6564 8566 6592 9114
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6656 8498 6684 9182
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6748 8090 6776 8978
rect 8128 8634 8156 11096
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 10244 8634 10272 11096
rect 12360 8634 12388 11096
rect 14476 8634 14504 11096
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 16592 8634 16620 11096
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16960 8634 16988 8774
rect 18708 8634 18736 11096
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 19076 8634 19104 8842
rect 20824 8634 20852 11096
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 22940 8634 22968 11096
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23216 8498 23244 9046
rect 23308 8498 23336 9318
rect 25056 8634 25084 11096
rect 27172 11070 27292 11096
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25136 8968 25188 8974
rect 25320 8968 25372 8974
rect 25188 8928 25320 8956
rect 25136 8910 25188 8916
rect 25320 8910 25372 8916
rect 25424 8906 25452 8978
rect 25412 8900 25464 8906
rect 25412 8842 25464 8848
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27356 8634 27384 11110
rect 29274 11096 29330 11152
rect 31390 11096 31446 11152
rect 33506 11096 33562 11152
rect 35622 11096 35678 11152
rect 37738 11096 37794 11152
rect 39854 11096 39910 11152
rect 41970 11096 42026 11152
rect 44086 11096 44142 11152
rect 29288 8634 29316 11096
rect 29828 8832 29880 8838
rect 29828 8774 29880 8780
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 27344 8628 27396 8634
rect 27344 8570 27396 8576
rect 29276 8628 29328 8634
rect 29276 8570 29328 8576
rect 29840 8498 29868 8774
rect 31404 8634 31432 11096
rect 32864 8900 32916 8906
rect 32864 8842 32916 8848
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 23204 8492 23256 8498
rect 23204 8434 23256 8440
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 32404 8492 32456 8498
rect 32404 8434 32456 8440
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 9968 8090 9996 8434
rect 11992 8090 12020 8434
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 1308 6734 1360 6740
rect 2502 6760 2558 6769
rect 2502 6695 2558 6704
rect 1124 6384 1176 6390
rect 1124 6326 1176 6332
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1032 5704 1084 5710
rect 1032 5646 1084 5652
rect 1306 5536 1362 5545
rect 1306 5471 1362 5480
rect 1320 5302 1348 5471
rect 1308 5296 1360 5302
rect 1308 5238 1360 5244
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 664 4616 716 4622
rect 664 4558 716 4564
rect 2318 4584 2374 4593
rect 848 4548 900 4554
rect 2318 4519 2320 4528
rect 848 4490 900 4496
rect 2372 4519 2374 4528
rect 2320 4490 2372 4496
rect 754 4448 810 4457
rect 754 4383 810 4392
rect 768 4010 796 4383
rect 756 4004 808 4010
rect 756 3946 808 3952
rect 860 56 888 4490
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 1306 4176 1362 4185
rect 1306 4111 1362 4120
rect 1860 4140 1912 4146
rect 1320 3670 1348 4111
rect 1860 4082 1912 4088
rect 1398 4040 1454 4049
rect 1398 3975 1454 3984
rect 1308 3664 1360 3670
rect 1412 3641 1440 3975
rect 1308 3606 1360 3612
rect 1398 3632 1454 3641
rect 1398 3567 1454 3576
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 1216 3120 1268 3126
rect 1216 3062 1268 3068
rect 1124 3052 1176 3058
rect 1124 2994 1176 3000
rect 1032 2916 1084 2922
rect 1032 2858 1084 2864
rect 110 0 166 56
rect 478 0 534 56
rect 846 0 902 56
rect 1044 42 1072 2858
rect 1136 2009 1164 2994
rect 1122 2000 1178 2009
rect 1122 1935 1178 1944
rect 1228 1465 1256 3062
rect 1780 2825 1808 3431
rect 1766 2816 1822 2825
rect 1766 2751 1822 2760
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 2281 1348 2314
rect 1306 2272 1362 2281
rect 1306 2207 1362 2216
rect 1872 2122 1900 4082
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2332 3194 2360 3538
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2424 2122 2452 4218
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 1872 2094 1992 2122
rect 1214 1456 1270 1465
rect 1214 1391 1270 1400
rect 1582 640 1638 649
rect 1582 575 1638 584
rect 1136 56 1256 82
rect 1596 56 1624 575
rect 1964 56 1992 2094
rect 2332 2094 2452 2122
rect 2332 56 2360 2094
rect 2608 1193 2636 2994
rect 2594 1184 2650 1193
rect 2594 1119 2650 1128
rect 2700 56 2728 7278
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 3240 5160 3292 5166
rect 3238 5128 3240 5137
rect 3292 5128 3294 5137
rect 3238 5063 3294 5072
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 2870 4040 2926 4049
rect 2870 3975 2926 3984
rect 2884 3369 2912 3975
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3436 3194 3464 4694
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3620 3040 3648 7686
rect 3712 3913 3740 7754
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3698 3904 3754 3913
rect 3698 3839 3754 3848
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 3436 3012 3648 3040
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 3436 218 3464 3012
rect 3712 2938 3740 3062
rect 3344 190 3464 218
rect 3528 2910 3740 2938
rect 3068 56 3188 82
rect 1136 54 1270 56
rect 1136 42 1164 54
rect 1044 14 1164 42
rect 1214 0 1270 54
rect 1582 0 1638 56
rect 1950 0 2006 56
rect 2318 0 2374 56
rect 2686 0 2742 56
rect 3054 54 3188 56
rect 3054 0 3110 54
rect 3160 42 3188 54
rect 3344 42 3372 190
rect 3528 82 3556 2910
rect 3436 56 3556 82
rect 3804 56 3832 7278
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4080 2854 4108 5306
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 4172 56 4200 6598
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4356 5273 4384 6258
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4540 5302 4568 6122
rect 4528 5296 4580 5302
rect 4342 5264 4398 5273
rect 4528 5238 4580 5244
rect 4342 5199 4398 5208
rect 5092 5001 5120 6258
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5914 5212 6054
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5078 4992 5134 5001
rect 5078 4927 5134 4936
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4540 56 4568 4762
rect 5552 4729 5580 6666
rect 6196 6458 6224 6666
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 5538 4720 5594 4729
rect 5538 4655 5594 4664
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4908 56 4936 4490
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 3058 5028 3334
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5276 56 5304 4082
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5644 56 5672 4014
rect 6104 2774 6132 5782
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6012 2746 6132 2774
rect 6012 56 6040 2746
rect 6196 1970 6224 3878
rect 6184 1964 6236 1970
rect 6184 1906 6236 1912
rect 6380 56 6408 5170
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4486 6500 4966
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6748 56 6776 3470
rect 7116 56 7144 5646
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 10152 5273 10180 7822
rect 12084 7818 12112 8026
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12176 6186 12204 7822
rect 13832 7750 13860 8434
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 14292 7546 14320 7822
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 10138 5264 10194 5273
rect 10138 5199 10194 5208
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11900 4706 11928 4762
rect 11900 4690 12112 4706
rect 7748 4684 7800 4690
rect 11900 4684 12124 4690
rect 11900 4678 12072 4684
rect 7748 4626 7800 4632
rect 12072 4626 12124 4632
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7208 1465 7236 4422
rect 7300 2514 7328 4422
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7194 1456 7250 1465
rect 7194 1391 7250 1400
rect 7484 56 7512 4490
rect 7760 2774 7788 4626
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 10888 4282 10916 4558
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 3738 7880 3878
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 7760 2746 7880 2774
rect 7852 56 7880 2746
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 8220 56 8248 2314
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 8574 2000 8630 2009
rect 8574 1935 8630 1944
rect 8588 56 8616 1935
rect 9312 1896 9364 1902
rect 9312 1838 9364 1844
rect 8944 264 8996 270
rect 8944 206 8996 212
rect 8956 56 8984 206
rect 9324 56 9352 1838
rect 9692 56 9720 4150
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9968 3534 9996 4014
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10782 3224 10838 3233
rect 10782 3159 10838 3168
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 10060 56 10088 2518
rect 10414 232 10470 241
rect 10414 167 10470 176
rect 10428 56 10456 167
rect 10796 56 10824 3159
rect 11072 2650 11100 4422
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 12084 2553 12112 4422
rect 12070 2544 12126 2553
rect 12070 2479 12126 2488
rect 11886 1592 11942 1601
rect 11886 1527 11942 1536
rect 11518 504 11574 513
rect 11518 439 11574 448
rect 11150 368 11206 377
rect 11150 303 11206 312
rect 11164 56 11192 303
rect 11532 56 11560 439
rect 11900 56 11928 1527
rect 12268 56 12296 6190
rect 12636 56 12664 7414
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 16488 5840 16540 5846
rect 16672 5840 16724 5846
rect 16540 5788 16672 5794
rect 16488 5782 16724 5788
rect 16500 5766 16712 5782
rect 16868 5642 16896 8434
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 21916 7812 21968 7818
rect 21916 7754 21968 7760
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 16488 5568 16540 5574
rect 16672 5568 16724 5574
rect 16540 5516 16672 5522
rect 16488 5510 16724 5516
rect 16500 5494 16712 5510
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 17328 5370 17356 6734
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 17224 5364 17276 5370
rect 15948 5324 16344 5352
rect 15948 5234 15976 5324
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13832 2378 13860 4558
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 14384 1766 14412 3674
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14372 1760 14424 1766
rect 14372 1702 14424 1708
rect 12992 1148 13044 1154
rect 12992 1090 13044 1096
rect 13004 56 13032 1090
rect 13728 196 13780 202
rect 13728 138 13780 144
rect 13372 66 13492 82
rect 13372 60 13504 66
rect 13372 56 13452 60
rect 3160 14 3372 42
rect 3422 54 3556 56
rect 3422 0 3478 54
rect 3790 0 3846 56
rect 4158 0 4214 56
rect 4526 0 4582 56
rect 4894 0 4950 56
rect 5262 0 5318 56
rect 5630 0 5686 56
rect 5998 0 6054 56
rect 6366 0 6422 56
rect 6734 0 6790 56
rect 7102 0 7158 56
rect 7470 0 7526 56
rect 7838 0 7894 56
rect 8206 0 8262 56
rect 8574 0 8630 56
rect 8942 0 8998 56
rect 9310 0 9366 56
rect 9678 0 9734 56
rect 10046 0 10102 56
rect 10414 0 10470 56
rect 10782 0 10838 56
rect 11150 0 11206 56
rect 11518 0 11574 56
rect 11886 0 11942 56
rect 12254 0 12310 56
rect 12622 0 12678 56
rect 12990 0 13046 56
rect 13358 54 13452 56
rect 13358 0 13414 54
rect 13740 56 13768 138
rect 14094 96 14150 105
rect 13452 2 13504 8
rect 13726 0 13782 56
rect 14476 56 14504 3402
rect 14660 1834 14688 3878
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 14738 3224 14794 3233
rect 15010 3227 15318 3236
rect 14738 3159 14794 3168
rect 14832 3188 14884 3194
rect 14752 2825 14780 3159
rect 14832 3130 14884 3136
rect 14738 2816 14794 2825
rect 14738 2751 14794 2760
rect 14648 1828 14700 1834
rect 14648 1770 14700 1776
rect 14844 56 14872 3130
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15384 3120 15436 3126
rect 15384 3062 15436 3068
rect 15212 2378 15240 3062
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 15200 2100 15252 2106
rect 15200 2042 15252 2048
rect 15212 56 15240 2042
rect 15396 649 15424 3062
rect 15948 2417 15976 4490
rect 15934 2408 15990 2417
rect 15934 2343 15990 2352
rect 16040 1902 16068 5170
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16132 5030 16160 5102
rect 16316 5098 16344 5324
rect 17224 5306 17276 5312
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16224 4826 16252 4966
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16408 4214 16436 4558
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16592 2582 16620 3470
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 16028 1896 16080 1902
rect 16028 1838 16080 1844
rect 16592 1329 16620 2246
rect 16578 1320 16634 1329
rect 16578 1255 16634 1264
rect 15382 640 15438 649
rect 15382 575 15438 584
rect 16304 400 16356 406
rect 16304 342 16356 348
rect 15936 332 15988 338
rect 15936 274 15988 280
rect 15568 196 15620 202
rect 15568 138 15620 144
rect 15580 56 15608 138
rect 15948 56 15976 274
rect 16316 56 16344 342
rect 16684 56 16712 4966
rect 17236 4622 17264 5306
rect 17972 4729 18000 6326
rect 18156 6322 18184 6598
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 17958 4720 18014 4729
rect 17958 4655 18014 4664
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17592 4548 17644 4554
rect 17592 4490 17644 4496
rect 17406 4176 17462 4185
rect 17406 4111 17462 4120
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17052 2038 17080 3334
rect 17040 2032 17092 2038
rect 17040 1974 17092 1980
rect 17040 1284 17092 1290
rect 17040 1226 17092 1232
rect 17052 56 17080 1226
rect 17420 56 17448 4111
rect 17604 1766 17632 4490
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17592 1760 17644 1766
rect 17592 1702 17644 1708
rect 17696 1562 17724 4422
rect 18248 2774 18276 7346
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18156 2746 18276 2774
rect 17774 1728 17830 1737
rect 17774 1663 17830 1672
rect 17684 1556 17736 1562
rect 17684 1498 17736 1504
rect 17788 56 17816 1663
rect 18156 56 18184 2746
rect 18524 56 18552 6326
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18708 3194 18736 3470
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 3194 18920 3334
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18880 3188 18932 3194
rect 18880 3130 18932 3136
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19168 2582 19196 2790
rect 19156 2576 19208 2582
rect 19156 2518 19208 2524
rect 18878 1864 18934 1873
rect 18878 1799 18934 1808
rect 18892 56 18920 1799
rect 19260 56 19288 2790
rect 19536 2446 19564 5102
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 19628 3534 19656 4014
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19720 2530 19748 7210
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 19812 2910 20392 2938
rect 19812 2825 19840 2910
rect 20364 2825 20392 2910
rect 19798 2816 19854 2825
rect 19798 2751 19854 2760
rect 20350 2816 20406 2825
rect 19950 2748 20258 2757
rect 20350 2751 20406 2760
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 19720 2514 20024 2530
rect 19720 2508 20036 2514
rect 19720 2502 19984 2508
rect 19984 2450 20036 2456
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19616 2304 19668 2310
rect 19616 2246 19668 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 19628 56 19656 2246
rect 19996 56 20024 2246
rect 20364 56 20392 2246
rect 20456 1154 20484 6258
rect 20548 2514 20576 7142
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 20640 2446 20668 6054
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 20444 1148 20496 1154
rect 20444 1090 20496 1096
rect 20732 56 20760 2246
rect 20916 1601 20944 4082
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21468 2582 21496 5510
rect 21456 2576 21508 2582
rect 21456 2518 21508 2524
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 20902 1592 20958 1601
rect 20902 1527 20958 1536
rect 21100 56 21220 82
rect 14094 0 14150 40
rect 14462 0 14518 56
rect 14830 0 14886 56
rect 15198 0 15254 56
rect 15566 0 15622 56
rect 15934 0 15990 56
rect 16302 0 16358 56
rect 16670 0 16726 56
rect 17038 0 17094 56
rect 17406 0 17462 56
rect 17774 0 17830 56
rect 18142 0 18198 56
rect 18510 0 18566 56
rect 18878 0 18934 56
rect 19246 0 19302 56
rect 19614 0 19670 56
rect 19982 0 20038 56
rect 20350 0 20406 56
rect 20718 0 20774 56
rect 21086 54 21220 56
rect 21086 0 21142 54
rect 21192 42 21220 54
rect 21376 42 21404 2246
rect 21468 56 21496 2246
rect 21744 1290 21772 7210
rect 21928 2446 21956 7754
rect 23584 7478 23612 7822
rect 32416 7750 32444 8434
rect 27896 7744 27948 7750
rect 27896 7686 27948 7692
rect 32404 7744 32456 7750
rect 32404 7686 32456 7692
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 26976 6384 27028 6390
rect 26976 6326 27028 6332
rect 22466 6216 22522 6225
rect 22466 6151 22522 6160
rect 23112 6180 23164 6186
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22284 4752 22336 4758
rect 22284 4694 22336 4700
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 21824 2304 21876 2310
rect 21824 2246 21876 2252
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 21732 1284 21784 1290
rect 21732 1226 21784 1232
rect 21836 56 21864 2246
rect 22204 56 22232 2246
rect 22296 1630 22324 4694
rect 22388 4078 22416 5510
rect 22480 5098 22508 6151
rect 23112 6122 23164 6128
rect 23124 5778 23152 6122
rect 26792 6112 26844 6118
rect 26792 6054 26844 6060
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 23112 5772 23164 5778
rect 23112 5714 23164 5720
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 22468 5092 22520 5098
rect 22468 5034 22520 5040
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 23400 2938 23428 4966
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 23204 2916 23256 2922
rect 23400 2910 23520 2938
rect 23204 2858 23256 2864
rect 22928 2576 22980 2582
rect 22928 2518 22980 2524
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22284 1624 22336 1630
rect 22284 1566 22336 1572
rect 22572 56 22600 2246
rect 22836 2100 22888 2106
rect 22836 2042 22888 2048
rect 22848 1698 22876 2042
rect 22836 1692 22888 1698
rect 22836 1634 22888 1640
rect 22940 56 22968 2518
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23032 1970 23060 2382
rect 23216 1970 23244 2858
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23400 2446 23428 2790
rect 23492 2774 23520 2910
rect 23492 2746 23612 2774
rect 23584 2514 23612 2746
rect 23572 2508 23624 2514
rect 23572 2450 23624 2456
rect 24412 2446 24440 3334
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23664 2304 23716 2310
rect 23664 2246 23716 2252
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 23020 1964 23072 1970
rect 23020 1906 23072 1912
rect 23204 1964 23256 1970
rect 23204 1906 23256 1912
rect 23308 56 23336 2246
rect 23676 56 23704 2246
rect 24044 56 24072 2246
rect 24136 1465 24164 2314
rect 24676 2304 24728 2310
rect 24676 2246 24728 2252
rect 24122 1456 24178 1465
rect 24122 1391 24178 1400
rect 24412 56 24532 82
rect 21192 14 21404 42
rect 21454 0 21510 56
rect 21822 0 21878 56
rect 22190 0 22246 56
rect 22558 0 22614 56
rect 22926 0 22982 56
rect 23294 0 23350 56
rect 23662 0 23718 56
rect 24030 0 24086 56
rect 24398 54 24532 56
rect 24398 0 24454 54
rect 24504 42 24532 54
rect 24688 42 24716 2246
rect 24780 56 24808 2518
rect 24964 2514 24992 4422
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24952 2508 25004 2514
rect 24952 2450 25004 2456
rect 25056 2009 25084 2926
rect 25148 2446 25176 5510
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25042 2000 25098 2009
rect 25042 1935 25098 1944
rect 25148 56 25176 2246
rect 25240 270 25268 2858
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25516 1902 25544 2382
rect 25608 1902 25636 4490
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25780 3120 25832 3126
rect 25780 3062 25832 3068
rect 25792 2825 25820 3062
rect 25778 2816 25834 2825
rect 25778 2751 25834 2760
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26804 2650 26832 6054
rect 26988 5710 27016 6326
rect 27344 6180 27396 6186
rect 27344 6122 27396 6128
rect 26976 5704 27028 5710
rect 26976 5646 27028 5652
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 26792 2644 26844 2650
rect 26792 2586 26844 2592
rect 26608 2576 26660 2582
rect 26608 2518 26660 2524
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 25504 1896 25556 1902
rect 25504 1838 25556 1844
rect 25596 1896 25648 1902
rect 25596 1838 25648 1844
rect 25228 264 25280 270
rect 25228 206 25280 212
rect 25516 56 25636 82
rect 24504 14 24716 42
rect 24766 0 24822 56
rect 25134 0 25190 56
rect 25502 54 25636 56
rect 25502 0 25558 54
rect 25608 42 25636 54
rect 25792 42 25820 2246
rect 25884 1834 25912 2382
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 25872 1828 25924 1834
rect 25872 1770 25924 1776
rect 25884 56 26004 82
rect 25608 14 25820 42
rect 25870 54 26004 56
rect 25870 0 25926 54
rect 25976 42 26004 54
rect 26160 42 26188 2246
rect 26252 56 26372 82
rect 25976 14 26188 42
rect 26238 54 26372 56
rect 26238 0 26294 54
rect 26344 42 26372 54
rect 26528 42 26556 2246
rect 26620 56 26648 2518
rect 27356 2446 27384 6122
rect 27436 3936 27488 3942
rect 27436 3878 27488 3884
rect 27448 2514 27476 3878
rect 27620 3392 27672 3398
rect 27620 3334 27672 3340
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 27436 2372 27488 2378
rect 27436 2314 27488 2320
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27356 218 27384 2246
rect 27264 190 27384 218
rect 26988 56 27108 82
rect 26344 14 26556 42
rect 26606 0 26662 56
rect 26974 54 27108 56
rect 26974 0 27030 54
rect 27080 42 27108 54
rect 27264 42 27292 190
rect 27448 82 27476 2314
rect 27632 513 27660 3334
rect 27712 2576 27764 2582
rect 27712 2518 27764 2524
rect 27618 504 27674 513
rect 27618 439 27674 448
rect 27356 56 27476 82
rect 27724 56 27752 2518
rect 27908 2446 27936 7686
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28080 2644 28132 2650
rect 28080 2586 28132 2592
rect 28092 2446 28120 2586
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 28184 1737 28212 7142
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 28816 6656 28868 6662
rect 28816 6598 28868 6604
rect 28724 3460 28776 3466
rect 28724 3402 28776 3408
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 28632 3392 28684 3398
rect 28632 3334 28684 3340
rect 28170 1728 28226 1737
rect 28170 1663 28226 1672
rect 28276 377 28304 3334
rect 28644 3058 28672 3334
rect 28632 3052 28684 3058
rect 28632 2994 28684 3000
rect 28448 2848 28500 2854
rect 28448 2790 28500 2796
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 28262 368 28318 377
rect 28262 303 28318 312
rect 28092 56 28212 82
rect 27080 14 27292 42
rect 27342 54 27476 56
rect 27342 0 27398 54
rect 27710 0 27766 56
rect 28078 54 28212 56
rect 28078 0 28134 54
rect 28184 42 28212 54
rect 28368 42 28396 2246
rect 28460 56 28488 2790
rect 28540 2508 28592 2514
rect 28540 2450 28592 2456
rect 28552 2038 28580 2450
rect 28736 2446 28764 3402
rect 28828 2774 28856 6598
rect 32876 6322 32904 8842
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 33520 8634 33548 11096
rect 34428 9240 34480 9246
rect 34428 9182 34480 9188
rect 34336 9036 34388 9042
rect 34336 8978 34388 8984
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33968 7540 34020 7546
rect 33968 7482 34020 7488
rect 33784 7472 33836 7478
rect 33784 7414 33836 7420
rect 33692 7200 33744 7206
rect 33692 7142 33744 7148
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 32864 6316 32916 6322
rect 32864 6258 32916 6264
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32772 5840 32824 5846
rect 32772 5782 32824 5788
rect 31116 5772 31168 5778
rect 31116 5714 31168 5720
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 3126 28948 3334
rect 28908 3120 28960 3126
rect 28908 3062 28960 3068
rect 28828 2746 28948 2774
rect 28816 2576 28868 2582
rect 28816 2518 28868 2524
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 28540 2032 28592 2038
rect 28540 1974 28592 1980
rect 28828 56 28856 2518
rect 28920 406 28948 2746
rect 28908 400 28960 406
rect 28908 342 28960 348
rect 29104 241 29132 3470
rect 29552 3392 29604 3398
rect 29552 3334 29604 3340
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 29564 2446 29592 3334
rect 29932 2446 29960 3334
rect 30300 2666 30328 4762
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 30012 2644 30064 2650
rect 30012 2586 30064 2592
rect 30208 2638 30328 2666
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29920 2440 29972 2446
rect 29920 2382 29972 2388
rect 29644 2372 29696 2378
rect 29644 2314 29696 2320
rect 29184 2304 29236 2310
rect 29184 2246 29236 2252
rect 29090 232 29146 241
rect 29090 167 29146 176
rect 29196 56 29224 2246
rect 29656 1170 29684 2314
rect 30024 1170 30052 2586
rect 30208 2514 30236 2638
rect 30288 2576 30340 2582
rect 30288 2518 30340 2524
rect 30196 2508 30248 2514
rect 30196 2450 30248 2456
rect 29564 1142 29684 1170
rect 29932 1142 30052 1170
rect 29564 56 29592 1142
rect 29932 56 29960 1142
rect 30300 56 30328 2518
rect 30576 2378 30604 2790
rect 30656 2440 30708 2446
rect 30656 2382 30708 2388
rect 30564 2372 30616 2378
rect 30564 2314 30616 2320
rect 30668 1562 30696 2382
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 30656 1556 30708 1562
rect 30656 1498 30708 1504
rect 30668 56 30788 82
rect 28184 14 28396 42
rect 28446 0 28502 56
rect 28814 0 28870 56
rect 29182 0 29238 56
rect 29550 0 29606 56
rect 29918 0 29974 56
rect 30286 0 30342 56
rect 30654 54 30788 56
rect 30654 0 30710 54
rect 30760 42 30788 54
rect 30944 42 30972 2246
rect 31036 56 31064 2790
rect 31128 270 31156 5714
rect 31484 5568 31536 5574
rect 31484 5510 31536 5516
rect 31496 4185 31524 5510
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31482 4176 31538 4185
rect 31482 4111 31538 4120
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31484 3052 31536 3058
rect 31484 2994 31536 3000
rect 31496 1873 31524 2994
rect 32784 2774 32812 5782
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 33416 3392 33468 3398
rect 33416 3334 33468 3340
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32692 2746 32812 2774
rect 31760 2576 31812 2582
rect 31760 2518 31812 2524
rect 31668 2304 31720 2310
rect 31668 2246 31720 2252
rect 31482 1864 31538 1873
rect 31482 1799 31538 1808
rect 31116 264 31168 270
rect 31116 206 31168 212
rect 31404 56 31524 82
rect 30760 14 30972 42
rect 31022 0 31078 56
rect 31390 54 31524 56
rect 31390 0 31446 54
rect 31496 42 31524 54
rect 31680 42 31708 2246
rect 31772 56 31800 2518
rect 32692 2446 32720 2746
rect 32772 2576 32824 2582
rect 32772 2518 32824 2524
rect 32862 2544 32918 2553
rect 32128 2440 32180 2446
rect 32496 2440 32548 2446
rect 32128 2382 32180 2388
rect 32494 2408 32496 2417
rect 32680 2440 32732 2446
rect 32548 2408 32550 2417
rect 32140 1834 32168 2382
rect 32680 2382 32732 2388
rect 32494 2343 32550 2352
rect 32588 2372 32640 2378
rect 32588 2314 32640 2320
rect 32404 2304 32456 2310
rect 32404 2246 32456 2252
rect 32128 1828 32180 1834
rect 32128 1770 32180 1776
rect 32140 56 32260 82
rect 31496 14 31708 42
rect 31758 0 31814 56
rect 32126 54 32260 56
rect 32126 0 32182 54
rect 32232 42 32260 54
rect 32416 42 32444 2246
rect 32600 1170 32628 2314
rect 32508 1142 32628 1170
rect 32784 1170 32812 2518
rect 32862 2479 32918 2488
rect 32876 2446 32904 2479
rect 32968 2446 32996 2790
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 33428 1766 33456 3334
rect 33520 2650 33548 6598
rect 33704 3058 33732 7142
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 33600 2848 33652 2854
rect 33600 2790 33652 2796
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 33416 1760 33468 1766
rect 33416 1702 33468 1708
rect 32784 1142 32904 1170
rect 32508 56 32536 1142
rect 32876 56 32904 1142
rect 33244 56 33364 82
rect 32232 14 32444 42
rect 32494 0 32550 56
rect 32862 0 32918 56
rect 33230 54 33364 56
rect 33230 0 33286 54
rect 33336 42 33364 54
rect 33520 42 33548 2246
rect 33612 56 33640 2790
rect 33796 2038 33824 7414
rect 33876 5024 33928 5030
rect 33876 4966 33928 4972
rect 33888 2514 33916 4966
rect 33876 2508 33928 2514
rect 33876 2450 33928 2456
rect 33980 2446 34008 7482
rect 34348 6118 34376 8978
rect 34440 7818 34468 9182
rect 35440 9172 35492 9178
rect 35440 9114 35492 9120
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 34428 7812 34480 7818
rect 34428 7754 34480 7760
rect 34716 7750 34744 8434
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34888 7880 34940 7886
rect 34888 7822 34940 7828
rect 34704 7744 34756 7750
rect 34704 7686 34756 7692
rect 34336 6112 34388 6118
rect 34336 6054 34388 6060
rect 34428 5568 34480 5574
rect 34428 5510 34480 5516
rect 34336 2576 34388 2582
rect 34336 2518 34388 2524
rect 33968 2440 34020 2446
rect 33968 2382 34020 2388
rect 34244 2304 34296 2310
rect 34244 2246 34296 2252
rect 33784 2032 33836 2038
rect 33784 1974 33836 1980
rect 33980 56 34100 82
rect 33336 14 33548 42
rect 33598 0 33654 56
rect 33966 54 34100 56
rect 33966 0 34022 54
rect 34072 42 34100 54
rect 34256 42 34284 2246
rect 34348 56 34376 2518
rect 34440 2446 34468 5510
rect 34808 5273 34836 7822
rect 34900 7546 34928 7822
rect 34888 7540 34940 7546
rect 34888 7482 34940 7488
rect 35452 7478 35480 9114
rect 35636 8634 35664 11096
rect 37464 9376 37516 9382
rect 37464 9318 37516 9324
rect 35624 8628 35676 8634
rect 35624 8570 35676 8576
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35820 7750 35848 8434
rect 36544 8424 36596 8430
rect 36544 8366 36596 8372
rect 36556 8090 36584 8366
rect 36452 8084 36504 8090
rect 36452 8026 36504 8032
rect 36544 8084 36596 8090
rect 36544 8026 36596 8032
rect 35992 7880 36044 7886
rect 35992 7822 36044 7828
rect 35808 7744 35860 7750
rect 35808 7686 35860 7692
rect 35440 7472 35492 7478
rect 35440 7414 35492 7420
rect 34794 5264 34850 5273
rect 34794 5199 34850 5208
rect 35072 4072 35124 4078
rect 35072 4014 35124 4020
rect 34520 3732 34572 3738
rect 34520 3674 34572 3680
rect 34428 2440 34480 2446
rect 34428 2382 34480 2388
rect 34532 2106 34560 3674
rect 34612 3528 34664 3534
rect 34612 3470 34664 3476
rect 34624 3380 34652 3470
rect 35084 3466 35112 4014
rect 35072 3460 35124 3466
rect 35072 3402 35124 3408
rect 34888 3392 34940 3398
rect 34624 3352 34888 3380
rect 34520 2100 34572 2106
rect 34520 2042 34572 2048
rect 34624 202 34652 3352
rect 34888 3334 34940 3340
rect 35808 2644 35860 2650
rect 35808 2586 35860 2592
rect 35716 2576 35768 2582
rect 35716 2518 35768 2524
rect 35624 2508 35676 2514
rect 35624 2450 35676 2456
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 35072 2372 35124 2378
rect 35072 2314 35124 2320
rect 34980 2304 35032 2310
rect 34980 2246 35032 2252
rect 34612 196 34664 202
rect 34612 138 34664 144
rect 34716 56 34836 82
rect 34072 14 34284 42
rect 34334 0 34390 56
rect 34702 54 34836 56
rect 34702 0 34758 54
rect 34808 42 34836 54
rect 34992 42 35020 2246
rect 35084 56 35112 2314
rect 35360 1630 35388 2382
rect 35636 2106 35664 2450
rect 35624 2100 35676 2106
rect 35624 2042 35676 2048
rect 35348 1624 35400 1630
rect 35348 1566 35400 1572
rect 35452 56 35572 82
rect 34808 14 35020 42
rect 35070 0 35126 56
rect 35438 54 35572 56
rect 35438 0 35494 54
rect 35544 42 35572 54
rect 35728 42 35756 2518
rect 35820 56 35848 2586
rect 36004 1290 36032 7822
rect 36464 7342 36492 8026
rect 36636 7812 36688 7818
rect 36636 7754 36688 7760
rect 36648 7478 36676 7754
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 36636 7472 36688 7478
rect 36636 7414 36688 7420
rect 36452 7336 36504 7342
rect 36452 7278 36504 7284
rect 36820 6452 36872 6458
rect 36820 6394 36872 6400
rect 36832 5846 36860 6394
rect 37188 5908 37240 5914
rect 37188 5850 37240 5856
rect 36820 5840 36872 5846
rect 36820 5782 36872 5788
rect 37200 5370 37228 5850
rect 37292 5681 37320 7482
rect 37476 6186 37504 9318
rect 37648 9104 37700 9110
rect 37648 9046 37700 9052
rect 37556 7744 37608 7750
rect 37556 7686 37608 7692
rect 37464 6180 37516 6186
rect 37464 6122 37516 6128
rect 37278 5672 37334 5681
rect 37278 5607 37334 5616
rect 37188 5364 37240 5370
rect 37188 5306 37240 5312
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 36268 3392 36320 3398
rect 36268 3334 36320 3340
rect 36280 3058 36308 3334
rect 36268 3052 36320 3058
rect 36268 2994 36320 3000
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 35992 1284 36044 1290
rect 35992 1226 36044 1232
rect 36188 56 36216 2790
rect 36556 2446 36584 3674
rect 36636 3188 36688 3194
rect 36636 3130 36688 3136
rect 36648 2446 36676 3130
rect 36912 2576 36964 2582
rect 36912 2518 36964 2524
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36636 2440 36688 2446
rect 36636 2382 36688 2388
rect 36820 2304 36872 2310
rect 36820 2246 36872 2252
rect 36556 56 36676 82
rect 35544 14 35756 42
rect 35806 0 35862 56
rect 36174 0 36230 56
rect 36542 54 36676 56
rect 36542 0 36598 54
rect 36648 42 36676 54
rect 36832 42 36860 2246
rect 36924 56 36952 2518
rect 37568 2514 37596 7686
rect 37660 6914 37688 9046
rect 37752 8634 37780 11096
rect 38568 8832 38620 8838
rect 38568 8774 38620 8780
rect 37740 8628 37792 8634
rect 37740 8570 37792 8576
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 38304 8090 38332 8434
rect 38292 8084 38344 8090
rect 38292 8026 38344 8032
rect 38384 7812 38436 7818
rect 38384 7754 38436 7760
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 37660 6886 37780 6914
rect 37752 6458 37780 6886
rect 37740 6452 37792 6458
rect 37740 6394 37792 6400
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 37648 2644 37700 2650
rect 37648 2586 37700 2592
rect 37556 2508 37608 2514
rect 37556 2450 37608 2456
rect 37556 2304 37608 2310
rect 37556 2246 37608 2252
rect 37292 56 37412 82
rect 36648 14 36860 42
rect 36910 0 36966 56
rect 37278 54 37412 56
rect 37278 0 37334 54
rect 37384 42 37412 54
rect 37568 42 37596 2246
rect 37660 56 37688 2586
rect 38016 2576 38068 2582
rect 38016 2518 38068 2524
rect 38028 56 38056 2518
rect 38200 2304 38252 2310
rect 38200 2246 38252 2252
rect 38212 1970 38240 2246
rect 38200 1964 38252 1970
rect 38200 1906 38252 1912
rect 38396 56 38424 7754
rect 38580 7206 38608 8774
rect 39010 8732 39318 8741
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 39868 8634 39896 11096
rect 41984 8634 42012 11096
rect 42982 9616 43038 9625
rect 42982 9551 43038 9560
rect 42524 9308 42576 9314
rect 42524 9250 42576 9256
rect 39856 8628 39908 8634
rect 39856 8570 39908 8576
rect 41972 8628 42024 8634
rect 41972 8570 42024 8576
rect 41602 8528 41658 8537
rect 39856 8492 39908 8498
rect 39856 8434 39908 8440
rect 39948 8492 40000 8498
rect 39948 8434 40000 8440
rect 40868 8492 40920 8498
rect 41602 8463 41658 8472
rect 40868 8434 40920 8440
rect 39764 8288 39816 8294
rect 39764 8230 39816 8236
rect 39776 7954 39804 8230
rect 39764 7948 39816 7954
rect 39764 7890 39816 7896
rect 39488 7880 39540 7886
rect 39488 7822 39540 7828
rect 39010 7644 39318 7653
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39396 7472 39448 7478
rect 39396 7414 39448 7420
rect 38752 7404 38804 7410
rect 38752 7346 38804 7352
rect 38568 7200 38620 7206
rect 38568 7142 38620 7148
rect 38660 4616 38712 4622
rect 38660 4558 38712 4564
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 38476 3936 38528 3942
rect 38476 3878 38528 3884
rect 38488 2446 38516 3878
rect 38476 2440 38528 2446
rect 38476 2382 38528 2388
rect 38580 134 38608 4082
rect 38568 128 38620 134
rect 38672 105 38700 4558
rect 38568 70 38620 76
rect 38658 96 38714 105
rect 37384 14 37596 42
rect 37646 0 37702 56
rect 38014 0 38070 56
rect 38382 0 38438 56
rect 38764 56 38792 7346
rect 39010 6556 39318 6565
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 38844 4480 38896 4486
rect 38844 4422 38896 4428
rect 38856 2378 38884 4422
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 38844 2372 38896 2378
rect 38844 2314 38896 2320
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 39132 56 39252 82
rect 38658 31 38714 40
rect 38750 0 38806 56
rect 39118 54 39252 56
rect 39118 0 39174 54
rect 39224 42 39252 54
rect 39408 42 39436 7414
rect 39500 338 39528 7822
rect 39672 7812 39724 7818
rect 39672 7754 39724 7760
rect 39684 5914 39712 7754
rect 39868 6662 39896 8434
rect 39960 8090 39988 8434
rect 40592 8356 40644 8362
rect 40592 8298 40644 8304
rect 39948 8084 40000 8090
rect 39948 8026 40000 8032
rect 40040 7880 40092 7886
rect 40040 7822 40092 7828
rect 40052 7002 40080 7822
rect 40040 6996 40092 7002
rect 40040 6938 40092 6944
rect 40604 6914 40632 8298
rect 40880 8090 40908 8434
rect 41616 8090 41644 8463
rect 40868 8084 40920 8090
rect 40868 8026 40920 8032
rect 41604 8084 41656 8090
rect 41604 8026 41656 8032
rect 42536 7886 42564 9250
rect 42800 8492 42852 8498
rect 42800 8434 42852 8440
rect 42812 8022 42840 8434
rect 42800 8016 42852 8022
rect 42800 7958 42852 7964
rect 42996 7886 43024 9551
rect 43350 9344 43406 9353
rect 43350 9279 43406 9288
rect 43260 8628 43312 8634
rect 43260 8570 43312 8576
rect 43272 8537 43300 8570
rect 43258 8528 43314 8537
rect 43258 8463 43314 8472
rect 43076 8288 43128 8294
rect 43076 8230 43128 8236
rect 43088 7954 43116 8230
rect 43364 8022 43392 9279
rect 43626 9072 43682 9081
rect 43626 9007 43682 9016
rect 43444 8492 43496 8498
rect 43444 8434 43496 8440
rect 43456 8090 43484 8434
rect 43536 8424 43588 8430
rect 43536 8366 43588 8372
rect 43444 8084 43496 8090
rect 43444 8026 43496 8032
rect 43352 8016 43404 8022
rect 43166 7984 43222 7993
rect 43076 7948 43128 7954
rect 43352 7958 43404 7964
rect 43166 7919 43222 7928
rect 43076 7890 43128 7896
rect 43180 7886 43208 7919
rect 40684 7880 40736 7886
rect 42064 7880 42116 7886
rect 40684 7822 40736 7828
rect 42062 7848 42064 7857
rect 42524 7880 42576 7886
rect 42116 7848 42118 7857
rect 40696 7546 40724 7822
rect 42524 7822 42576 7828
rect 42984 7880 43036 7886
rect 42984 7822 43036 7828
rect 43168 7880 43220 7886
rect 43168 7822 43220 7828
rect 42062 7783 42118 7792
rect 42076 7750 42104 7783
rect 42064 7744 42116 7750
rect 42064 7686 42116 7692
rect 40684 7540 40736 7546
rect 40684 7482 40736 7488
rect 42708 7540 42760 7546
rect 42708 7482 42760 7488
rect 40604 6886 40724 6914
rect 39856 6656 39908 6662
rect 39856 6598 39908 6604
rect 40696 6458 40724 6886
rect 41512 6792 41564 6798
rect 41512 6734 41564 6740
rect 40684 6452 40736 6458
rect 40684 6394 40736 6400
rect 41328 6180 41380 6186
rect 41328 6122 41380 6128
rect 40960 6112 41012 6118
rect 40960 6054 41012 6060
rect 41052 6112 41104 6118
rect 41052 6054 41104 6060
rect 39672 5908 39724 5914
rect 39672 5850 39724 5856
rect 40592 3460 40644 3466
rect 40592 3402 40644 3408
rect 40224 2100 40276 2106
rect 40224 2042 40276 2048
rect 39488 332 39540 338
rect 39488 274 39540 280
rect 39856 264 39908 270
rect 39486 232 39542 241
rect 39856 206 39908 212
rect 39486 167 39542 176
rect 39500 56 39528 167
rect 39868 56 39896 206
rect 40236 56 40264 2042
rect 40604 56 40632 3402
rect 40972 56 41000 6054
rect 41064 4593 41092 6054
rect 41050 4584 41106 4593
rect 41050 4519 41106 4528
rect 41052 4480 41104 4486
rect 41052 4422 41104 4428
rect 41236 4480 41288 4486
rect 41236 4422 41288 4428
rect 41064 66 41092 4422
rect 41248 2446 41276 4422
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 41052 60 41104 66
rect 39224 14 39436 42
rect 39486 0 39542 56
rect 39854 0 39910 56
rect 40222 0 40278 56
rect 40590 0 40646 56
rect 40958 0 41014 56
rect 41340 56 41368 6122
rect 41524 5778 41552 6734
rect 41604 6384 41656 6390
rect 41604 6326 41656 6332
rect 41512 5772 41564 5778
rect 41512 5714 41564 5720
rect 41420 5636 41472 5642
rect 41420 5578 41472 5584
rect 41432 5137 41460 5578
rect 41418 5128 41474 5137
rect 41418 5063 41474 5072
rect 41510 4040 41566 4049
rect 41510 3975 41566 3984
rect 41524 3194 41552 3975
rect 41512 3188 41564 3194
rect 41512 3130 41564 3136
rect 41616 2938 41644 6326
rect 42340 6316 42392 6322
rect 42340 6258 42392 6264
rect 42064 6248 42116 6254
rect 42064 6190 42116 6196
rect 41878 3496 41934 3505
rect 41878 3431 41934 3440
rect 41892 3194 41920 3431
rect 41880 3188 41932 3194
rect 41880 3130 41932 3136
rect 41694 3088 41750 3097
rect 41694 3023 41696 3032
rect 41748 3023 41750 3032
rect 41696 2994 41748 3000
rect 41616 2910 41736 2938
rect 41512 2372 41564 2378
rect 41512 2314 41564 2320
rect 41524 1698 41552 2314
rect 41512 1692 41564 1698
rect 41512 1634 41564 1640
rect 41708 56 41736 2910
rect 42076 56 42104 6190
rect 42248 3460 42300 3466
rect 42248 3402 42300 3408
rect 42260 3194 42288 3402
rect 42352 3210 42380 6258
rect 42430 4720 42486 4729
rect 42430 4655 42432 4664
rect 42484 4655 42486 4664
rect 42432 4626 42484 4632
rect 42248 3188 42300 3194
rect 42352 3182 42472 3210
rect 42248 3130 42300 3136
rect 42444 56 42472 3182
rect 42720 474 42748 7482
rect 43076 7404 43128 7410
rect 43076 7346 43128 7352
rect 42984 7200 43036 7206
rect 42984 7142 43036 7148
rect 42892 6724 42944 6730
rect 42892 6666 42944 6672
rect 42798 6352 42854 6361
rect 42798 6287 42800 6296
rect 42852 6287 42854 6296
rect 42800 6258 42852 6264
rect 42904 3346 42932 6666
rect 42812 3318 42932 3346
rect 42708 468 42760 474
rect 42708 410 42760 416
rect 42812 56 42840 3318
rect 42996 2938 43024 7142
rect 42904 2910 43024 2938
rect 42904 1630 42932 2910
rect 42984 2848 43036 2854
rect 42984 2790 43036 2796
rect 42996 2514 43024 2790
rect 43088 2774 43116 7346
rect 43260 6248 43312 6254
rect 43260 6190 43312 6196
rect 43166 5808 43222 5817
rect 43166 5743 43168 5752
rect 43220 5743 43222 5752
rect 43168 5714 43220 5720
rect 43272 5370 43300 6190
rect 43260 5364 43312 5370
rect 43260 5306 43312 5312
rect 43548 4826 43576 8366
rect 43640 7546 43668 9007
rect 43718 8800 43774 8809
rect 43718 8735 43774 8744
rect 43732 8090 43760 8735
rect 44100 8634 44128 11096
rect 44640 8968 44692 8974
rect 44640 8910 44692 8916
rect 44088 8628 44140 8634
rect 44088 8570 44140 8576
rect 43812 8492 43864 8498
rect 43812 8434 43864 8440
rect 43720 8084 43772 8090
rect 43720 8026 43772 8032
rect 43628 7540 43680 7546
rect 43628 7482 43680 7488
rect 43824 6458 43852 8434
rect 43950 8188 44258 8197
rect 43950 8186 43956 8188
rect 44012 8186 44036 8188
rect 44092 8186 44116 8188
rect 44172 8186 44196 8188
rect 44252 8186 44258 8188
rect 44012 8134 44014 8186
rect 44194 8134 44196 8186
rect 43950 8132 43956 8134
rect 44012 8132 44036 8134
rect 44092 8132 44116 8134
rect 44172 8132 44196 8134
rect 44252 8132 44258 8134
rect 43950 8123 44258 8132
rect 44548 7880 44600 7886
rect 44548 7822 44600 7828
rect 44272 7744 44324 7750
rect 44456 7744 44508 7750
rect 44272 7686 44324 7692
rect 44454 7712 44456 7721
rect 44508 7712 44510 7721
rect 44284 7449 44312 7686
rect 44454 7647 44510 7656
rect 44270 7440 44326 7449
rect 44270 7375 44326 7384
rect 44364 7404 44416 7410
rect 44364 7346 44416 7352
rect 43950 7100 44258 7109
rect 43950 7098 43956 7100
rect 44012 7098 44036 7100
rect 44092 7098 44116 7100
rect 44172 7098 44196 7100
rect 44252 7098 44258 7100
rect 44012 7046 44014 7098
rect 44194 7046 44196 7098
rect 43950 7044 43956 7046
rect 44012 7044 44036 7046
rect 44092 7044 44116 7046
rect 44172 7044 44196 7046
rect 44252 7044 44258 7046
rect 43950 7035 44258 7044
rect 44088 6656 44140 6662
rect 44086 6624 44088 6633
rect 44140 6624 44142 6633
rect 44086 6559 44142 6568
rect 43812 6452 43864 6458
rect 43812 6394 43864 6400
rect 44086 6216 44142 6225
rect 44086 6151 44088 6160
rect 44140 6151 44142 6160
rect 44088 6122 44140 6128
rect 43950 6012 44258 6021
rect 43950 6010 43956 6012
rect 44012 6010 44036 6012
rect 44092 6010 44116 6012
rect 44172 6010 44196 6012
rect 44252 6010 44258 6012
rect 44012 5958 44014 6010
rect 44194 5958 44196 6010
rect 43950 5956 43956 5958
rect 44012 5956 44036 5958
rect 44092 5956 44116 5958
rect 44172 5956 44196 5958
rect 44252 5956 44258 5958
rect 43950 5947 44258 5956
rect 43810 5672 43866 5681
rect 43810 5607 43866 5616
rect 43626 5264 43682 5273
rect 43626 5199 43682 5208
rect 43536 4820 43588 4826
rect 43536 4762 43588 4768
rect 43444 4140 43496 4146
rect 43444 4082 43496 4088
rect 43260 4072 43312 4078
rect 43260 4014 43312 4020
rect 43272 3738 43300 4014
rect 43260 3732 43312 3738
rect 43260 3674 43312 3680
rect 43258 3632 43314 3641
rect 43258 3567 43314 3576
rect 43352 3596 43404 3602
rect 43272 3058 43300 3567
rect 43352 3538 43404 3544
rect 43364 3058 43392 3538
rect 43456 3194 43484 4082
rect 43444 3188 43496 3194
rect 43444 3130 43496 3136
rect 43168 3052 43220 3058
rect 43168 2994 43220 3000
rect 43260 3052 43312 3058
rect 43260 2994 43312 3000
rect 43352 3052 43404 3058
rect 43352 2994 43404 3000
rect 43180 2961 43208 2994
rect 43166 2952 43222 2961
rect 43166 2887 43168 2896
rect 43220 2887 43222 2896
rect 43168 2858 43220 2864
rect 43272 2854 43300 2994
rect 43260 2848 43312 2854
rect 43260 2790 43312 2796
rect 43640 2774 43668 5199
rect 43088 2746 43208 2774
rect 42984 2508 43036 2514
rect 42984 2450 43036 2456
rect 42984 2304 43036 2310
rect 42984 2246 43036 2252
rect 42996 1737 43024 2246
rect 42982 1728 43038 1737
rect 42982 1663 43038 1672
rect 42892 1624 42944 1630
rect 42892 1566 42944 1572
rect 43180 56 43208 2746
rect 43548 2746 43668 2774
rect 43260 2440 43312 2446
rect 43260 2382 43312 2388
rect 43272 1834 43300 2382
rect 43352 2304 43404 2310
rect 43352 2246 43404 2252
rect 43260 1828 43312 1834
rect 43260 1770 43312 1776
rect 43364 1465 43392 2246
rect 43350 1456 43406 1465
rect 43350 1391 43406 1400
rect 43548 56 43576 2746
rect 43628 2440 43680 2446
rect 43628 2382 43680 2388
rect 43640 1329 43668 2382
rect 43824 1442 43852 5607
rect 44086 5128 44142 5137
rect 44086 5063 44088 5072
rect 44140 5063 44142 5072
rect 44088 5034 44140 5040
rect 43950 4924 44258 4933
rect 43950 4922 43956 4924
rect 44012 4922 44036 4924
rect 44092 4922 44116 4924
rect 44172 4922 44196 4924
rect 44252 4922 44258 4924
rect 44012 4870 44014 4922
rect 44194 4870 44196 4922
rect 43950 4868 43956 4870
rect 44012 4868 44036 4870
rect 44092 4868 44116 4870
rect 44172 4868 44196 4870
rect 44252 4868 44258 4870
rect 43950 4859 44258 4868
rect 44376 4758 44404 7346
rect 44456 7200 44508 7206
rect 44454 7168 44456 7177
rect 44508 7168 44510 7177
rect 44454 7103 44510 7112
rect 44454 6896 44510 6905
rect 44454 6831 44510 6840
rect 44468 6662 44496 6831
rect 44456 6656 44508 6662
rect 44456 6598 44508 6604
rect 44456 6452 44508 6458
rect 44456 6394 44508 6400
rect 44468 6361 44496 6394
rect 44454 6352 44510 6361
rect 44454 6287 44510 6296
rect 44456 5840 44508 5846
rect 44454 5808 44456 5817
rect 44508 5808 44510 5817
rect 44454 5743 44510 5752
rect 44456 5364 44508 5370
rect 44456 5306 44508 5312
rect 44468 5273 44496 5306
rect 44454 5264 44510 5273
rect 44454 5199 44510 5208
rect 44560 5030 44588 7822
rect 44652 6914 44680 8910
rect 44916 8560 44968 8566
rect 44916 8502 44968 8508
rect 44732 8356 44784 8362
rect 44732 8298 44784 8304
rect 44744 8265 44772 8298
rect 44730 8256 44786 8265
rect 44730 8191 44786 8200
rect 44928 7993 44956 8502
rect 44914 7984 44970 7993
rect 44914 7919 44970 7928
rect 44916 6996 44968 7002
rect 44916 6938 44968 6944
rect 44652 6886 44772 6914
rect 44640 5908 44692 5914
rect 44640 5850 44692 5856
rect 44548 5024 44600 5030
rect 44548 4966 44600 4972
rect 44364 4752 44416 4758
rect 44456 4752 44508 4758
rect 44364 4694 44416 4700
rect 44454 4720 44456 4729
rect 44508 4720 44510 4729
rect 44454 4655 44510 4664
rect 43904 4616 43956 4622
rect 43904 4558 43956 4564
rect 43916 4282 43944 4558
rect 44088 4480 44140 4486
rect 44086 4448 44088 4457
rect 44140 4448 44142 4457
rect 44086 4383 44142 4392
rect 43904 4276 43956 4282
rect 43904 4218 43956 4224
rect 44454 4176 44510 4185
rect 44454 4111 44510 4120
rect 44086 4040 44142 4049
rect 44468 4010 44496 4111
rect 44086 3975 44088 3984
rect 44140 3975 44142 3984
rect 44456 4004 44508 4010
rect 44088 3946 44140 3952
rect 44456 3946 44508 3952
rect 43950 3836 44258 3845
rect 43950 3834 43956 3836
rect 44012 3834 44036 3836
rect 44092 3834 44116 3836
rect 44172 3834 44196 3836
rect 44252 3834 44258 3836
rect 44012 3782 44014 3834
rect 44194 3782 44196 3834
rect 43950 3780 43956 3782
rect 44012 3780 44036 3782
rect 44092 3780 44116 3782
rect 44172 3780 44196 3782
rect 44252 3780 44258 3782
rect 43950 3771 44258 3780
rect 44456 3664 44508 3670
rect 44454 3632 44456 3641
rect 44508 3632 44510 3641
rect 44454 3567 44510 3576
rect 44088 3392 44140 3398
rect 44086 3360 44088 3369
rect 44140 3360 44142 3369
rect 44086 3295 44142 3304
rect 44652 3210 44680 5850
rect 44744 3534 44772 6886
rect 44824 5772 44876 5778
rect 44824 5714 44876 5720
rect 44836 4622 44864 5714
rect 44824 4616 44876 4622
rect 44824 4558 44876 4564
rect 44732 3528 44784 3534
rect 44732 3470 44784 3476
rect 44652 3182 44772 3210
rect 44640 3120 44692 3126
rect 44546 3088 44602 3097
rect 44640 3062 44692 3068
rect 44546 3023 44602 3032
rect 44364 2848 44416 2854
rect 44456 2848 44508 2854
rect 44364 2790 44416 2796
rect 44454 2816 44456 2825
rect 44508 2816 44510 2825
rect 43950 2748 44258 2757
rect 43950 2746 43956 2748
rect 44012 2746 44036 2748
rect 44092 2746 44116 2748
rect 44172 2746 44196 2748
rect 44252 2746 44258 2748
rect 44012 2694 44014 2746
rect 44194 2694 44196 2746
rect 43950 2692 43956 2694
rect 44012 2692 44036 2694
rect 44092 2692 44116 2694
rect 44172 2692 44196 2694
rect 44252 2692 44258 2694
rect 43950 2683 44258 2692
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 44192 2553 44220 2586
rect 44178 2544 44234 2553
rect 44178 2479 44234 2488
rect 44088 2304 44140 2310
rect 44086 2272 44088 2281
rect 44140 2272 44142 2281
rect 44086 2207 44142 2216
rect 44376 2009 44404 2790
rect 44454 2751 44510 2760
rect 44560 2650 44588 3023
rect 44548 2644 44600 2650
rect 44548 2586 44600 2592
rect 44652 2446 44680 3062
rect 44640 2440 44692 2446
rect 44640 2382 44692 2388
rect 44362 2000 44418 2009
rect 44362 1935 44418 1944
rect 44744 1442 44772 3182
rect 44928 2774 44956 6938
rect 45192 5568 45244 5574
rect 45190 5536 45192 5545
rect 45244 5536 45246 5545
rect 45190 5471 45246 5480
rect 45744 4548 45796 4554
rect 45744 4490 45796 4496
rect 44928 2746 45048 2774
rect 44824 2576 44876 2582
rect 44824 2518 44876 2524
rect 43824 1414 43944 1442
rect 43626 1320 43682 1329
rect 43626 1255 43682 1264
rect 43916 56 43944 1414
rect 44652 1414 44772 1442
rect 44272 1284 44324 1290
rect 44272 1226 44324 1232
rect 44284 56 44312 1226
rect 44652 56 44680 1414
rect 44836 1193 44864 2518
rect 44822 1184 44878 1193
rect 44822 1119 44878 1128
rect 45020 56 45048 2746
rect 45376 468 45428 474
rect 45376 410 45428 416
rect 45388 56 45416 410
rect 45756 56 45784 4490
rect 41052 2 41104 8
rect 41326 0 41382 56
rect 41694 0 41750 56
rect 42062 0 42118 56
rect 42430 0 42486 56
rect 42798 0 42854 56
rect 43166 0 43222 56
rect 43534 0 43590 56
rect 43902 0 43958 56
rect 44270 0 44326 56
rect 44638 0 44694 56
rect 45006 0 45062 56
rect 45374 0 45430 56
rect 45742 0 45798 56
<< via2 >>
rect 1214 9560 1270 9616
rect 754 9288 810 9344
rect 1030 8744 1086 8800
rect 2870 9016 2926 9072
rect 1306 8200 1362 8256
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2502 7928 2558 7984
rect 2686 7948 2742 7984
rect 2686 7928 2688 7948
rect 2688 7928 2740 7948
rect 2740 7928 2742 7948
rect 1214 7792 1270 7848
rect 1214 7656 1270 7712
rect 1122 7112 1178 7168
rect 1030 6568 1086 6624
rect 662 6024 718 6080
rect 386 1672 442 1728
rect 1306 7384 1362 7440
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1306 6840 1362 6896
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 2502 6704 2558 6760
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1306 5480 1362 5536
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2318 4548 2374 4584
rect 2318 4528 2320 4548
rect 2320 4528 2372 4548
rect 2372 4528 2374 4548
rect 754 4392 810 4448
rect 1306 4120 1362 4176
rect 1398 3984 1454 4040
rect 1398 3576 1454 3632
rect 1766 3440 1822 3496
rect 1122 1944 1178 2000
rect 1766 2760 1822 2816
rect 1306 2216 1362 2272
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 1214 1400 1270 1456
rect 1582 584 1638 640
rect 2594 1128 2650 1184
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 3238 5108 3240 5128
rect 3240 5108 3292 5128
rect 3292 5108 3294 5128
rect 3238 5072 3294 5108
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 2870 3984 2926 4040
rect 2870 3304 2926 3360
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 3698 3848 3754 3904
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 4342 5208 4398 5264
rect 5078 4936 5134 4992
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 5538 4664 5594 4720
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 10138 5208 10194 5264
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7194 1400 7250 1456
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 8574 1944 8630 2000
rect 10782 3168 10838 3224
rect 10414 176 10470 232
rect 12070 2488 12126 2544
rect 11886 1536 11942 1592
rect 11518 448 11574 504
rect 11150 312 11206 368
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 14094 40 14150 96
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 14738 3168 14794 3224
rect 14738 2760 14794 2816
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 15934 2352 15990 2408
rect 16578 1264 16634 1320
rect 15382 584 15438 640
rect 17958 4664 18014 4720
rect 17406 4120 17462 4176
rect 17774 1672 17830 1728
rect 18878 1808 18934 1864
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 19798 2760 19854 2816
rect 20350 2760 20406 2816
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 20902 1536 20958 1592
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 22466 6160 22522 6216
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 24122 1400 24178 1456
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25042 1944 25098 2000
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25778 2760 25834 2816
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 27618 448 27674 504
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 28170 1672 28226 1728
rect 28262 312 28318 368
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 29090 176 29146 232
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31482 4120 31538 4176
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 31482 1808 31538 1864
rect 32494 2388 32496 2408
rect 32496 2388 32548 2408
rect 32548 2388 32550 2408
rect 32494 2352 32550 2388
rect 32862 2488 32918 2544
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 34794 5208 34850 5264
rect 37278 5616 37334 5672
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 42982 9560 43038 9616
rect 41602 8472 41658 8528
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 38658 40 38714 96
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 43350 9288 43406 9344
rect 43258 8472 43314 8528
rect 43626 9016 43682 9072
rect 43166 7928 43222 7984
rect 42062 7828 42064 7848
rect 42064 7828 42116 7848
rect 42116 7828 42118 7848
rect 42062 7792 42118 7828
rect 39486 176 39542 232
rect 41050 4528 41106 4584
rect 41418 5072 41474 5128
rect 41510 3984 41566 4040
rect 41878 3440 41934 3496
rect 41694 3052 41750 3088
rect 41694 3032 41696 3052
rect 41696 3032 41748 3052
rect 41748 3032 41750 3052
rect 42430 4684 42486 4720
rect 42430 4664 42432 4684
rect 42432 4664 42484 4684
rect 42484 4664 42486 4684
rect 42798 6316 42854 6352
rect 42798 6296 42800 6316
rect 42800 6296 42852 6316
rect 42852 6296 42854 6316
rect 43166 5772 43222 5808
rect 43166 5752 43168 5772
rect 43168 5752 43220 5772
rect 43220 5752 43222 5772
rect 43718 8744 43774 8800
rect 43956 8186 44012 8188
rect 44036 8186 44092 8188
rect 44116 8186 44172 8188
rect 44196 8186 44252 8188
rect 43956 8134 44002 8186
rect 44002 8134 44012 8186
rect 44036 8134 44066 8186
rect 44066 8134 44078 8186
rect 44078 8134 44092 8186
rect 44116 8134 44130 8186
rect 44130 8134 44142 8186
rect 44142 8134 44172 8186
rect 44196 8134 44206 8186
rect 44206 8134 44252 8186
rect 43956 8132 44012 8134
rect 44036 8132 44092 8134
rect 44116 8132 44172 8134
rect 44196 8132 44252 8134
rect 44454 7692 44456 7712
rect 44456 7692 44508 7712
rect 44508 7692 44510 7712
rect 44454 7656 44510 7692
rect 44270 7384 44326 7440
rect 43956 7098 44012 7100
rect 44036 7098 44092 7100
rect 44116 7098 44172 7100
rect 44196 7098 44252 7100
rect 43956 7046 44002 7098
rect 44002 7046 44012 7098
rect 44036 7046 44066 7098
rect 44066 7046 44078 7098
rect 44078 7046 44092 7098
rect 44116 7046 44130 7098
rect 44130 7046 44142 7098
rect 44142 7046 44172 7098
rect 44196 7046 44206 7098
rect 44206 7046 44252 7098
rect 43956 7044 44012 7046
rect 44036 7044 44092 7046
rect 44116 7044 44172 7046
rect 44196 7044 44252 7046
rect 44086 6604 44088 6624
rect 44088 6604 44140 6624
rect 44140 6604 44142 6624
rect 44086 6568 44142 6604
rect 44086 6180 44142 6216
rect 44086 6160 44088 6180
rect 44088 6160 44140 6180
rect 44140 6160 44142 6180
rect 43956 6010 44012 6012
rect 44036 6010 44092 6012
rect 44116 6010 44172 6012
rect 44196 6010 44252 6012
rect 43956 5958 44002 6010
rect 44002 5958 44012 6010
rect 44036 5958 44066 6010
rect 44066 5958 44078 6010
rect 44078 5958 44092 6010
rect 44116 5958 44130 6010
rect 44130 5958 44142 6010
rect 44142 5958 44172 6010
rect 44196 5958 44206 6010
rect 44206 5958 44252 6010
rect 43956 5956 44012 5958
rect 44036 5956 44092 5958
rect 44116 5956 44172 5958
rect 44196 5956 44252 5958
rect 43810 5616 43866 5672
rect 43626 5208 43682 5264
rect 43258 3576 43314 3632
rect 43166 2916 43222 2952
rect 43166 2896 43168 2916
rect 43168 2896 43220 2916
rect 43220 2896 43222 2916
rect 42982 1672 43038 1728
rect 43350 1400 43406 1456
rect 44086 5092 44142 5128
rect 44086 5072 44088 5092
rect 44088 5072 44140 5092
rect 44140 5072 44142 5092
rect 43956 4922 44012 4924
rect 44036 4922 44092 4924
rect 44116 4922 44172 4924
rect 44196 4922 44252 4924
rect 43956 4870 44002 4922
rect 44002 4870 44012 4922
rect 44036 4870 44066 4922
rect 44066 4870 44078 4922
rect 44078 4870 44092 4922
rect 44116 4870 44130 4922
rect 44130 4870 44142 4922
rect 44142 4870 44172 4922
rect 44196 4870 44206 4922
rect 44206 4870 44252 4922
rect 43956 4868 44012 4870
rect 44036 4868 44092 4870
rect 44116 4868 44172 4870
rect 44196 4868 44252 4870
rect 44454 7148 44456 7168
rect 44456 7148 44508 7168
rect 44508 7148 44510 7168
rect 44454 7112 44510 7148
rect 44454 6840 44510 6896
rect 44454 6296 44510 6352
rect 44454 5788 44456 5808
rect 44456 5788 44508 5808
rect 44508 5788 44510 5808
rect 44454 5752 44510 5788
rect 44454 5208 44510 5264
rect 44730 8200 44786 8256
rect 44914 7928 44970 7984
rect 44454 4700 44456 4720
rect 44456 4700 44508 4720
rect 44508 4700 44510 4720
rect 44454 4664 44510 4700
rect 44086 4428 44088 4448
rect 44088 4428 44140 4448
rect 44140 4428 44142 4448
rect 44086 4392 44142 4428
rect 44454 4120 44510 4176
rect 44086 4004 44142 4040
rect 44086 3984 44088 4004
rect 44088 3984 44140 4004
rect 44140 3984 44142 4004
rect 43956 3834 44012 3836
rect 44036 3834 44092 3836
rect 44116 3834 44172 3836
rect 44196 3834 44252 3836
rect 43956 3782 44002 3834
rect 44002 3782 44012 3834
rect 44036 3782 44066 3834
rect 44066 3782 44078 3834
rect 44078 3782 44092 3834
rect 44116 3782 44130 3834
rect 44130 3782 44142 3834
rect 44142 3782 44172 3834
rect 44196 3782 44206 3834
rect 44206 3782 44252 3834
rect 43956 3780 44012 3782
rect 44036 3780 44092 3782
rect 44116 3780 44172 3782
rect 44196 3780 44252 3782
rect 44454 3612 44456 3632
rect 44456 3612 44508 3632
rect 44508 3612 44510 3632
rect 44454 3576 44510 3612
rect 44086 3340 44088 3360
rect 44088 3340 44140 3360
rect 44140 3340 44142 3360
rect 44086 3304 44142 3340
rect 44546 3032 44602 3088
rect 44454 2796 44456 2816
rect 44456 2796 44508 2816
rect 44508 2796 44510 2816
rect 43956 2746 44012 2748
rect 44036 2746 44092 2748
rect 44116 2746 44172 2748
rect 44196 2746 44252 2748
rect 43956 2694 44002 2746
rect 44002 2694 44012 2746
rect 44036 2694 44066 2746
rect 44066 2694 44078 2746
rect 44078 2694 44092 2746
rect 44116 2694 44130 2746
rect 44130 2694 44142 2746
rect 44142 2694 44172 2746
rect 44196 2694 44206 2746
rect 44206 2694 44252 2746
rect 43956 2692 44012 2694
rect 44036 2692 44092 2694
rect 44116 2692 44172 2694
rect 44196 2692 44252 2694
rect 44178 2488 44234 2544
rect 44086 2252 44088 2272
rect 44088 2252 44140 2272
rect 44140 2252 44142 2272
rect 44086 2216 44142 2252
rect 44454 2760 44510 2796
rect 44362 1944 44418 2000
rect 45190 5516 45192 5536
rect 45192 5516 45244 5536
rect 45244 5516 45246 5536
rect 45190 5480 45246 5516
rect 43626 1264 43682 1320
rect 44822 1128 44878 1184
<< metal3 >>
rect 0 9618 120 9648
rect 1209 9618 1275 9621
rect 0 9616 1275 9618
rect 0 9560 1214 9616
rect 1270 9560 1275 9616
rect 0 9558 1275 9560
rect 0 9528 120 9558
rect 1209 9555 1275 9558
rect 42977 9618 43043 9621
rect 45880 9618 46000 9648
rect 42977 9616 46000 9618
rect 42977 9560 42982 9616
rect 43038 9560 46000 9616
rect 42977 9558 46000 9560
rect 42977 9555 43043 9558
rect 45880 9528 46000 9558
rect 0 9346 120 9376
rect 749 9346 815 9349
rect 0 9344 815 9346
rect 0 9288 754 9344
rect 810 9288 815 9344
rect 0 9286 815 9288
rect 0 9256 120 9286
rect 749 9283 815 9286
rect 43345 9346 43411 9349
rect 45880 9346 46000 9376
rect 43345 9344 46000 9346
rect 43345 9288 43350 9344
rect 43406 9288 46000 9344
rect 43345 9286 46000 9288
rect 43345 9283 43411 9286
rect 45880 9256 46000 9286
rect 0 9074 120 9104
rect 2865 9074 2931 9077
rect 0 9072 2931 9074
rect 0 9016 2870 9072
rect 2926 9016 2931 9072
rect 0 9014 2931 9016
rect 0 8984 120 9014
rect 2865 9011 2931 9014
rect 43621 9074 43687 9077
rect 45880 9074 46000 9104
rect 43621 9072 46000 9074
rect 43621 9016 43626 9072
rect 43682 9016 46000 9072
rect 43621 9014 46000 9016
rect 43621 9011 43687 9014
rect 45880 8984 46000 9014
rect 0 8802 120 8832
rect 1025 8802 1091 8805
rect 0 8800 1091 8802
rect 0 8744 1030 8800
rect 1086 8744 1091 8800
rect 0 8742 1091 8744
rect 0 8712 120 8742
rect 1025 8739 1091 8742
rect 43713 8802 43779 8805
rect 45880 8802 46000 8832
rect 43713 8800 46000 8802
rect 43713 8744 43718 8800
rect 43774 8744 46000 8800
rect 43713 8742 46000 8744
rect 43713 8739 43779 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 45880 8712 46000 8742
rect 39006 8671 39322 8672
rect 0 8530 120 8560
rect 41597 8530 41663 8533
rect 0 8528 41663 8530
rect 0 8472 41602 8528
rect 41658 8472 41663 8528
rect 0 8470 41663 8472
rect 0 8440 120 8470
rect 41597 8467 41663 8470
rect 43253 8530 43319 8533
rect 45880 8530 46000 8560
rect 43253 8528 46000 8530
rect 43253 8472 43258 8528
rect 43314 8472 46000 8528
rect 43253 8470 46000 8472
rect 43253 8467 43319 8470
rect 45880 8440 46000 8470
rect 0 8258 120 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 0 8168 120 8198
rect 1301 8195 1367 8198
rect 44725 8258 44791 8261
rect 45880 8258 46000 8288
rect 44725 8256 46000 8258
rect 44725 8200 44730 8256
rect 44786 8200 46000 8256
rect 44725 8198 46000 8200
rect 44725 8195 44791 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 37946 8127 38262 8128
rect 43946 8192 44262 8193
rect 43946 8128 43952 8192
rect 44016 8128 44032 8192
rect 44096 8128 44112 8192
rect 44176 8128 44192 8192
rect 44256 8128 44262 8192
rect 45880 8168 46000 8198
rect 43946 8127 44262 8128
rect 0 7986 120 8016
rect 2497 7986 2563 7989
rect 0 7984 2563 7986
rect 0 7928 2502 7984
rect 2558 7928 2563 7984
rect 0 7926 2563 7928
rect 0 7896 120 7926
rect 2497 7923 2563 7926
rect 2681 7986 2747 7989
rect 43161 7986 43227 7989
rect 2681 7984 43227 7986
rect 2681 7928 2686 7984
rect 2742 7928 43166 7984
rect 43222 7928 43227 7984
rect 2681 7926 43227 7928
rect 2681 7923 2747 7926
rect 43161 7923 43227 7926
rect 44909 7986 44975 7989
rect 45880 7986 46000 8016
rect 44909 7984 46000 7986
rect 44909 7928 44914 7984
rect 44970 7928 46000 7984
rect 44909 7926 46000 7928
rect 44909 7923 44975 7926
rect 45880 7896 46000 7926
rect 1209 7850 1275 7853
rect 42057 7850 42123 7853
rect 1209 7848 42123 7850
rect 1209 7792 1214 7848
rect 1270 7792 42062 7848
rect 42118 7792 42123 7848
rect 1209 7790 42123 7792
rect 1209 7787 1275 7790
rect 42057 7787 42123 7790
rect 0 7714 120 7744
rect 1209 7714 1275 7717
rect 0 7712 1275 7714
rect 0 7656 1214 7712
rect 1270 7656 1275 7712
rect 0 7654 1275 7656
rect 0 7624 120 7654
rect 1209 7651 1275 7654
rect 44449 7714 44515 7717
rect 45880 7714 46000 7744
rect 44449 7712 46000 7714
rect 44449 7656 44454 7712
rect 44510 7656 46000 7712
rect 44449 7654 46000 7656
rect 44449 7651 44515 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 45880 7624 46000 7654
rect 39006 7583 39322 7584
rect 0 7442 120 7472
rect 1301 7442 1367 7445
rect 0 7440 1367 7442
rect 0 7384 1306 7440
rect 1362 7384 1367 7440
rect 0 7382 1367 7384
rect 0 7352 120 7382
rect 1301 7379 1367 7382
rect 44265 7442 44331 7445
rect 45880 7442 46000 7472
rect 44265 7440 46000 7442
rect 44265 7384 44270 7440
rect 44326 7384 46000 7440
rect 44265 7382 46000 7384
rect 44265 7379 44331 7382
rect 45880 7352 46000 7382
rect 0 7170 120 7200
rect 1117 7170 1183 7173
rect 0 7168 1183 7170
rect 0 7112 1122 7168
rect 1178 7112 1183 7168
rect 0 7110 1183 7112
rect 0 7080 120 7110
rect 1117 7107 1183 7110
rect 44449 7170 44515 7173
rect 45880 7170 46000 7200
rect 44449 7168 46000 7170
rect 44449 7112 44454 7168
rect 44510 7112 46000 7168
rect 44449 7110 46000 7112
rect 44449 7107 44515 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 37946 7039 38262 7040
rect 43946 7104 44262 7105
rect 43946 7040 43952 7104
rect 44016 7040 44032 7104
rect 44096 7040 44112 7104
rect 44176 7040 44192 7104
rect 44256 7040 44262 7104
rect 45880 7080 46000 7110
rect 43946 7039 44262 7040
rect 0 6898 120 6928
rect 1301 6898 1367 6901
rect 0 6896 1367 6898
rect 0 6840 1306 6896
rect 1362 6840 1367 6896
rect 0 6838 1367 6840
rect 0 6808 120 6838
rect 1301 6835 1367 6838
rect 44449 6898 44515 6901
rect 45880 6898 46000 6928
rect 44449 6896 46000 6898
rect 44449 6840 44454 6896
rect 44510 6840 46000 6896
rect 44449 6838 46000 6840
rect 44449 6835 44515 6838
rect 45880 6808 46000 6838
rect 2497 6762 2563 6765
rect 2497 6760 12450 6762
rect 2497 6704 2502 6760
rect 2558 6704 12450 6760
rect 2497 6702 12450 6704
rect 2497 6699 2563 6702
rect 0 6626 120 6656
rect 1025 6626 1091 6629
rect 0 6624 1091 6626
rect 0 6568 1030 6624
rect 1086 6568 1091 6624
rect 0 6566 1091 6568
rect 0 6536 120 6566
rect 1025 6563 1091 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 0 6354 120 6384
rect 12390 6354 12450 6702
rect 44081 6626 44147 6629
rect 45880 6626 46000 6656
rect 44081 6624 46000 6626
rect 44081 6568 44086 6624
rect 44142 6568 46000 6624
rect 44081 6566 46000 6568
rect 44081 6563 44147 6566
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 45880 6536 46000 6566
rect 39006 6495 39322 6496
rect 42793 6354 42859 6357
rect 0 6294 2790 6354
rect 12390 6352 42859 6354
rect 12390 6296 42798 6352
rect 42854 6296 42859 6352
rect 12390 6294 42859 6296
rect 0 6264 120 6294
rect 2730 6218 2790 6294
rect 42793 6291 42859 6294
rect 44449 6354 44515 6357
rect 45880 6354 46000 6384
rect 44449 6352 46000 6354
rect 44449 6296 44454 6352
rect 44510 6296 46000 6352
rect 44449 6294 46000 6296
rect 44449 6291 44515 6294
rect 45880 6264 46000 6294
rect 22461 6218 22527 6221
rect 2730 6216 22527 6218
rect 2730 6160 22466 6216
rect 22522 6160 22527 6216
rect 2730 6158 22527 6160
rect 22461 6155 22527 6158
rect 44081 6218 44147 6221
rect 44081 6216 45018 6218
rect 44081 6160 44086 6216
rect 44142 6160 45018 6216
rect 44081 6158 45018 6160
rect 44081 6155 44147 6158
rect 0 6082 120 6112
rect 657 6082 723 6085
rect 0 6080 723 6082
rect 0 6024 662 6080
rect 718 6024 723 6080
rect 0 6022 723 6024
rect 44958 6082 45018 6158
rect 45880 6082 46000 6112
rect 44958 6022 46000 6082
rect 0 5992 120 6022
rect 657 6019 723 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 37946 5951 38262 5952
rect 43946 6016 44262 6017
rect 43946 5952 43952 6016
rect 44016 5952 44032 6016
rect 44096 5952 44112 6016
rect 44176 5952 44192 6016
rect 44256 5952 44262 6016
rect 45880 5992 46000 6022
rect 43946 5951 44262 5952
rect 0 5810 120 5840
rect 43161 5810 43227 5813
rect 0 5808 43227 5810
rect 0 5752 43166 5808
rect 43222 5752 43227 5808
rect 0 5750 43227 5752
rect 0 5720 120 5750
rect 43161 5747 43227 5750
rect 44449 5810 44515 5813
rect 45880 5810 46000 5840
rect 44449 5808 46000 5810
rect 44449 5752 44454 5808
rect 44510 5752 46000 5808
rect 44449 5750 46000 5752
rect 44449 5747 44515 5750
rect 45880 5720 46000 5750
rect 37273 5674 37339 5677
rect 43805 5674 43871 5677
rect 37273 5672 43871 5674
rect 37273 5616 37278 5672
rect 37334 5616 43810 5672
rect 43866 5616 43871 5672
rect 37273 5614 43871 5616
rect 37273 5611 37339 5614
rect 43805 5611 43871 5614
rect 0 5538 120 5568
rect 1301 5538 1367 5541
rect 0 5536 1367 5538
rect 0 5480 1306 5536
rect 1362 5480 1367 5536
rect 0 5478 1367 5480
rect 0 5448 120 5478
rect 1301 5475 1367 5478
rect 45185 5538 45251 5541
rect 45880 5538 46000 5568
rect 45185 5536 46000 5538
rect 45185 5480 45190 5536
rect 45246 5480 46000 5536
rect 45185 5478 46000 5480
rect 45185 5475 45251 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 45880 5448 46000 5478
rect 39006 5407 39322 5408
rect 0 5266 120 5296
rect 4337 5266 4403 5269
rect 0 5264 4403 5266
rect 0 5208 4342 5264
rect 4398 5208 4403 5264
rect 0 5206 4403 5208
rect 0 5176 120 5206
rect 4337 5203 4403 5206
rect 10133 5266 10199 5269
rect 30966 5266 30972 5268
rect 10133 5264 30972 5266
rect 10133 5208 10138 5264
rect 10194 5208 30972 5264
rect 10133 5206 30972 5208
rect 10133 5203 10199 5206
rect 30966 5204 30972 5206
rect 31036 5204 31042 5268
rect 34789 5266 34855 5269
rect 43621 5266 43687 5269
rect 34789 5264 43687 5266
rect 34789 5208 34794 5264
rect 34850 5208 43626 5264
rect 43682 5208 43687 5264
rect 34789 5206 43687 5208
rect 34789 5203 34855 5206
rect 43621 5203 43687 5206
rect 44449 5266 44515 5269
rect 45880 5266 46000 5296
rect 44449 5264 46000 5266
rect 44449 5208 44454 5264
rect 44510 5208 46000 5264
rect 44449 5206 46000 5208
rect 44449 5203 44515 5206
rect 45880 5176 46000 5206
rect 3233 5130 3299 5133
rect 41413 5130 41479 5133
rect 1718 5070 2514 5130
rect 0 4994 120 5024
rect 1718 4994 1778 5070
rect 0 4934 1778 4994
rect 2454 4994 2514 5070
rect 3233 5128 41479 5130
rect 3233 5072 3238 5128
rect 3294 5072 41418 5128
rect 41474 5072 41479 5128
rect 3233 5070 41479 5072
rect 3233 5067 3299 5070
rect 41413 5067 41479 5070
rect 44081 5130 44147 5133
rect 44081 5128 45018 5130
rect 44081 5072 44086 5128
rect 44142 5072 45018 5128
rect 44081 5070 45018 5072
rect 44081 5067 44147 5070
rect 5073 4994 5139 4997
rect 2454 4992 5139 4994
rect 2454 4936 5078 4992
rect 5134 4936 5139 4992
rect 2454 4934 5139 4936
rect 44958 4994 45018 5070
rect 45880 4994 46000 5024
rect 44958 4934 46000 4994
rect 0 4904 120 4934
rect 5073 4931 5139 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 37946 4863 38262 4864
rect 43946 4928 44262 4929
rect 43946 4864 43952 4928
rect 44016 4864 44032 4928
rect 44096 4864 44112 4928
rect 44176 4864 44192 4928
rect 44256 4864 44262 4928
rect 45880 4904 46000 4934
rect 43946 4863 44262 4864
rect 0 4722 120 4752
rect 5533 4722 5599 4725
rect 0 4720 5599 4722
rect 0 4664 5538 4720
rect 5594 4664 5599 4720
rect 0 4662 5599 4664
rect 0 4632 120 4662
rect 5533 4659 5599 4662
rect 17953 4722 18019 4725
rect 42425 4722 42491 4725
rect 17953 4720 42491 4722
rect 17953 4664 17958 4720
rect 18014 4664 42430 4720
rect 42486 4664 42491 4720
rect 17953 4662 42491 4664
rect 17953 4659 18019 4662
rect 42425 4659 42491 4662
rect 44449 4722 44515 4725
rect 45880 4722 46000 4752
rect 44449 4720 46000 4722
rect 44449 4664 44454 4720
rect 44510 4664 46000 4720
rect 44449 4662 46000 4664
rect 44449 4659 44515 4662
rect 45880 4632 46000 4662
rect 2313 4586 2379 4589
rect 41045 4586 41111 4589
rect 2313 4584 41111 4586
rect 2313 4528 2318 4584
rect 2374 4528 41050 4584
rect 41106 4528 41111 4584
rect 2313 4526 41111 4528
rect 2313 4523 2379 4526
rect 41045 4523 41111 4526
rect 0 4450 120 4480
rect 749 4450 815 4453
rect 0 4448 815 4450
rect 0 4392 754 4448
rect 810 4392 815 4448
rect 0 4390 815 4392
rect 0 4360 120 4390
rect 749 4387 815 4390
rect 44081 4450 44147 4453
rect 45880 4450 46000 4480
rect 44081 4448 46000 4450
rect 44081 4392 44086 4448
rect 44142 4392 46000 4448
rect 44081 4390 46000 4392
rect 44081 4387 44147 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 45880 4360 46000 4390
rect 39006 4319 39322 4320
rect 0 4178 120 4208
rect 1301 4178 1367 4181
rect 0 4176 1367 4178
rect 0 4120 1306 4176
rect 1362 4120 1367 4176
rect 0 4118 1367 4120
rect 0 4088 120 4118
rect 1301 4115 1367 4118
rect 17401 4178 17467 4181
rect 31477 4178 31543 4181
rect 17401 4176 31543 4178
rect 17401 4120 17406 4176
rect 17462 4120 31482 4176
rect 31538 4120 31543 4176
rect 17401 4118 31543 4120
rect 17401 4115 17467 4118
rect 31477 4115 31543 4118
rect 44449 4178 44515 4181
rect 45880 4178 46000 4208
rect 44449 4176 46000 4178
rect 44449 4120 44454 4176
rect 44510 4120 46000 4176
rect 44449 4118 46000 4120
rect 44449 4115 44515 4118
rect 45880 4088 46000 4118
rect 1393 4042 1459 4045
rect 2865 4042 2931 4045
rect 41505 4042 41571 4045
rect 1393 4040 2514 4042
rect 1393 3984 1398 4040
rect 1454 3984 2514 4040
rect 1393 3982 2514 3984
rect 1393 3979 1459 3982
rect 0 3906 120 3936
rect 2454 3906 2514 3982
rect 2865 4040 41571 4042
rect 2865 3984 2870 4040
rect 2926 3984 41510 4040
rect 41566 3984 41571 4040
rect 2865 3982 41571 3984
rect 2865 3979 2931 3982
rect 41505 3979 41571 3982
rect 44081 4042 44147 4045
rect 44081 4040 45018 4042
rect 44081 3984 44086 4040
rect 44142 3984 45018 4040
rect 44081 3982 45018 3984
rect 44081 3979 44147 3982
rect 3693 3906 3759 3909
rect 0 3846 1778 3906
rect 2454 3904 3759 3906
rect 2454 3848 3698 3904
rect 3754 3848 3759 3904
rect 2454 3846 3759 3848
rect 44958 3906 45018 3982
rect 45880 3906 46000 3936
rect 44958 3846 46000 3906
rect 0 3816 120 3846
rect 0 3634 120 3664
rect 1393 3634 1459 3637
rect 0 3632 1459 3634
rect 0 3576 1398 3632
rect 1454 3576 1459 3632
rect 0 3574 1459 3576
rect 1718 3634 1778 3846
rect 3693 3843 3759 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 37946 3775 38262 3776
rect 43946 3840 44262 3841
rect 43946 3776 43952 3840
rect 44016 3776 44032 3840
rect 44096 3776 44112 3840
rect 44176 3776 44192 3840
rect 44256 3776 44262 3840
rect 45880 3816 46000 3846
rect 43946 3775 44262 3776
rect 43253 3634 43319 3637
rect 1718 3632 43319 3634
rect 1718 3576 43258 3632
rect 43314 3576 43319 3632
rect 1718 3574 43319 3576
rect 0 3544 120 3574
rect 1393 3571 1459 3574
rect 43253 3571 43319 3574
rect 44449 3634 44515 3637
rect 45880 3634 46000 3664
rect 44449 3632 46000 3634
rect 44449 3576 44454 3632
rect 44510 3576 46000 3632
rect 44449 3574 46000 3576
rect 44449 3571 44515 3574
rect 45880 3544 46000 3574
rect 1761 3498 1827 3501
rect 41873 3498 41939 3501
rect 1761 3496 41939 3498
rect 1761 3440 1766 3496
rect 1822 3440 41878 3496
rect 41934 3440 41939 3496
rect 1761 3438 41939 3440
rect 1761 3435 1827 3438
rect 41873 3435 41939 3438
rect 0 3362 120 3392
rect 2865 3362 2931 3365
rect 0 3360 2931 3362
rect 0 3304 2870 3360
rect 2926 3304 2931 3360
rect 0 3302 2931 3304
rect 0 3272 120 3302
rect 2865 3299 2931 3302
rect 44081 3362 44147 3365
rect 45880 3362 46000 3392
rect 44081 3360 46000 3362
rect 44081 3304 44086 3360
rect 44142 3304 46000 3360
rect 44081 3302 46000 3304
rect 44081 3299 44147 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 45880 3272 46000 3302
rect 39006 3231 39322 3232
rect 10777 3226 10843 3229
rect 14733 3226 14799 3229
rect 10777 3224 14799 3226
rect 10777 3168 10782 3224
rect 10838 3168 14738 3224
rect 14794 3168 14799 3224
rect 10777 3166 14799 3168
rect 10777 3163 10843 3166
rect 14733 3163 14799 3166
rect 0 3090 120 3120
rect 41689 3090 41755 3093
rect 0 3088 41755 3090
rect 0 3032 41694 3088
rect 41750 3032 41755 3088
rect 0 3030 41755 3032
rect 0 3000 120 3030
rect 41689 3027 41755 3030
rect 44541 3090 44607 3093
rect 45880 3090 46000 3120
rect 44541 3088 46000 3090
rect 44541 3032 44546 3088
rect 44602 3032 46000 3088
rect 44541 3030 46000 3032
rect 44541 3027 44607 3030
rect 45880 3000 46000 3030
rect 43161 2954 43227 2957
rect 9630 2952 43227 2954
rect 9630 2896 43166 2952
rect 43222 2896 43227 2952
rect 9630 2894 43227 2896
rect 0 2818 120 2848
rect 1761 2818 1827 2821
rect 0 2816 1827 2818
rect 0 2760 1766 2816
rect 1822 2760 1827 2816
rect 0 2758 1827 2760
rect 0 2728 120 2758
rect 1761 2755 1827 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 0 2546 120 2576
rect 9630 2546 9690 2894
rect 43161 2891 43227 2894
rect 14733 2818 14799 2821
rect 19793 2818 19859 2821
rect 14733 2816 19859 2818
rect 14733 2760 14738 2816
rect 14794 2760 19798 2816
rect 19854 2760 19859 2816
rect 14733 2758 19859 2760
rect 14733 2755 14799 2758
rect 19793 2755 19859 2758
rect 20345 2818 20411 2821
rect 25773 2818 25839 2821
rect 20345 2816 25839 2818
rect 20345 2760 20350 2816
rect 20406 2760 25778 2816
rect 25834 2760 25839 2816
rect 20345 2758 25839 2760
rect 20345 2755 20411 2758
rect 25773 2755 25839 2758
rect 44449 2818 44515 2821
rect 45880 2818 46000 2848
rect 44449 2816 46000 2818
rect 44449 2760 44454 2816
rect 44510 2760 46000 2816
rect 44449 2758 46000 2760
rect 44449 2755 44515 2758
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 37946 2687 38262 2688
rect 43946 2752 44262 2753
rect 43946 2688 43952 2752
rect 44016 2688 44032 2752
rect 44096 2688 44112 2752
rect 44176 2688 44192 2752
rect 44256 2688 44262 2752
rect 45880 2728 46000 2758
rect 43946 2687 44262 2688
rect 0 2486 9690 2546
rect 12065 2546 12131 2549
rect 32857 2546 32923 2549
rect 12065 2544 32923 2546
rect 12065 2488 12070 2544
rect 12126 2488 32862 2544
rect 32918 2488 32923 2544
rect 12065 2486 32923 2488
rect 0 2456 120 2486
rect 12065 2483 12131 2486
rect 32857 2483 32923 2486
rect 44173 2546 44239 2549
rect 45880 2546 46000 2576
rect 44173 2544 46000 2546
rect 44173 2488 44178 2544
rect 44234 2488 46000 2544
rect 44173 2486 46000 2488
rect 44173 2483 44239 2486
rect 45880 2456 46000 2486
rect 15929 2410 15995 2413
rect 32489 2410 32555 2413
rect 15929 2408 32555 2410
rect 15929 2352 15934 2408
rect 15990 2352 32494 2408
rect 32550 2352 32555 2408
rect 15929 2350 32555 2352
rect 15929 2347 15995 2350
rect 32489 2347 32555 2350
rect 0 2274 120 2304
rect 1301 2274 1367 2277
rect 0 2272 1367 2274
rect 0 2216 1306 2272
rect 1362 2216 1367 2272
rect 0 2214 1367 2216
rect 0 2184 120 2214
rect 1301 2211 1367 2214
rect 44081 2274 44147 2277
rect 45880 2274 46000 2304
rect 44081 2272 46000 2274
rect 44081 2216 44086 2272
rect 44142 2216 46000 2272
rect 44081 2214 46000 2216
rect 44081 2211 44147 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 45880 2184 46000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 1117 2002 1183 2005
rect 0 2000 1183 2002
rect 0 1944 1122 2000
rect 1178 1944 1183 2000
rect 0 1942 1183 1944
rect 0 1912 120 1942
rect 1117 1939 1183 1942
rect 8569 2002 8635 2005
rect 25037 2002 25103 2005
rect 8569 2000 25103 2002
rect 8569 1944 8574 2000
rect 8630 1944 25042 2000
rect 25098 1944 25103 2000
rect 8569 1942 25103 1944
rect 8569 1939 8635 1942
rect 25037 1939 25103 1942
rect 44357 2002 44423 2005
rect 45880 2002 46000 2032
rect 44357 2000 46000 2002
rect 44357 1944 44362 2000
rect 44418 1944 46000 2000
rect 44357 1942 46000 1944
rect 44357 1939 44423 1942
rect 45880 1912 46000 1942
rect 18873 1866 18939 1869
rect 31477 1866 31543 1869
rect 18873 1864 31543 1866
rect 18873 1808 18878 1864
rect 18934 1808 31482 1864
rect 31538 1808 31543 1864
rect 18873 1806 31543 1808
rect 18873 1803 18939 1806
rect 31477 1803 31543 1806
rect 0 1730 120 1760
rect 381 1730 447 1733
rect 0 1728 447 1730
rect 0 1672 386 1728
rect 442 1672 447 1728
rect 0 1670 447 1672
rect 0 1640 120 1670
rect 381 1667 447 1670
rect 17769 1730 17835 1733
rect 28165 1730 28231 1733
rect 17769 1728 28231 1730
rect 17769 1672 17774 1728
rect 17830 1672 28170 1728
rect 28226 1672 28231 1728
rect 17769 1670 28231 1672
rect 17769 1667 17835 1670
rect 28165 1667 28231 1670
rect 42977 1730 43043 1733
rect 45880 1730 46000 1760
rect 42977 1728 46000 1730
rect 42977 1672 42982 1728
rect 43038 1672 46000 1728
rect 42977 1670 46000 1672
rect 42977 1667 43043 1670
rect 45880 1640 46000 1670
rect 11881 1594 11947 1597
rect 20897 1594 20963 1597
rect 11881 1592 20963 1594
rect 11881 1536 11886 1592
rect 11942 1536 20902 1592
rect 20958 1536 20963 1592
rect 11881 1534 20963 1536
rect 11881 1531 11947 1534
rect 20897 1531 20963 1534
rect 0 1458 120 1488
rect 1209 1458 1275 1461
rect 0 1456 1275 1458
rect 0 1400 1214 1456
rect 1270 1400 1275 1456
rect 0 1398 1275 1400
rect 0 1368 120 1398
rect 1209 1395 1275 1398
rect 7189 1458 7255 1461
rect 24117 1458 24183 1461
rect 7189 1456 24183 1458
rect 7189 1400 7194 1456
rect 7250 1400 24122 1456
rect 24178 1400 24183 1456
rect 7189 1398 24183 1400
rect 7189 1395 7255 1398
rect 24117 1395 24183 1398
rect 43345 1458 43411 1461
rect 45880 1458 46000 1488
rect 43345 1456 46000 1458
rect 43345 1400 43350 1456
rect 43406 1400 46000 1456
rect 43345 1398 46000 1400
rect 43345 1395 43411 1398
rect 45880 1368 46000 1398
rect 16573 1322 16639 1325
rect 43621 1322 43687 1325
rect 16573 1320 43687 1322
rect 16573 1264 16578 1320
rect 16634 1264 43626 1320
rect 43682 1264 43687 1320
rect 16573 1262 43687 1264
rect 16573 1259 16639 1262
rect 43621 1259 43687 1262
rect 0 1186 120 1216
rect 2589 1186 2655 1189
rect 0 1184 2655 1186
rect 0 1128 2594 1184
rect 2650 1128 2655 1184
rect 0 1126 2655 1128
rect 0 1096 120 1126
rect 2589 1123 2655 1126
rect 44817 1186 44883 1189
rect 45880 1186 46000 1216
rect 44817 1184 46000 1186
rect 44817 1128 44822 1184
rect 44878 1128 46000 1184
rect 44817 1126 46000 1128
rect 44817 1123 44883 1126
rect 45880 1096 46000 1126
rect 1577 642 1643 645
rect 15377 642 15443 645
rect 1577 640 15443 642
rect 1577 584 1582 640
rect 1638 584 15382 640
rect 15438 584 15443 640
rect 1577 582 15443 584
rect 1577 579 1643 582
rect 15377 579 15443 582
rect 11513 506 11579 509
rect 27613 506 27679 509
rect 11513 504 27679 506
rect 11513 448 11518 504
rect 11574 448 27618 504
rect 27674 448 27679 504
rect 11513 446 27679 448
rect 11513 443 11579 446
rect 27613 443 27679 446
rect 11145 370 11211 373
rect 28257 370 28323 373
rect 11145 368 28323 370
rect 11145 312 11150 368
rect 11206 312 28262 368
rect 28318 312 28323 368
rect 11145 310 28323 312
rect 11145 307 11211 310
rect 28257 307 28323 310
rect 10409 234 10475 237
rect 29085 234 29151 237
rect 10409 232 29151 234
rect 10409 176 10414 232
rect 10470 176 29090 232
rect 29146 176 29151 232
rect 10409 174 29151 176
rect 10409 171 10475 174
rect 29085 171 29151 174
rect 30966 172 30972 236
rect 31036 234 31042 236
rect 39481 234 39547 237
rect 31036 232 39547 234
rect 31036 176 39486 232
rect 39542 176 39547 232
rect 31036 174 39547 176
rect 31036 172 31042 174
rect 39481 171 39547 174
rect 14089 98 14155 101
rect 38653 98 38719 101
rect 14089 96 38719 98
rect 14089 40 14094 96
rect 14150 40 38658 96
rect 38714 40 38719 96
rect 14089 38 38719 40
rect 14089 35 14155 38
rect 38653 35 38719 38
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 43952 8188 44016 8192
rect 43952 8132 43956 8188
rect 43956 8132 44012 8188
rect 44012 8132 44016 8188
rect 43952 8128 44016 8132
rect 44032 8188 44096 8192
rect 44032 8132 44036 8188
rect 44036 8132 44092 8188
rect 44092 8132 44096 8188
rect 44032 8128 44096 8132
rect 44112 8188 44176 8192
rect 44112 8132 44116 8188
rect 44116 8132 44172 8188
rect 44172 8132 44176 8188
rect 44112 8128 44176 8132
rect 44192 8188 44256 8192
rect 44192 8132 44196 8188
rect 44196 8132 44252 8188
rect 44252 8132 44256 8188
rect 44192 8128 44256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 43952 7100 44016 7104
rect 43952 7044 43956 7100
rect 43956 7044 44012 7100
rect 44012 7044 44016 7100
rect 43952 7040 44016 7044
rect 44032 7100 44096 7104
rect 44032 7044 44036 7100
rect 44036 7044 44092 7100
rect 44092 7044 44096 7100
rect 44032 7040 44096 7044
rect 44112 7100 44176 7104
rect 44112 7044 44116 7100
rect 44116 7044 44172 7100
rect 44172 7044 44176 7100
rect 44112 7040 44176 7044
rect 44192 7100 44256 7104
rect 44192 7044 44196 7100
rect 44196 7044 44252 7100
rect 44252 7044 44256 7100
rect 44192 7040 44256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 43952 6012 44016 6016
rect 43952 5956 43956 6012
rect 43956 5956 44012 6012
rect 44012 5956 44016 6012
rect 43952 5952 44016 5956
rect 44032 6012 44096 6016
rect 44032 5956 44036 6012
rect 44036 5956 44092 6012
rect 44092 5956 44096 6012
rect 44032 5952 44096 5956
rect 44112 6012 44176 6016
rect 44112 5956 44116 6012
rect 44116 5956 44172 6012
rect 44172 5956 44176 6012
rect 44112 5952 44176 5956
rect 44192 6012 44256 6016
rect 44192 5956 44196 6012
rect 44196 5956 44252 6012
rect 44252 5956 44256 6012
rect 44192 5952 44256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 30972 5204 31036 5268
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 43952 4924 44016 4928
rect 43952 4868 43956 4924
rect 43956 4868 44012 4924
rect 44012 4868 44016 4924
rect 43952 4864 44016 4868
rect 44032 4924 44096 4928
rect 44032 4868 44036 4924
rect 44036 4868 44092 4924
rect 44092 4868 44096 4924
rect 44032 4864 44096 4868
rect 44112 4924 44176 4928
rect 44112 4868 44116 4924
rect 44116 4868 44172 4924
rect 44172 4868 44176 4924
rect 44112 4864 44176 4868
rect 44192 4924 44256 4928
rect 44192 4868 44196 4924
rect 44196 4868 44252 4924
rect 44252 4868 44256 4924
rect 44192 4864 44256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 43952 3836 44016 3840
rect 43952 3780 43956 3836
rect 43956 3780 44012 3836
rect 44012 3780 44016 3836
rect 43952 3776 44016 3780
rect 44032 3836 44096 3840
rect 44032 3780 44036 3836
rect 44036 3780 44092 3836
rect 44092 3780 44096 3836
rect 44032 3776 44096 3780
rect 44112 3836 44176 3840
rect 44112 3780 44116 3836
rect 44116 3780 44172 3836
rect 44172 3780 44176 3836
rect 44112 3776 44176 3780
rect 44192 3836 44256 3840
rect 44192 3780 44196 3836
rect 44196 3780 44252 3836
rect 44252 3780 44256 3836
rect 44192 3776 44256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 43952 2748 44016 2752
rect 43952 2692 43956 2748
rect 43956 2692 44012 2748
rect 44012 2692 44016 2748
rect 43952 2688 44016 2692
rect 44032 2748 44096 2752
rect 44032 2692 44036 2748
rect 44036 2692 44092 2748
rect 44092 2692 44096 2748
rect 44032 2688 44096 2692
rect 44112 2748 44176 2752
rect 44112 2692 44116 2748
rect 44116 2692 44172 2748
rect 44172 2692 44176 2748
rect 44112 2688 44176 2692
rect 44192 2748 44256 2752
rect 44192 2692 44196 2748
rect 44196 2692 44252 2748
rect 44252 2692 44256 2748
rect 44192 2688 44256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
rect 30972 172 31036 236
<< metal4 >>
rect 1944 8192 2264 11152
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11152
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11152
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11152
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11152
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11152
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11152
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11152
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11152
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11152
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 31944 8192 32264 11152
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 30971 5268 31037 5269
rect 30971 5204 30972 5268
rect 31036 5204 31037 5268
rect 30971 5203 31037 5204
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 30974 237 31034 5203
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 30971 236 31037 237
rect 30971 172 30972 236
rect 31036 172 31037 236
rect 30971 171 31037 172
rect 31944 0 32264 2688
rect 33004 8736 33324 11152
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11152
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11152
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
rect 43944 8192 44264 11152
rect 43944 8128 43952 8192
rect 44016 8128 44032 8192
rect 44096 8128 44112 8192
rect 44176 8128 44192 8192
rect 44256 8128 44264 8192
rect 43944 7104 44264 8128
rect 43944 7040 43952 7104
rect 44016 7040 44032 7104
rect 44096 7040 44112 7104
rect 44176 7040 44192 7104
rect 44256 7040 44264 7104
rect 43944 6016 44264 7040
rect 43944 5952 43952 6016
rect 44016 5952 44032 6016
rect 44096 5952 44112 6016
rect 44176 5952 44192 6016
rect 44256 5952 44264 6016
rect 43944 4928 44264 5952
rect 43944 4864 43952 4928
rect 44016 4864 44032 4928
rect 44096 4864 44112 4928
rect 44176 4864 44192 4928
rect 44256 4864 44264 4928
rect 43944 3840 44264 4864
rect 43944 3776 43952 3840
rect 44016 3776 44032 3840
rect 44096 3776 44112 3840
rect 44176 3776 44192 3840
rect 44256 3776 44264 3840
rect 43944 2752 44264 3776
rect 43944 2688 43952 2752
rect 44016 2688 44032 2752
rect 44096 2688 44112 2752
rect 44176 2688 44192 2752
rect 44256 2688 44264 2752
rect 43944 0 44264 2688
use sky130_fd_sc_hd__clkbuf_2  _000_
timestamp -3599
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _001_
timestamp -3599
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _002_
timestamp -3599
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _003_
timestamp -3599
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _004_
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _005_
timestamp -3599
transform 1 0 42964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _006_
timestamp -3599
transform -1 0 42964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _007_
timestamp -3599
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _008_
timestamp -3599
transform -1 0 42320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _009_
timestamp -3599
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _010_
timestamp -3599
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _011_
timestamp -3599
transform -1 0 43148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _012_
timestamp -3599
transform -1 0 43424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _013_
timestamp -3599
transform 1 0 5888 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _014_
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _015_
timestamp -3599
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _016_
timestamp -3599
transform 1 0 2944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _017_
timestamp -3599
transform -1 0 43608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _018_
timestamp -3599
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _019_
timestamp -3599
transform -1 0 43332 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _020_
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _021_
timestamp -3599
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _022_
timestamp -3599
transform -1 0 42872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _023_
timestamp -3599
transform 1 0 3128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _024_
timestamp -3599
transform -1 0 42688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _025_
timestamp -3599
transform -1 0 43148 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _026_
timestamp -3599
transform -1 0 42780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _027_
timestamp -3599
transform -1 0 42044 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _028_
timestamp -3599
transform -1 0 41584 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _029_
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _030_
timestamp -3599
transform 1 0 2392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp -3599
transform -1 0 42320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _032_
timestamp -3599
transform -1 0 35788 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _033_
timestamp -3599
transform -1 0 35788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp -3599
transform 1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp -3599
transform 1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp -3599
transform 1 0 16560 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _038_
timestamp -3599
transform -1 0 37168 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _039_
timestamp -3599
transform -1 0 37536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _040_
timestamp -3599
transform -1 0 38456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _041_
timestamp -3599
transform -1 0 39652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _042_
timestamp -3599
transform -1 0 40940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _043_
timestamp -3599
transform -1 0 41492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _044_
timestamp -3599
transform -1 0 41492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform 1 0 32384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform 1 0 35788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform 1 0 38088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform 1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 40940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp -3599
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp -3599
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp -3599
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp -3599
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp -3599
transform -1 0 18400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp -3599
transform -1 0 14628 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp -3599
transform -1 0 17664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp -3599
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp -3599
transform 1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp -3599
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp -3599
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp -3599
transform -1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp -3599
transform -1 0 16560 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp -3599
transform -1 0 19872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp -3599
transform -1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp -3599
transform -1 0 22632 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp -3599
transform 1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _069_
timestamp -3599
transform 1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _070_
timestamp -3599
transform 1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp -3599
transform -1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp -3599
transform -1 0 23276 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp -3599
transform -1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp -3599
transform -1 0 26036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform -1 0 27324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp -3599
transform -1 0 28060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform -1 0 28704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp -3599
transform -1 0 29256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp -3599
transform -1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _080_
timestamp -3599
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _081_
timestamp -3599
transform 1 0 16376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _082_
timestamp -3599
transform 1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp -3599
transform -1 0 30636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform -1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _085_
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _086_
timestamp -3599
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp -3599
transform 1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform -1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform -1 0 27232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform -1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp -3599
transform -1 0 29072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp -3599
transform -1 0 31924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _093_
timestamp -3599
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp -3599
transform -1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp -3599
transform -1 0 31924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp -3599
transform 1 0 39284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp -3599
transform -1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform -1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _099_
timestamp -3599
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _100_
timestamp -3599
transform 1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp -3599
transform 1 0 39100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp -3599
transform 1 0 38364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp -3599
transform 1 0 41216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform -1 0 36800 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 43700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 42688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 43148 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 43148 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 43056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform 1 0 42412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 42872 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 42872 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 41584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 42504 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 43884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform 1 0 41860 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 41860 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 41676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 27784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform 1 0 22816 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform 1 0 30176 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform -1 0 28980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform -1 0 41216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform 1 0 28612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform -1 0 35144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 31648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 23368 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 31648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6
timestamp -3599
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp -3599
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12
timestamp -3599
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19
timestamp -3599
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22
timestamp -3599
transform 1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25
timestamp -3599
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp -3599
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35
timestamp -3599
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp -3599
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp -3599
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47
timestamp -3599
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50
timestamp -3599
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60
timestamp -3599
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp -3599
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp -3599
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp -3599
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78
timestamp -3599
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_88
timestamp -3599
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91
timestamp -3599
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp -3599
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp -3599
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100
timestamp -3599
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103
timestamp -3599
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106
timestamp -3599
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_116
timestamp -3599
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp -3599
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_122
timestamp -3599
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp -3599
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_128
timestamp -3599
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_131
timestamp -3599
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_134
timestamp -3599
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_144
timestamp -3599
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_147
timestamp -3599
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_150
timestamp -3599
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_153
timestamp -3599
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp -3599
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_159
timestamp -3599
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_162
timestamp -3599
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_172
timestamp -3599
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_175
timestamp -3599
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_178
timestamp -3599
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp -3599
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_184
timestamp -3599
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp -3599
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_190
timestamp -3599
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp -3599
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_413
timestamp -3599
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_416
timestamp -3599
transform 1 0 39376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp -3599
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_421
timestamp -3599
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_424
timestamp -3599
transform 1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_427
timestamp -3599
transform 1 0 40388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_430
timestamp -3599
transform 1 0 40664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_433
timestamp -3599
transform 1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_436
timestamp -3599
transform 1 0 41216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_439
timestamp -3599
transform 1 0 41492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_442
timestamp -3599
transform 1 0 41768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp -3599
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6
timestamp -3599
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp -3599
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp -3599
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_30
timestamp -3599
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_33
timestamp -3599
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_36
timestamp -3599
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_39
timestamp -3599
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_48
timestamp -3599
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -3599
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_60
timestamp -3599
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_63
timestamp -3599
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_66
timestamp -3599
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp -3599
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_72
timestamp -3599
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_75
timestamp -3599
transform 1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp -3599
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp -3599
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_84
timestamp -3599
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_87
timestamp -3599
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_90
timestamp -3599
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_93
timestamp -3599
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_96
timestamp -3599
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_99
timestamp -3599
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp -3599
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_108
timestamp -3599
transform 1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_116
timestamp -3599
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp -3599
transform 1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_122
timestamp -3599
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp -3599
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_128
timestamp -3599
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_131
timestamp -3599
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_134
timestamp -3599
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_137
timestamp -3599
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_140
timestamp -3599
transform 1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp -3599
transform 1 0 14260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_146
timestamp -3599
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_149
timestamp -3599
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp -3599
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_155
timestamp -3599
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_158
timestamp -3599
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_164
timestamp -3599
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_172
timestamp -3599
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp -3599
transform 1 0 17204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_180
timestamp -3599
transform 1 0 17664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_183
timestamp -3599
transform 1 0 17940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_186
timestamp -3599
transform 1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_189
timestamp -3599
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_192
timestamp -3599
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_195
timestamp -3599
transform 1 0 19044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_202
timestamp -3599
transform 1 0 19688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp -3599
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_211
timestamp -3599
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_214
timestamp -3599
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_217
timestamp -3599
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp -3599
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -3599
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_228
timestamp -3599
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_231
timestamp -3599
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_234
timestamp -3599
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_237
timestamp -3599
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_240
timestamp -3599
transform 1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_243
timestamp -3599
transform 1 0 23460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_246
timestamp -3599
transform 1 0 23736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_249
timestamp -3599
transform 1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_252
timestamp -3599
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_255
timestamp -3599
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_258
timestamp -3599
transform 1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_261
timestamp -3599
transform 1 0 25116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_264
timestamp -3599
transform 1 0 25392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_267
timestamp -3599
transform 1 0 25668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_270
timestamp -3599
transform 1 0 25944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_273
timestamp -3599
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_276
timestamp -3599
transform 1 0 26496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_284
timestamp -3599
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_287
timestamp -3599
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_290
timestamp -3599
transform 1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_293
timestamp -3599
transform 1 0 28060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_296
timestamp -3599
transform 1 0 28336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_302
timestamp -3599
transform 1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_305
timestamp -3599
transform 1 0 29164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_308
timestamp -3599
transform 1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_311
timestamp -3599
transform 1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_314
timestamp -3599
transform 1 0 29992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_324
timestamp -3599
transform 1 0 30912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp -3599
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_340
timestamp -3599
transform 1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_343
timestamp -3599
transform 1 0 32660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_346
timestamp -3599
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_349
timestamp -3599
transform 1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_352
timestamp -3599
transform 1 0 33488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_358
timestamp -3599
transform 1 0 34040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_361
timestamp -3599
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_364
timestamp -3599
transform 1 0 34592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_367
timestamp -3599
transform 1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_370
timestamp -3599
transform 1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_373
timestamp -3599
transform 1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_376
timestamp -3599
transform 1 0 35696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_379
timestamp -3599
transform 1 0 35972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_386
timestamp -3599
transform 1 0 36616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_389
timestamp -3599
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_393
timestamp -3599
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_396
timestamp -3599
transform 1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_399
timestamp -3599
transform 1 0 37812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_402
timestamp -3599
transform 1 0 38088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_405
timestamp -3599
transform 1 0 38364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_408
timestamp -3599
transform 1 0 38640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_411
timestamp -3599
transform 1 0 38916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_414
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_417
timestamp -3599
transform 1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_420
timestamp -3599
transform 1 0 39744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_423
timestamp -3599
transform 1 0 40020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_426
timestamp -3599
transform 1 0 40296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_429
timestamp -3599
transform 1 0 40572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_432
timestamp -3599
transform 1 0 40848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_435
timestamp -3599
transform 1 0 41124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_438
timestamp -3599
transform 1 0 41400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_6
timestamp -3599
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_9
timestamp -3599
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_12
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_18
timestamp -3599
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_21
timestamp -3599
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_24
timestamp -3599
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp -3599
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_35
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_38
timestamp -3599
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp -3599
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_44
timestamp -3599
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_47
timestamp -3599
transform 1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp -3599
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp -3599
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp -3599
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_59
timestamp -3599
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_62
timestamp -3599
transform 1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_65
timestamp -3599
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp -3599
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_71
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_74
timestamp -3599
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_80
timestamp -3599
transform 1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_88
timestamp -3599
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_91
timestamp -3599
transform 1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_94
timestamp -3599
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp -3599
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_100
timestamp -3599
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_103
timestamp -3599
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_106
timestamp -3599
transform 1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp -3599
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_112
timestamp -3599
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_115
timestamp -3599
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_118
timestamp -3599
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_121
timestamp -3599
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_124
timestamp -3599
transform 1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_127
timestamp -3599
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_130
timestamp -3599
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_136
timestamp -3599
transform 1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_144
timestamp -3599
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_147
timestamp -3599
transform 1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp -3599
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_153
timestamp -3599
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_156
timestamp -3599
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_159
timestamp -3599
transform 1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_162
timestamp -3599
transform 1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_165
timestamp -3599
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_171
timestamp -3599
transform 1 0 16836 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_175
timestamp -3599
transform 1 0 17204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_178
timestamp -3599
transform 1 0 17480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_181
timestamp -3599
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_184
timestamp -3599
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp -3599
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_190
timestamp -3599
transform 1 0 18584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp -3599
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_200
timestamp -3599
transform 1 0 19504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_204
timestamp -3599
transform 1 0 19872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_207
timestamp -3599
transform 1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_210
timestamp -3599
transform 1 0 20424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_213
timestamp -3599
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_216
timestamp -3599
transform 1 0 20976 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_219
timestamp -3599
transform 1 0 21252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_222
timestamp -3599
transform 1 0 21528 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_225
timestamp -3599
transform 1 0 21804 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_228
timestamp -3599
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_231
timestamp -3599
transform 1 0 22356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_234
timestamp -3599
transform 1 0 22632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_237
timestamp -3599
transform 1 0 22908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_240
timestamp -3599
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_243
timestamp -3599
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_246
timestamp -3599
transform 1 0 23736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp -3599
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_256
timestamp -3599
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_259
timestamp -3599
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_262
timestamp -3599
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_265
timestamp -3599
transform 1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_268
timestamp -3599
transform 1 0 25760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_271
timestamp -3599
transform 1 0 26036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_274
timestamp -3599
transform 1 0 26312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_277
timestamp -3599
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_280
timestamp -3599
transform 1 0 26864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_283
timestamp -3599
transform 1 0 27140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_286
timestamp -3599
transform 1 0 27416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_293
timestamp -3599
transform 1 0 28060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_300
timestamp -3599
transform 1 0 28704 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp -3599
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_312
timestamp -3599
transform 1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_315
timestamp -3599
transform 1 0 30084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_318
timestamp -3599
transform 1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_321
timestamp -3599
transform 1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_324
timestamp -3599
transform 1 0 30912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_327
timestamp -3599
transform 1 0 31188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_330
timestamp -3599
transform 1 0 31464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_333
timestamp -3599
transform 1 0 31740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_336
timestamp -3599
transform 1 0 32016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_339
timestamp -3599
transform 1 0 32292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_342
timestamp -3599
transform 1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_345
timestamp -3599
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_348
timestamp -3599
transform 1 0 33120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_351
timestamp -3599
transform 1 0 33396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_354
timestamp -3599
transform 1 0 33672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_357
timestamp -3599
transform 1 0 33948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_360
timestamp -3599
transform 1 0 34224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp -3599
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_370
timestamp -3599
transform 1 0 35144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_373
timestamp -3599
transform 1 0 35420 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_377
timestamp -3599
transform 1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_380
timestamp -3599
transform 1 0 36064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_383
timestamp -3599
transform 1 0 36340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_386
timestamp -3599
transform 1 0 36616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_389
timestamp -3599
transform 1 0 36892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_392
timestamp -3599
transform 1 0 37168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_395
timestamp -3599
transform 1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_398
timestamp -3599
transform 1 0 37720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_401
timestamp -3599
transform 1 0 37996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_404
timestamp -3599
transform 1 0 38272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_407
timestamp -3599
transform 1 0 38548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_410
timestamp -3599
transform 1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_413
timestamp -3599
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_416
timestamp -3599
transform 1 0 39376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp -3599
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_421
timestamp -3599
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_424
timestamp -3599
transform 1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_427
timestamp -3599
transform 1 0 40388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_430
timestamp -3599
transform 1 0 40664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_433
timestamp -3599
transform 1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_436
timestamp -3599
transform 1 0 41216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_439
timestamp -3599
transform 1 0 41492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_442
timestamp -3599
transform 1 0 41768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_445
timestamp -3599
transform 1 0 42044 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_448
timestamp -3599
transform 1 0 42320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_451
timestamp -3599
transform 1 0 42596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_457
timestamp -3599
transform 1 0 43148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_460
timestamp -3599
transform 1 0 43424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_463
timestamp -3599
transform 1 0 43700 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_6
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_9
timestamp -3599
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_12
timestamp -3599
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_18
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_21
timestamp -3599
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_24
timestamp -3599
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp -3599
transform 1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_30
timestamp -3599
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_33
timestamp -3599
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_36
timestamp -3599
transform 1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_39
timestamp -3599
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_45
timestamp -3599
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_48
timestamp -3599
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp -3599
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_60
timestamp -3599
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_63
timestamp -3599
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_66
timestamp -3599
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_69
timestamp -3599
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_74
timestamp -3599
transform 1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_77
timestamp -3599
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_80
timestamp -3599
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_83
timestamp -3599
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_86
timestamp -3599
transform 1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_89
timestamp -3599
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_92
timestamp -3599
transform 1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_98
timestamp -3599
transform 1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_101
timestamp -3599
transform 1 0 10396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_104
timestamp -3599
transform 1 0 10672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_107
timestamp -3599
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp -3599
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_116
timestamp -3599
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp -3599
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_122
timestamp -3599
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_125
timestamp -3599
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_128
timestamp -3599
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_131
timestamp -3599
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_134
timestamp -3599
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_137
timestamp -3599
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_140
timestamp -3599
transform 1 0 13984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_143
timestamp -3599
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_146
timestamp -3599
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_149
timestamp -3599
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_152
timestamp -3599
transform 1 0 15088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_155
timestamp -3599
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_158
timestamp -3599
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_164
timestamp -3599
transform 1 0 16192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_172
timestamp -3599
transform 1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_175
timestamp -3599
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_178
timestamp -3599
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp -3599
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp -3599
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_187
timestamp -3599
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_190
timestamp -3599
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_193
timestamp -3599
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_196
timestamp -3599
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_199
timestamp -3599
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_202
timestamp -3599
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_205
timestamp -3599
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_208
timestamp -3599
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_211
timestamp -3599
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_214
timestamp -3599
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp -3599
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp -3599
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_228
timestamp -3599
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_231
timestamp -3599
transform 1 0 22356 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_234
timestamp -3599
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_237
timestamp -3599
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_240
timestamp -3599
transform 1 0 23184 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_243
timestamp -3599
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_246
timestamp -3599
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_249
timestamp -3599
transform 1 0 24012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_252
timestamp -3599
transform 1 0 24288 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_255
timestamp -3599
transform 1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_258
timestamp -3599
transform 1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_261
timestamp -3599
transform 1 0 25116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_264
timestamp -3599
transform 1 0 25392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_267
timestamp -3599
transform 1 0 25668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_270
timestamp -3599
transform 1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_273
timestamp -3599
transform 1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_276
timestamp -3599
transform 1 0 26496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_281
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_285
timestamp -3599
transform 1 0 27324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_288
timestamp -3599
transform 1 0 27600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_291
timestamp -3599
transform 1 0 27876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_294
timestamp -3599
transform 1 0 28152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_297
timestamp -3599
transform 1 0 28428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_300
timestamp -3599
transform 1 0 28704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_303
timestamp -3599
transform 1 0 28980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_306
timestamp -3599
transform 1 0 29256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_309
timestamp -3599
transform 1 0 29532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_312
timestamp -3599
transform 1 0 29808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_315
timestamp -3599
transform 1 0 30084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_318
timestamp -3599
transform 1 0 30360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_321
timestamp -3599
transform 1 0 30636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_324
timestamp -3599
transform 1 0 30912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_327
timestamp -3599
transform 1 0 31188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_330
timestamp -3599
transform 1 0 31464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp -3599
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_340
timestamp -3599
transform 1 0 32384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_343
timestamp -3599
transform 1 0 32660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_346
timestamp -3599
transform 1 0 32936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_349
timestamp -3599
transform 1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_352
timestamp -3599
transform 1 0 33488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_355
timestamp -3599
transform 1 0 33764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_358
timestamp -3599
transform 1 0 34040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_361
timestamp -3599
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_364
timestamp -3599
transform 1 0 34592 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_367
timestamp -3599
transform 1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_370
timestamp -3599
transform 1 0 35144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_373
timestamp -3599
transform 1 0 35420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_376
timestamp -3599
transform 1 0 35696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_379
timestamp -3599
transform 1 0 35972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_382
timestamp -3599
transform 1 0 36248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_388
timestamp -3599
transform 1 0 36800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_393
timestamp -3599
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_396
timestamp -3599
transform 1 0 37536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_399
timestamp -3599
transform 1 0 37812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_402
timestamp -3599
transform 1 0 38088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_408
timestamp -3599
transform 1 0 38640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_411
timestamp -3599
transform 1 0 38916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_414
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_417
timestamp -3599
transform 1 0 39468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_420
timestamp -3599
transform 1 0 39744 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_423
timestamp -3599
transform 1 0 40020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_426
timestamp -3599
transform 1 0 40296 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_429
timestamp -3599
transform 1 0 40572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_432
timestamp -3599
transform 1 0 40848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_435
timestamp -3599
transform 1 0 41124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_438
timestamp -3599
transform 1 0 41400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_441
timestamp -3599
transform 1 0 41676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_444
timestamp -3599
transform 1 0 41952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp -3599
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_449
timestamp -3599
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_452
timestamp -3599
transform 1 0 42688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_460
timestamp -3599
transform 1 0 43424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_463
timestamp -3599
transform 1 0 43700 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_6
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp -3599
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_14
timestamp -3599
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_17
timestamp -3599
transform 1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_20
timestamp -3599
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_23
timestamp -3599
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp -3599
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp -3599
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_35
timestamp -3599
transform 1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp -3599
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_44
timestamp -3599
transform 1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_47
timestamp -3599
transform 1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_50
timestamp -3599
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp -3599
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_59
timestamp -3599
transform 1 0 6532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp -3599
transform 1 0 6900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_68
timestamp -3599
transform 1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_71
timestamp -3599
transform 1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_74
timestamp -3599
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_80
timestamp -3599
transform 1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_88
timestamp -3599
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_91
timestamp -3599
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_94
timestamp -3599
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_100
timestamp -3599
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_103
timestamp -3599
transform 1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp -3599
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_112
timestamp -3599
transform 1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_115
timestamp -3599
transform 1 0 11684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_120
timestamp -3599
transform 1 0 12144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_123
timestamp -3599
transform 1 0 12420 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_126
timestamp -3599
transform 1 0 12696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_130
timestamp -3599
transform 1 0 13064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_133
timestamp -3599
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_136
timestamp -3599
transform 1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_144
timestamp -3599
transform 1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_147
timestamp -3599
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp -3599
transform 1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_153
timestamp -3599
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp -3599
transform 1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_159
timestamp -3599
transform 1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_162
timestamp -3599
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_165
timestamp -3599
transform 1 0 16284 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_169
timestamp -3599
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_172
timestamp -3599
transform 1 0 16928 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_175
timestamp -3599
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_178
timestamp -3599
transform 1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_181
timestamp -3599
transform 1 0 17756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_184
timestamp -3599
transform 1 0 18032 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_187
timestamp -3599
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_190
timestamp -3599
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp -3599
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_200
timestamp -3599
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_203
timestamp -3599
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_206
timestamp -3599
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp -3599
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_212
timestamp -3599
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_215
timestamp -3599
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_218
timestamp -3599
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp -3599
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_224
timestamp -3599
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_227
timestamp -3599
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_230
timestamp -3599
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_233
timestamp -3599
transform 1 0 22540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_236
timestamp -3599
transform 1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_239
timestamp -3599
transform 1 0 23092 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_245
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_248
timestamp -3599
transform 1 0 23920 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_256
timestamp -3599
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_259
timestamp -3599
transform 1 0 24932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_262
timestamp -3599
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_265
timestamp -3599
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_268
timestamp -3599
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_271
timestamp -3599
transform 1 0 26036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_274
timestamp -3599
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_277
timestamp -3599
transform 1 0 26588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_280
timestamp -3599
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_283
timestamp -3599
transform 1 0 27140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_286
timestamp -3599
transform 1 0 27416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_289
timestamp -3599
transform 1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_292
timestamp -3599
transform 1 0 27968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_295
timestamp -3599
transform 1 0 28244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_298
timestamp -3599
transform 1 0 28520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_301
timestamp -3599
transform 1 0 28796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_304
timestamp -3599
transform 1 0 29072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_312
timestamp -3599
transform 1 0 29808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_315
timestamp -3599
transform 1 0 30084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_318
timestamp -3599
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_324
timestamp -3599
transform 1 0 30912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_327
timestamp -3599
transform 1 0 31188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_330
timestamp -3599
transform 1 0 31464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp -3599
transform 1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_336
timestamp -3599
transform 1 0 32016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_339
timestamp -3599
transform 1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_342
timestamp -3599
transform 1 0 32568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_345
timestamp -3599
transform 1 0 32844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_348
timestamp -3599
transform 1 0 33120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_351
timestamp -3599
transform 1 0 33396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_354
timestamp -3599
transform 1 0 33672 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_357
timestamp -3599
transform 1 0 33948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_360
timestamp -3599
transform 1 0 34224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp -3599
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_365
timestamp -3599
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_368
timestamp -3599
transform 1 0 34960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_371
timestamp -3599
transform 1 0 35236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_374
timestamp -3599
transform 1 0 35512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_377
timestamp -3599
transform 1 0 35788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_380
timestamp -3599
transform 1 0 36064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_383
timestamp -3599
transform 1 0 36340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_386
timestamp -3599
transform 1 0 36616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_389
timestamp -3599
transform 1 0 36892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_392
timestamp -3599
transform 1 0 37168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_395
timestamp -3599
transform 1 0 37444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_398
timestamp -3599
transform 1 0 37720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_401
timestamp -3599
transform 1 0 37996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_404
timestamp -3599
transform 1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_407
timestamp -3599
transform 1 0 38548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_410
timestamp -3599
transform 1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_416
timestamp -3599
transform 1 0 39376 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp -3599
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_421
timestamp -3599
transform 1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_424
timestamp -3599
transform 1 0 40112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_427
timestamp -3599
transform 1 0 40388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_430
timestamp -3599
transform 1 0 40664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_433
timestamp -3599
transform 1 0 40940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_439
timestamp -3599
transform 1 0 41492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_442
timestamp -3599
transform 1 0 41768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_445
timestamp -3599
transform 1 0 42044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_448
timestamp -3599
transform 1 0 42320 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_454
timestamp -3599
transform 1 0 42872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_457
timestamp -3599
transform 1 0 43148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_460
timestamp -3599
transform 1 0 43424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_6
timestamp -3599
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_9
timestamp -3599
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp -3599
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_18
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp -3599
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_33
timestamp -3599
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_36
timestamp -3599
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_42
timestamp -3599
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_45
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_48
timestamp -3599
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_60
timestamp -3599
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_63
timestamp -3599
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_66
timestamp -3599
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_72
timestamp -3599
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp -3599
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_84
timestamp -3599
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_87
timestamp -3599
transform 1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_90
timestamp -3599
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp -3599
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_96
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_99
timestamp -3599
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_102
timestamp -3599
transform 1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_108
timestamp -3599
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_116
timestamp -3599
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp -3599
transform 1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_122
timestamp -3599
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp -3599
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_128
timestamp -3599
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_131
timestamp -3599
transform 1 0 13156 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_134
timestamp -3599
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_137
timestamp -3599
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_140
timestamp -3599
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp -3599
transform 1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_146
timestamp -3599
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp -3599
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_152
timestamp -3599
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_155
timestamp -3599
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_158
timestamp -3599
transform 1 0 15640 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp -3599
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_172
timestamp -3599
transform 1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_175
timestamp -3599
transform 1 0 17204 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_178
timestamp -3599
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_181
timestamp -3599
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp -3599
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_187
timestamp -3599
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_190
timestamp -3599
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_193
timestamp -3599
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_196
timestamp -3599
transform 1 0 19136 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_199
timestamp -3599
transform 1 0 19412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_202
timestamp -3599
transform 1 0 19688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_205
timestamp -3599
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_208
timestamp -3599
transform 1 0 20240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_213
timestamp -3599
transform 1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_216
timestamp -3599
transform 1 0 20976 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_219
timestamp -3599
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp -3599
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_228
timestamp -3599
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_231
timestamp -3599
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_234
timestamp -3599
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_237
timestamp -3599
transform 1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_240
timestamp -3599
transform 1 0 23184 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_243
timestamp -3599
transform 1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_246
timestamp -3599
transform 1 0 23736 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_249
timestamp -3599
transform 1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_252
timestamp -3599
transform 1 0 24288 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_255
timestamp -3599
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_258
timestamp -3599
transform 1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_261
timestamp -3599
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_264
timestamp -3599
transform 1 0 25392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_267
timestamp -3599
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_270
timestamp -3599
transform 1 0 25944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_276
timestamp -3599
transform 1 0 26496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_284
timestamp -3599
transform 1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_287
timestamp -3599
transform 1 0 27508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_290
timestamp -3599
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_293
timestamp -3599
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_296
timestamp -3599
transform 1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_299
timestamp -3599
transform 1 0 28612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_302
timestamp -3599
transform 1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_305
timestamp -3599
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_308
timestamp -3599
transform 1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_311
timestamp -3599
transform 1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_314
timestamp -3599
transform 1 0 29992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_317
timestamp -3599
transform 1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_320
timestamp -3599
transform 1 0 30544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_323
timestamp -3599
transform 1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_326
timestamp -3599
transform 1 0 31096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_329
timestamp -3599
transform 1 0 31372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp -3599
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_337
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_340
timestamp -3599
transform 1 0 32384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_343
timestamp -3599
transform 1 0 32660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_346
timestamp -3599
transform 1 0 32936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_349
timestamp -3599
transform 1 0 33212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_352
timestamp -3599
transform 1 0 33488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_355
timestamp -3599
transform 1 0 33764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_358
timestamp -3599
transform 1 0 34040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_361
timestamp -3599
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_364
timestamp -3599
transform 1 0 34592 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_367
timestamp -3599
transform 1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_370
timestamp -3599
transform 1 0 35144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_373
timestamp -3599
transform 1 0 35420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_376
timestamp -3599
transform 1 0 35696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_379
timestamp -3599
transform 1 0 35972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_382
timestamp -3599
transform 1 0 36248 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_388
timestamp -3599
transform 1 0 36800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_393
timestamp -3599
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_396
timestamp -3599
transform 1 0 37536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_399
timestamp -3599
transform 1 0 37812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_402
timestamp -3599
transform 1 0 38088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_405
timestamp -3599
transform 1 0 38364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_408
timestamp -3599
transform 1 0 38640 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_411
timestamp -3599
transform 1 0 38916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_414
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_417
timestamp -3599
transform 1 0 39468 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_420
timestamp -3599
transform 1 0 39744 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_423
timestamp -3599
transform 1 0 40020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_426
timestamp -3599
transform 1 0 40296 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_429
timestamp -3599
transform 1 0 40572 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_432
timestamp -3599
transform 1 0 40848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_435
timestamp -3599
transform 1 0 41124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_438
timestamp -3599
transform 1 0 41400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_441
timestamp -3599
transform 1 0 41676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_444
timestamp -3599
transform 1 0 41952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp -3599
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_459
timestamp -3599
transform 1 0 43332 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_462
timestamp -3599
transform 1 0 43608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_6
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_13
timestamp -3599
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_16
timestamp -3599
transform 1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_19
timestamp -3599
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_22
timestamp -3599
transform 1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp -3599
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_38
timestamp -3599
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_44
timestamp -3599
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_47
timestamp -3599
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_50
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp -3599
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp -3599
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_59
timestamp -3599
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_62
timestamp -3599
transform 1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_65
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_68
timestamp -3599
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_71
timestamp -3599
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_74
timestamp -3599
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_77
timestamp -3599
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_80
timestamp -3599
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_88
timestamp -3599
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_91
timestamp -3599
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_94
timestamp -3599
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_97
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_100
timestamp -3599
transform 1 0 10304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_103
timestamp -3599
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_106
timestamp -3599
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_109
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_112
timestamp -3599
transform 1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_115
timestamp -3599
transform 1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_118
timestamp -3599
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp -3599
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_124
timestamp -3599
transform 1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_127
timestamp -3599
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_130
timestamp -3599
transform 1 0 13064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_136
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_144
timestamp -3599
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_147
timestamp -3599
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp -3599
transform 1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_153
timestamp -3599
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp -3599
transform 1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_159
timestamp -3599
transform 1 0 15732 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_162
timestamp -3599
transform 1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_171
timestamp -3599
transform 1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_174
timestamp -3599
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_177
timestamp -3599
transform 1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_180
timestamp -3599
transform 1 0 17664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_183
timestamp -3599
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_186
timestamp -3599
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_189
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_192
timestamp -3599
transform 1 0 18768 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_200
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_203
timestamp -3599
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_206
timestamp -3599
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_212
timestamp -3599
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp -3599
transform 1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_218
timestamp -3599
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_221
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_224
timestamp -3599
transform 1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_227
timestamp -3599
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_230
timestamp -3599
transform 1 0 22264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_234
timestamp -3599
transform 1 0 22632 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_237
timestamp -3599
transform 1 0 22908 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_240
timestamp -3599
transform 1 0 23184 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_243
timestamp -3599
transform 1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_246
timestamp -3599
transform 1 0 23736 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp -3599
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_256
timestamp -3599
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_259
timestamp -3599
transform 1 0 24932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_262
timestamp -3599
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_268
timestamp -3599
transform 1 0 25760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_271
timestamp -3599
transform 1 0 26036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_274
timestamp -3599
transform 1 0 26312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_277
timestamp -3599
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_280
timestamp -3599
transform 1 0 26864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_284
timestamp -3599
transform 1 0 27232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_287
timestamp -3599
transform 1 0 27508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_290
timestamp -3599
transform 1 0 27784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_293
timestamp -3599
transform 1 0 28060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_296
timestamp -3599
transform 1 0 28336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_299
timestamp -3599
transform 1 0 28612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_302
timestamp -3599
transform 1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_305
timestamp -3599
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_312
timestamp -3599
transform 1 0 29808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_315
timestamp -3599
transform 1 0 30084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_318
timestamp -3599
transform 1 0 30360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_321
timestamp -3599
transform 1 0 30636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_324
timestamp -3599
transform 1 0 30912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_327
timestamp -3599
transform 1 0 31188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_335
timestamp -3599
transform 1 0 31924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_338
timestamp -3599
transform 1 0 32200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_341
timestamp -3599
transform 1 0 32476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_344
timestamp -3599
transform 1 0 32752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_347
timestamp -3599
transform 1 0 33028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_350
timestamp -3599
transform 1 0 33304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_353
timestamp -3599
transform 1 0 33580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_356
timestamp -3599
transform 1 0 33856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_359
timestamp -3599
transform 1 0 34132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp -3599
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_365
timestamp -3599
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_368
timestamp -3599
transform 1 0 34960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_371
timestamp -3599
transform 1 0 35236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_374
timestamp -3599
transform 1 0 35512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_377
timestamp -3599
transform 1 0 35788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_380
timestamp -3599
transform 1 0 36064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_383
timestamp -3599
transform 1 0 36340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_386
timestamp -3599
transform 1 0 36616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_389
timestamp -3599
transform 1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_392
timestamp -3599
transform 1 0 37168 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_395
timestamp -3599
transform 1 0 37444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_398
timestamp -3599
transform 1 0 37720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_401
timestamp -3599
transform 1 0 37996 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_404
timestamp -3599
transform 1 0 38272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_407
timestamp -3599
transform 1 0 38548 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_410
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_413
timestamp -3599
transform 1 0 39100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_416
timestamp -3599
transform 1 0 39376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp -3599
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_421
timestamp -3599
transform 1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_424
timestamp -3599
transform 1 0 40112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_427
timestamp -3599
transform 1 0 40388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_430
timestamp -3599
transform 1 0 40664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_433
timestamp -3599
transform 1 0 40940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_436
timestamp -3599
transform 1 0 41216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_439
timestamp -3599
transform 1 0 41492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_442
timestamp -3599
transform 1 0 41768 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_445
timestamp -3599
transform 1 0 42044 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_448
timestamp -3599
transform 1 0 42320 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_451
timestamp -3599
transform 1 0 42596 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_454
timestamp -3599
transform 1 0 42872 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_462
timestamp -3599
transform 1 0 43608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_6
timestamp -3599
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_9
timestamp -3599
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_12
timestamp -3599
transform 1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_18
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_21
timestamp -3599
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_30
timestamp -3599
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_33
timestamp -3599
transform 1 0 4140 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_38
timestamp -3599
transform 1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_41
timestamp -3599
transform 1 0 4876 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_46
timestamp -3599
transform 1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_49
timestamp -3599
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_52
timestamp -3599
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_60
timestamp -3599
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_63
timestamp -3599
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_66
timestamp -3599
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp -3599
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_75
timestamp -3599
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_78
timestamp -3599
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_81
timestamp -3599
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_84
timestamp -3599
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_87
timestamp -3599
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_90
timestamp -3599
transform 1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_93
timestamp -3599
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_96
timestamp -3599
transform 1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_99
timestamp -3599
transform 1 0 10212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_102
timestamp -3599
transform 1 0 10488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_105
timestamp -3599
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_108
timestamp -3599
transform 1 0 11040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_116
timestamp -3599
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp -3599
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp -3599
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_125
timestamp -3599
transform 1 0 12604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_128
timestamp -3599
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_131
timestamp -3599
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_134
timestamp -3599
transform 1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_137
timestamp -3599
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_140
timestamp -3599
transform 1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_143
timestamp -3599
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_146
timestamp -3599
transform 1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_149
timestamp -3599
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_152
timestamp -3599
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_155
timestamp -3599
transform 1 0 15364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_158
timestamp -3599
transform 1 0 15640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_164
timestamp -3599
transform 1 0 16192 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_172
timestamp -3599
transform 1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_175
timestamp -3599
transform 1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_178
timestamp -3599
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp -3599
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp -3599
transform 1 0 18032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_188
timestamp -3599
transform 1 0 18400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_191
timestamp -3599
transform 1 0 18676 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_194
timestamp -3599
transform 1 0 18952 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_197
timestamp -3599
transform 1 0 19228 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_200
timestamp -3599
transform 1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_203
timestamp -3599
transform 1 0 19780 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_206
timestamp -3599
transform 1 0 20056 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_209
timestamp -3599
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_212
timestamp -3599
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_215
timestamp -3599
transform 1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_218
timestamp -3599
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp -3599
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_228
timestamp -3599
transform 1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_231
timestamp -3599
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_234
timestamp -3599
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_241
timestamp -3599
transform 1 0 23276 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_244
timestamp -3599
transform 1 0 23552 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_247
timestamp -3599
transform 1 0 23828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_250
timestamp -3599
transform 1 0 24104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_253
timestamp -3599
transform 1 0 24380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_256
timestamp -3599
transform 1 0 24656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_259
timestamp -3599
transform 1 0 24932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_262
timestamp -3599
transform 1 0 25208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_265
timestamp -3599
transform 1 0 25484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_271
timestamp -3599
transform 1 0 26036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_274
timestamp -3599
transform 1 0 26312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp -3599
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_284
timestamp -3599
transform 1 0 27232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_287
timestamp -3599
transform 1 0 27508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_290
timestamp -3599
transform 1 0 27784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_296
timestamp -3599
transform 1 0 28336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_299
timestamp -3599
transform 1 0 28612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_302
timestamp -3599
transform 1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_305
timestamp -3599
transform 1 0 29164 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_308
timestamp -3599
transform 1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_311
timestamp -3599
transform 1 0 29716 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_314
timestamp -3599
transform 1 0 29992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_317
timestamp -3599
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_320
timestamp -3599
transform 1 0 30544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_323
timestamp -3599
transform 1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_326
timestamp -3599
transform 1 0 31096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_332
timestamp -3599
transform 1 0 31648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_340
timestamp -3599
transform 1 0 32384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_343
timestamp -3599
transform 1 0 32660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_346
timestamp -3599
transform 1 0 32936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_349
timestamp -3599
transform 1 0 33212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_352
timestamp -3599
transform 1 0 33488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_355
timestamp -3599
transform 1 0 33764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_358
timestamp -3599
transform 1 0 34040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_361
timestamp -3599
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_364
timestamp -3599
transform 1 0 34592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_367
timestamp -3599
transform 1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_370
timestamp -3599
transform 1 0 35144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_373
timestamp -3599
transform 1 0 35420 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_376
timestamp -3599
transform 1 0 35696 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_379
timestamp -3599
transform 1 0 35972 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_382
timestamp -3599
transform 1 0 36248 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_385
timestamp -3599
transform 1 0 36524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_388
timestamp -3599
transform 1 0 36800 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_396
timestamp -3599
transform 1 0 37536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_399
timestamp -3599
transform 1 0 37812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_402
timestamp -3599
transform 1 0 38088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_406
timestamp -3599
transform 1 0 38456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_409
timestamp -3599
transform 1 0 38732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_412
timestamp -3599
transform 1 0 39008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_415
timestamp -3599
transform 1 0 39284 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_419
timestamp -3599
transform 1 0 39652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_422
timestamp -3599
transform 1 0 39928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_425
timestamp -3599
transform 1 0 40204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_428
timestamp -3599
transform 1 0 40480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_433
timestamp -3599
transform 1 0 40940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_436
timestamp -3599
transform 1 0 41216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_439
timestamp -3599
transform 1 0 41492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_442
timestamp -3599
transform 1 0 41768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_445
timestamp -3599
transform 1 0 42044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_449
timestamp -3599
transform 1 0 42412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_457
timestamp -3599
transform 1 0 43148 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_460
timestamp -3599
transform 1 0 43424 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_463
timestamp -3599
transform 1 0 43700 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_6
timestamp -3599
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_9
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_12
timestamp -3599
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_19
timestamp -3599
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_22
timestamp -3599
transform 1 0 3128 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp -3599
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp -3599
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_35
timestamp -3599
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp -3599
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp -3599
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_47
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_50
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_56
timestamp -3599
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_59
timestamp -3599
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_68
timestamp -3599
transform 1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_71
timestamp -3599
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_74
timestamp -3599
transform 1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_77
timestamp -3599
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_80
timestamp -3599
transform 1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_88
timestamp -3599
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_91
timestamp -3599
transform 1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_94
timestamp -3599
transform 1 0 9752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp -3599
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_100
timestamp -3599
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_103
timestamp -3599
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_106
timestamp -3599
transform 1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_109
timestamp -3599
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_112
timestamp -3599
transform 1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_115
timestamp -3599
transform 1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_118
timestamp -3599
transform 1 0 11960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_121
timestamp -3599
transform 1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_124
timestamp -3599
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_127
timestamp -3599
transform 1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_130
timestamp -3599
transform 1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_133
timestamp -3599
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_136
timestamp -3599
transform 1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_144
timestamp -3599
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_147
timestamp -3599
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp -3599
transform 1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp -3599
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_159
timestamp -3599
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_162
timestamp -3599
transform 1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp -3599
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp -3599
transform 1 0 16560 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_171
timestamp -3599
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_174
timestamp -3599
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_180
timestamp -3599
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_183
timestamp -3599
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_186
timestamp -3599
transform 1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_192
timestamp -3599
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_200
timestamp -3599
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_203
timestamp -3599
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_206
timestamp -3599
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp -3599
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_212
timestamp -3599
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_215
timestamp -3599
transform 1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_218
timestamp -3599
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_221
timestamp -3599
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_224
timestamp -3599
transform 1 0 21712 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_227
timestamp -3599
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_230
timestamp -3599
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_233
timestamp -3599
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_236
timestamp -3599
transform 1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_239
timestamp -3599
transform 1 0 23092 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_242
timestamp -3599
transform 1 0 23368 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_245
timestamp -3599
transform 1 0 23644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_248
timestamp -3599
transform 1 0 23920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_256
timestamp -3599
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_259
timestamp -3599
transform 1 0 24932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_262
timestamp -3599
transform 1 0 25208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_265
timestamp -3599
transform 1 0 25484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_268
timestamp -3599
transform 1 0 25760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_271
timestamp -3599
transform 1 0 26036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_274
timestamp -3599
transform 1 0 26312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_277
timestamp -3599
transform 1 0 26588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_280
timestamp -3599
transform 1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_283
timestamp -3599
transform 1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_286
timestamp -3599
transform 1 0 27416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_289
timestamp -3599
transform 1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_292
timestamp -3599
transform 1 0 27968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_295
timestamp -3599
transform 1 0 28244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_298
timestamp -3599
transform 1 0 28520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_301
timestamp -3599
transform 1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_304
timestamp -3599
transform 1 0 29072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_312
timestamp -3599
transform 1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_315
timestamp -3599
transform 1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_318
timestamp -3599
transform 1 0 30360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_321
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_324
timestamp -3599
transform 1 0 30912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_327
timestamp -3599
transform 1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_335
timestamp -3599
transform 1 0 31924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_338
timestamp -3599
transform 1 0 32200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_341
timestamp -3599
transform 1 0 32476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_344
timestamp -3599
transform 1 0 32752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_347
timestamp -3599
transform 1 0 33028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_350
timestamp -3599
transform 1 0 33304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_353
timestamp -3599
transform 1 0 33580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_356
timestamp -3599
transform 1 0 33856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_359
timestamp -3599
transform 1 0 34132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp -3599
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_365
timestamp -3599
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_368
timestamp -3599
transform 1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_371
timestamp -3599
transform 1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_374
timestamp -3599
transform 1 0 35512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_377
timestamp -3599
transform 1 0 35788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_380
timestamp -3599
transform 1 0 36064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_383
timestamp -3599
transform 1 0 36340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_386
timestamp -3599
transform 1 0 36616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_389
timestamp -3599
transform 1 0 36892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_392
timestamp -3599
transform 1 0 37168 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_395
timestamp -3599
transform 1 0 37444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_398
timestamp -3599
transform 1 0 37720 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_401
timestamp -3599
transform 1 0 37996 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_404
timestamp -3599
transform 1 0 38272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_407
timestamp -3599
transform 1 0 38548 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_410
timestamp -3599
transform 1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_413
timestamp -3599
transform 1 0 39100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_416
timestamp -3599
transform 1 0 39376 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp -3599
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_421
timestamp -3599
transform 1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_424
timestamp -3599
transform 1 0 40112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_427
timestamp -3599
transform 1 0 40388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_430
timestamp -3599
transform 1 0 40664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_433
timestamp -3599
transform 1 0 40940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_439
timestamp -3599
transform 1 0 41492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_442
timestamp -3599
transform 1 0 41768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_445
timestamp -3599
transform 1 0 42044 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_448
timestamp -3599
transform 1 0 42320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_451
timestamp -3599
transform 1 0 42596 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_454
timestamp -3599
transform 1 0 42872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_457
timestamp -3599
transform 1 0 43148 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_460
timestamp -3599
transform 1 0 43424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_463
timestamp -3599
transform 1 0 43700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6
timestamp -3599
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_9
timestamp -3599
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_12
timestamp -3599
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp -3599
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_18
timestamp -3599
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_21
timestamp -3599
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_24
timestamp -3599
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp -3599
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_30
timestamp -3599
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_33
timestamp -3599
transform 1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_36
timestamp -3599
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_39
timestamp -3599
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_42
timestamp -3599
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_45
timestamp -3599
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_48
timestamp -3599
transform 1 0 5520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_51
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp -3599
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_60
timestamp -3599
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_63
timestamp -3599
transform 1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_66
timestamp -3599
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_72
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_75
timestamp -3599
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_78
timestamp -3599
transform 1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp -3599
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_84
timestamp -3599
transform 1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_87
timestamp -3599
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_90
timestamp -3599
transform 1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_93
timestamp -3599
transform 1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_96
timestamp -3599
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_99
timestamp -3599
transform 1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_102
timestamp -3599
transform 1 0 10488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_108
timestamp -3599
transform 1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_116
timestamp -3599
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_122
timestamp -3599
transform 1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_125
timestamp -3599
transform 1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_128
timestamp -3599
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_131
timestamp -3599
transform 1 0 13156 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_134
timestamp -3599
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp -3599
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_140
timestamp -3599
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_143
timestamp -3599
transform 1 0 14260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_147
timestamp -3599
transform 1 0 14628 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_150
timestamp -3599
transform 1 0 14904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_153
timestamp -3599
transform 1 0 15180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_156
timestamp -3599
transform 1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_159
timestamp -3599
transform 1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_162
timestamp -3599
transform 1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp -3599
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_172
timestamp -3599
transform 1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_175
timestamp -3599
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_178
timestamp -3599
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_181
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_184
timestamp -3599
transform 1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_187
timestamp -3599
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_190
timestamp -3599
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp -3599
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_196
timestamp -3599
transform 1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_199
timestamp -3599
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_202
timestamp -3599
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_205
timestamp -3599
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_208
timestamp -3599
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_211
timestamp -3599
transform 1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_214
timestamp -3599
transform 1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_217
timestamp -3599
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_220
timestamp -3599
transform 1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_228
timestamp -3599
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_231
timestamp -3599
transform 1 0 22356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_234
timestamp -3599
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_237
timestamp -3599
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_240
timestamp -3599
transform 1 0 23184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_243
timestamp -3599
transform 1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_246
timestamp -3599
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_249
timestamp -3599
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_252
timestamp -3599
transform 1 0 24288 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_255
timestamp -3599
transform 1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_258
timestamp -3599
transform 1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_261
timestamp -3599
transform 1 0 25116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_264
timestamp -3599
transform 1 0 25392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_267
timestamp -3599
transform 1 0 25668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_270
timestamp -3599
transform 1 0 25944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_275
timestamp -3599
transform 1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp -3599
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_284
timestamp -3599
transform 1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_287
timestamp -3599
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_290
timestamp -3599
transform 1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_293
timestamp -3599
transform 1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_296
timestamp -3599
transform 1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_304
timestamp -3599
transform 1 0 29072 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_307
timestamp -3599
transform 1 0 29348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_310
timestamp -3599
transform 1 0 29624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_313
timestamp -3599
transform 1 0 29900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_316
timestamp -3599
transform 1 0 30176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_319
timestamp -3599
transform 1 0 30452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_322
timestamp -3599
transform 1 0 30728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_325
timestamp -3599
transform 1 0 31004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_328
timestamp -3599
transform 1 0 31280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_331
timestamp -3599
transform 1 0 31556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp -3599
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_340
timestamp -3599
transform 1 0 32384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_343
timestamp -3599
transform 1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_346
timestamp -3599
transform 1 0 32936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_349
timestamp -3599
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_352
timestamp -3599
transform 1 0 33488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_355
timestamp -3599
transform 1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_358
timestamp -3599
transform 1 0 34040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp -3599
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_364
timestamp -3599
transform 1 0 34592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_367
timestamp -3599
transform 1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_370
timestamp -3599
transform 1 0 35144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_377
timestamp -3599
transform 1 0 35788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_380
timestamp -3599
transform 1 0 36064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_383
timestamp -3599
transform 1 0 36340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_386
timestamp -3599
transform 1 0 36616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp -3599
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_396
timestamp -3599
transform 1 0 37536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_399
timestamp -3599
transform 1 0 37812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_402
timestamp -3599
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_405
timestamp -3599
transform 1 0 38364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_408
timestamp -3599
transform 1 0 38640 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_411
timestamp -3599
transform 1 0 38916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_414
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_417
timestamp -3599
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_420
timestamp -3599
transform 1 0 39744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_423
timestamp -3599
transform 1 0 40020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_426
timestamp -3599
transform 1 0 40296 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_429
timestamp -3599
transform 1 0 40572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_432
timestamp -3599
transform 1 0 40848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_435
timestamp -3599
transform 1 0 41124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_439
timestamp -3599
transform 1 0 41492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_442
timestamp -3599
transform 1 0 41768 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp -3599
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_449
timestamp -3599
transform 1 0 42412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_452
timestamp -3599
transform 1 0 42688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_455
timestamp -3599
transform 1 0 42964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_458
timestamp -3599
transform 1 0 43240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_461
timestamp -3599
transform 1 0 43516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_6
timestamp -3599
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_9
timestamp -3599
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_12
timestamp -3599
transform 1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp -3599
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp -3599
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_35
timestamp -3599
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_38
timestamp -3599
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_44
timestamp -3599
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_47
timestamp -3599
transform 1 0 5428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_50
timestamp -3599
transform 1 0 5704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_57
timestamp -3599
transform 1 0 6348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_60
timestamp -3599
transform 1 0 6624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_63
timestamp -3599
transform 1 0 6900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_66
timestamp -3599
transform 1 0 7176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_69
timestamp -3599
transform 1 0 7452 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_72
timestamp -3599
transform 1 0 7728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_75
timestamp -3599
transform 1 0 8004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_78
timestamp -3599
transform 1 0 8280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp -3599
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_88
timestamp -3599
transform 1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_91
timestamp -3599
transform 1 0 9476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_99
timestamp -3599
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_102
timestamp -3599
transform 1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp -3599
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_108
timestamp -3599
transform 1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_111
timestamp -3599
transform 1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_114
timestamp -3599
transform 1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_117
timestamp -3599
transform 1 0 11868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_124
timestamp -3599
transform 1 0 12512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_127
timestamp -3599
transform 1 0 12788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_130
timestamp -3599
transform 1 0 13064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_133
timestamp -3599
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_136
timestamp -3599
transform 1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_144
timestamp -3599
transform 1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_147
timestamp -3599
transform 1 0 14628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp -3599
transform 1 0 14904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_153
timestamp -3599
transform 1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_156
timestamp -3599
transform 1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_159
timestamp -3599
transform 1 0 15732 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_162
timestamp -3599
transform 1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp -3599
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_168
timestamp -3599
transform 1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_171
timestamp -3599
transform 1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_174
timestamp -3599
transform 1 0 17112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_177
timestamp -3599
transform 1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_180
timestamp -3599
transform 1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_183
timestamp -3599
transform 1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_186
timestamp -3599
transform 1 0 18216 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_192
timestamp -3599
transform 1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_200
timestamp -3599
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_203
timestamp -3599
transform 1 0 19780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_206
timestamp -3599
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp -3599
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_212
timestamp -3599
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp -3599
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_218
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_221
timestamp -3599
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_224
timestamp -3599
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_227
timestamp -3599
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp -3599
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_233
timestamp -3599
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_236
timestamp -3599
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_239
timestamp -3599
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_242
timestamp -3599
transform 1 0 23368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_247
timestamp -3599
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp -3599
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_256
timestamp -3599
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_259
timestamp -3599
transform 1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_262
timestamp -3599
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_265
timestamp -3599
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_268
timestamp -3599
transform 1 0 25760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_271
timestamp -3599
transform 1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_274
timestamp -3599
transform 1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_277
timestamp -3599
transform 1 0 26588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_280
timestamp -3599
transform 1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_283
timestamp -3599
transform 1 0 27140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_286
timestamp -3599
transform 1 0 27416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_289
timestamp -3599
transform 1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_292
timestamp -3599
transform 1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_295
timestamp -3599
transform 1 0 28244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_298
timestamp -3599
transform 1 0 28520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_301
timestamp -3599
transform 1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_304
timestamp -3599
transform 1 0 29072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_312
timestamp -3599
transform 1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_315
timestamp -3599
transform 1 0 30084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_318
timestamp -3599
transform 1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_321
timestamp -3599
transform 1 0 30636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_324
timestamp -3599
transform 1 0 30912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_327
timestamp -3599
transform 1 0 31188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_330
timestamp -3599
transform 1 0 31464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_333
timestamp -3599
transform 1 0 31740 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_336
timestamp -3599
transform 1 0 32016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_339
timestamp -3599
transform 1 0 32292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_343
timestamp -3599
transform 1 0 32660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_346
timestamp -3599
transform 1 0 32936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_349
timestamp -3599
transform 1 0 33212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_352
timestamp -3599
transform 1 0 33488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_355
timestamp -3599
transform 1 0 33764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_358
timestamp -3599
transform 1 0 34040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp -3599
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_368
timestamp -3599
transform 1 0 34960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_371
timestamp -3599
transform 1 0 35236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_380
timestamp -3599
transform 1 0 36064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_383
timestamp -3599
transform 1 0 36340 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_388
timestamp -3599
transform 1 0 36800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_391
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_394
timestamp -3599
transform 1 0 37352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_397
timestamp -3599
transform 1 0 37628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_400
timestamp -3599
transform 1 0 37904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_405
timestamp -3599
transform 1 0 38364 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_408
timestamp -3599
transform 1 0 38640 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_411
timestamp -3599
transform 1 0 38916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_414
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp -3599
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_424
timestamp -3599
transform 1 0 40112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_427
timestamp -3599
transform 1 0 40388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_433
timestamp -3599
transform 1 0 40940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_436
timestamp -3599
transform 1 0 41216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6
timestamp -3599
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_11
timestamp -3599
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_14
timestamp -3599
transform 1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_17
timestamp -3599
transform 1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_20
timestamp -3599
transform 1 0 2944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_23
timestamp -3599
transform 1 0 3220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp -3599
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_35
timestamp -3599
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_38
timestamp -3599
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_41
timestamp -3599
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_44
timestamp -3599
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_47
timestamp -3599
transform 1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_50
timestamp -3599
transform 1 0 5704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp -3599
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_61
timestamp -3599
transform 1 0 6716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_64
timestamp -3599
transform 1 0 6992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_67
timestamp -3599
transform 1 0 7268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_70
timestamp -3599
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_73
timestamp -3599
transform 1 0 7820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_76
timestamp -3599
transform 1 0 8096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_81
timestamp -3599
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_88
timestamp -3599
transform 1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_91
timestamp -3599
transform 1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_94
timestamp -3599
transform 1 0 9752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_97
timestamp -3599
transform 1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_104
timestamp -3599
transform 1 0 10672 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_107
timestamp -3599
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp -3599
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_116
timestamp -3599
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp -3599
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_122
timestamp -3599
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_127
timestamp -3599
transform 1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_130
timestamp -3599
transform 1 0 13064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp -3599
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_136
timestamp -3599
transform 1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_139
timestamp -3599
transform 1 0 13892 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_144
timestamp -3599
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_150
timestamp -3599
transform 1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_153
timestamp -3599
transform 1 0 15180 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_156
timestamp -3599
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_159
timestamp -3599
transform 1 0 15732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_162
timestamp -3599
transform 1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp -3599
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_173
timestamp -3599
transform 1 0 17020 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_176
timestamp -3599
transform 1 0 17296 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_179
timestamp -3599
transform 1 0 17572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_182
timestamp -3599
transform 1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_185
timestamp -3599
transform 1 0 18124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_188
timestamp -3599
transform 1 0 18400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_191
timestamp -3599
transform 1 0 18676 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_200
timestamp -3599
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_203
timestamp -3599
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_206
timestamp -3599
transform 1 0 20056 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_209
timestamp -3599
transform 1 0 20332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_212
timestamp -3599
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_219
timestamp -3599
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_228
timestamp -3599
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_231
timestamp -3599
transform 1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_234
timestamp -3599
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_237
timestamp -3599
transform 1 0 22908 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_242
timestamp -3599
transform 1 0 23368 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_245
timestamp -3599
transform 1 0 23644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_248
timestamp -3599
transform 1 0 23920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_251
timestamp -3599
transform 1 0 24196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_253
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_256
timestamp -3599
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_259
timestamp -3599
transform 1 0 24932 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_265
timestamp -3599
transform 1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_268
timestamp -3599
transform 1 0 25760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_271
timestamp -3599
transform 1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_274
timestamp -3599
transform 1 0 26312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp -3599
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_288
timestamp -3599
transform 1 0 27600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_291
timestamp -3599
transform 1 0 27876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_294
timestamp -3599
transform 1 0 28152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_297
timestamp -3599
transform 1 0 28428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_300
timestamp -3599
transform 1 0 28704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_303
timestamp -3599
transform 1 0 28980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_306
timestamp -3599
transform 1 0 29256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_313
timestamp -3599
transform 1 0 29900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_316
timestamp -3599
transform 1 0 30176 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_319
timestamp -3599
transform 1 0 30452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_322
timestamp -3599
transform 1 0 30728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_325
timestamp -3599
transform 1 0 31004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_328
timestamp -3599
transform 1 0 31280 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp -3599
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_340
timestamp -3599
transform 1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_343
timestamp -3599
transform 1 0 32660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_346
timestamp -3599
transform 1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_349
timestamp -3599
transform 1 0 33212 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_352
timestamp -3599
transform 1 0 33488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_357
timestamp -3599
transform 1 0 33948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_360
timestamp -3599
transform 1 0 34224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_363
timestamp -3599
transform 1 0 34500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_365
timestamp -3599
transform 1 0 34684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_368
timestamp -3599
transform 1 0 34960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_371
timestamp -3599
transform 1 0 35236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_374
timestamp -3599
transform 1 0 35512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_380
timestamp -3599
transform 1 0 36064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_383
timestamp -3599
transform 1 0 36340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_386
timestamp -3599
transform 1 0 36616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_393
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_396
timestamp -3599
transform 1 0 37536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_403
timestamp -3599
transform 1 0 38180 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_406
timestamp -3599
transform 1 0 38456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_409
timestamp -3599
transform 1 0 38732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_412
timestamp -3599
transform 1 0 39008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_415
timestamp -3599
transform 1 0 39284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_418
timestamp -3599
transform 1 0 39560 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_421
timestamp -3599
transform 1 0 39836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_426
timestamp -3599
transform 1 0 40296 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_429
timestamp -3599
transform 1 0 40572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_432
timestamp -3599
transform 1 0 40848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_435
timestamp -3599
transform 1 0 41124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_438
timestamp -3599
transform 1 0 41400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_441
timestamp -3599
transform 1 0 41676 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_444
timestamp -3599
transform 1 0 41952 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp -3599
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_453
timestamp -3599
transform 1 0 42780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_472
timestamp -3599
transform 1 0 44528 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 43884 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 44252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 43884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 43884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 44252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 43884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 44252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 43884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 44252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 43884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 44252 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 44252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 43884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 44252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 43792 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 43424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 43056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 43516 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 43884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 43148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 42780 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 43884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 43884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform -1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 44252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 43884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 44252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform -1 0 4324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform -1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform -1 0 27600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform -1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform -1 0 31832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform -1 0 33948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform -1 0 36064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform -1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 39928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 42412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 44160 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform -1 0 8556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform -1 0 12788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform -1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform -1 0 17020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform -1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform -1 0 23368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 19320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 19872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 21896 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 23368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 23736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 31372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 31096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform -1 0 28888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 36248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 37628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform -1 0 39100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform 1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform 1 0 33672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 36524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 36524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 44896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 44896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 44896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 44896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp -3599
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp -3599
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_46
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_47
timestamp -3599
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_54
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_55
timestamp -3599
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_59
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_62
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_63
timestamp -3599
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_67
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp -3599
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_73
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_77
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp -3599
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_82
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_86
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_87
timestamp -3599
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_89
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_90
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_91
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_92
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_93
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_94
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_95
timestamp -3599
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_96
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_97
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_98
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_103
timestamp -3599
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_106
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_107
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_108
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_109
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_110
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_111
timestamp -3599
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_112
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_114
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_115
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_116
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_118
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_119
timestamp -3599
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_122
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_123
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_124
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_125
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_127
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_128
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_129
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_130
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_131
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp -3599
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp -3599
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1096 120 1216 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 45880 1096 46000 1216 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 45880 3816 46000 3936 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 45880 4088 46000 4208 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 45880 4360 46000 4480 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 45880 4632 46000 4752 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 45880 4904 46000 5024 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 45880 5176 46000 5296 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 45880 5448 46000 5568 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 45880 5720 46000 5840 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 45880 5992 46000 6112 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 45880 6264 46000 6384 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 45880 1368 46000 1488 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 45880 6536 46000 6656 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 45880 6808 46000 6928 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 45880 7080 46000 7200 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 45880 7352 46000 7472 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 45880 7624 46000 7744 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 45880 7896 46000 8016 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 45880 8168 46000 8288 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 45880 8440 46000 8560 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 45880 8712 46000 8832 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 45880 8984 46000 9104 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 45880 1640 46000 1760 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 45880 9256 46000 9376 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 45880 9528 46000 9648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 45880 1912 46000 2032 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 45880 2184 46000 2304 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 45880 2456 46000 2576 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 45880 2728 46000 2848 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 45880 3000 46000 3120 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 45880 3272 46000 3392 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 45880 3544 46000 3664 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 38750 0 38806 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 42430 0 42486 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 42798 0 42854 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 43166 0 43222 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 43534 0 43590 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 43902 0 43958 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 44270 0 44326 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 44638 0 44694 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 45006 0 45062 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 45374 0 45430 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 45742 0 45798 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 39118 0 39174 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 39486 0 39542 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 39854 0 39910 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 40222 0 40278 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 40590 0 40646 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 40958 0 41014 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 41326 0 41382 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 41694 0 41750 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 42062 0 42118 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 3882 11096 3938 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 25042 11096 25098 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 27158 11096 27214 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 29274 11096 29330 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 31390 11096 31446 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 33506 11096 33562 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 35622 11096 35678 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 37738 11096 37794 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 39854 11096 39910 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 41970 11096 42026 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 44086 11096 44142 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 5998 11096 6054 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 8114 11096 8170 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 10230 11096 10286 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 12346 11096 12402 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 14462 11096 14518 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 16578 11096 16634 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 18694 11096 18750 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 20810 11096 20866 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 22926 11096 22982 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 110 0 166 56 0 FreeSans 224 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal2 s 478 0 534 56 0 FreeSans 224 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal2 s 846 0 902 56 0 FreeSans 224 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal2 s 1214 0 1270 56 0 FreeSans 224 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal2 s 4526 0 4582 56 0 FreeSans 224 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal2 s 4894 0 4950 56 0 FreeSans 224 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal2 s 5262 0 5318 56 0 FreeSans 224 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal2 s 5630 0 5686 56 0 FreeSans 224 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal2 s 5998 0 6054 56 0 FreeSans 224 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal2 s 6366 0 6422 56 0 FreeSans 224 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal2 s 6734 0 6790 56 0 FreeSans 224 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal2 s 7102 0 7158 56 0 FreeSans 224 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal2 s 1582 0 1638 56 0 FreeSans 224 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal2 s 1950 0 2006 56 0 FreeSans 224 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal2 s 2318 0 2374 56 0 FreeSans 224 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal2 s 2686 0 2742 56 0 FreeSans 224 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal2 s 3054 0 3110 56 0 FreeSans 224 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal2 s 3422 0 3478 56 0 FreeSans 224 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal2 s 3790 0 3846 56 0 FreeSans 224 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal2 s 4158 0 4214 56 0 FreeSans 224 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal2 s 7470 0 7526 56 0 FreeSans 224 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal2 s 11150 0 11206 56 0 FreeSans 224 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal2 s 11518 0 11574 56 0 FreeSans 224 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal2 s 11886 0 11942 56 0 FreeSans 224 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal2 s 12254 0 12310 56 0 FreeSans 224 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal2 s 12622 0 12678 56 0 FreeSans 224 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal2 s 12990 0 13046 56 0 FreeSans 224 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal2 s 7838 0 7894 56 0 FreeSans 224 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal2 s 8206 0 8262 56 0 FreeSans 224 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal2 s 8574 0 8630 56 0 FreeSans 224 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal2 s 8942 0 8998 56 0 FreeSans 224 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal2 s 9310 0 9366 56 0 FreeSans 224 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal2 s 9678 0 9734 56 0 FreeSans 224 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal2 s 10046 0 10102 56 0 FreeSans 224 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal2 s 10414 0 10470 56 0 FreeSans 224 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal2 s 10782 0 10838 56 0 FreeSans 224 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal2 s 13358 0 13414 56 0 FreeSans 224 0 0 0 NN4END[0]
port 140 nsew signal input
flabel metal2 s 17038 0 17094 56 0 FreeSans 224 0 0 0 NN4END[10]
port 141 nsew signal input
flabel metal2 s 17406 0 17462 56 0 FreeSans 224 0 0 0 NN4END[11]
port 142 nsew signal input
flabel metal2 s 17774 0 17830 56 0 FreeSans 224 0 0 0 NN4END[12]
port 143 nsew signal input
flabel metal2 s 18142 0 18198 56 0 FreeSans 224 0 0 0 NN4END[13]
port 144 nsew signal input
flabel metal2 s 18510 0 18566 56 0 FreeSans 224 0 0 0 NN4END[14]
port 145 nsew signal input
flabel metal2 s 18878 0 18934 56 0 FreeSans 224 0 0 0 NN4END[15]
port 146 nsew signal input
flabel metal2 s 13726 0 13782 56 0 FreeSans 224 0 0 0 NN4END[1]
port 147 nsew signal input
flabel metal2 s 14094 0 14150 56 0 FreeSans 224 0 0 0 NN4END[2]
port 148 nsew signal input
flabel metal2 s 14462 0 14518 56 0 FreeSans 224 0 0 0 NN4END[3]
port 149 nsew signal input
flabel metal2 s 14830 0 14886 56 0 FreeSans 224 0 0 0 NN4END[4]
port 150 nsew signal input
flabel metal2 s 15198 0 15254 56 0 FreeSans 224 0 0 0 NN4END[5]
port 151 nsew signal input
flabel metal2 s 15566 0 15622 56 0 FreeSans 224 0 0 0 NN4END[6]
port 152 nsew signal input
flabel metal2 s 15934 0 15990 56 0 FreeSans 224 0 0 0 NN4END[7]
port 153 nsew signal input
flabel metal2 s 16302 0 16358 56 0 FreeSans 224 0 0 0 NN4END[8]
port 154 nsew signal input
flabel metal2 s 16670 0 16726 56 0 FreeSans 224 0 0 0 NN4END[9]
port 155 nsew signal input
flabel metal2 s 19246 0 19302 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 156 nsew signal output
flabel metal2 s 19614 0 19670 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 157 nsew signal output
flabel metal2 s 19982 0 20038 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 158 nsew signal output
flabel metal2 s 20350 0 20406 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 159 nsew signal output
flabel metal2 s 20718 0 20774 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 160 nsew signal output
flabel metal2 s 21086 0 21142 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 161 nsew signal output
flabel metal2 s 21454 0 21510 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 162 nsew signal output
flabel metal2 s 21822 0 21878 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 163 nsew signal output
flabel metal2 s 22190 0 22246 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 164 nsew signal output
flabel metal2 s 22558 0 22614 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 165 nsew signal output
flabel metal2 s 22926 0 22982 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 166 nsew signal output
flabel metal2 s 23294 0 23350 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 167 nsew signal output
flabel metal2 s 23662 0 23718 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 168 nsew signal output
flabel metal2 s 24030 0 24086 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 169 nsew signal output
flabel metal2 s 24398 0 24454 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 170 nsew signal output
flabel metal2 s 24766 0 24822 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 171 nsew signal output
flabel metal2 s 25134 0 25190 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 172 nsew signal output
flabel metal2 s 25502 0 25558 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 173 nsew signal output
flabel metal2 s 25870 0 25926 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 174 nsew signal output
flabel metal2 s 26238 0 26294 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 175 nsew signal output
flabel metal2 s 26606 0 26662 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 176 nsew signal output
flabel metal2 s 30286 0 30342 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 177 nsew signal output
flabel metal2 s 30654 0 30710 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 178 nsew signal output
flabel metal2 s 31022 0 31078 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 179 nsew signal output
flabel metal2 s 31390 0 31446 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 180 nsew signal output
flabel metal2 s 31758 0 31814 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 181 nsew signal output
flabel metal2 s 32126 0 32182 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 182 nsew signal output
flabel metal2 s 26974 0 27030 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 183 nsew signal output
flabel metal2 s 27342 0 27398 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 184 nsew signal output
flabel metal2 s 27710 0 27766 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 185 nsew signal output
flabel metal2 s 28078 0 28134 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 186 nsew signal output
flabel metal2 s 28446 0 28502 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 187 nsew signal output
flabel metal2 s 28814 0 28870 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 188 nsew signal output
flabel metal2 s 29182 0 29238 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 189 nsew signal output
flabel metal2 s 29550 0 29606 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 190 nsew signal output
flabel metal2 s 29918 0 29974 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 191 nsew signal output
flabel metal2 s 32494 0 32550 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 192 nsew signal output
flabel metal2 s 36174 0 36230 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 193 nsew signal output
flabel metal2 s 36542 0 36598 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 194 nsew signal output
flabel metal2 s 36910 0 36966 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 195 nsew signal output
flabel metal2 s 37278 0 37334 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 196 nsew signal output
flabel metal2 s 37646 0 37702 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 197 nsew signal output
flabel metal2 s 38014 0 38070 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 198 nsew signal output
flabel metal2 s 32862 0 32918 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 199 nsew signal output
flabel metal2 s 33230 0 33286 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 200 nsew signal output
flabel metal2 s 33598 0 33654 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 201 nsew signal output
flabel metal2 s 33966 0 34022 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 202 nsew signal output
flabel metal2 s 34334 0 34390 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 203 nsew signal output
flabel metal2 s 34702 0 34758 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 204 nsew signal output
flabel metal2 s 35070 0 35126 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 205 nsew signal output
flabel metal2 s 35438 0 35494 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 206 nsew signal output
flabel metal2 s 35806 0 35862 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 207 nsew signal output
flabel metal2 s 38382 0 38438 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 1766 11096 1822 11152 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3004 0 3324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 11092 3324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 11092 9324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 11092 15324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 11092 21324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 11092 27324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 11092 33324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11152 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 11092 39324 11152 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 11092 2264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 11092 8264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 11092 14264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 11092 20264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 11092 26264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 11092 32264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 11092 38264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 0 44264 11152 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 0 44264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 43944 11092 44264 11152 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 23000 8704 23000 8704 0 VGND
rlabel metal1 23000 8160 23000 8160 0 VPWR
rlabel metal3 1356 1156 1356 1156 0 FrameData[0]
rlabel metal3 919 3876 919 3876 0 FrameData[10]
rlabel metal3 712 4148 712 4148 0 FrameData[11]
rlabel metal3 436 4420 436 4420 0 FrameData[12]
rlabel metal2 5566 5695 5566 5695 0 FrameData[13]
rlabel metal3 919 4964 919 4964 0 FrameData[14]
rlabel metal2 4370 5763 4370 5763 0 FrameData[15]
rlabel metal3 712 5508 712 5508 0 FrameData[16]
rlabel via2 43194 5763 43194 5763 0 FrameData[17]
rlabel metal3 390 6052 390 6052 0 FrameData[18]
rlabel metal1 43056 5202 43056 5202 0 FrameData[19]
rlabel metal3 666 1428 666 1428 0 FrameData[1]
rlabel metal3 574 6596 574 6596 0 FrameData[20]
rlabel metal3 712 6868 712 6868 0 FrameData[21]
rlabel via2 42458 4675 42458 4675 0 FrameData[22]
rlabel metal3 712 7412 712 7412 0 FrameData[23]
rlabel metal1 1978 6834 1978 6834 0 FrameData[24]
rlabel via2 42826 6307 42826 6307 0 FrameData[25]
rlabel metal3 712 8228 712 8228 0 FrameData[26]
rlabel metal2 41630 8279 41630 8279 0 FrameData[27]
rlabel metal3 574 8772 574 8772 0 FrameData[28]
rlabel metal2 2898 8415 2898 8415 0 FrameData[29]
rlabel metal3 252 1700 252 1700 0 FrameData[2]
rlabel metal3 436 9316 436 9316 0 FrameData[30]
rlabel metal3 666 9588 666 9588 0 FrameData[31]
rlabel metal3 620 1972 620 1972 0 FrameData[3]
rlabel metal3 712 2244 712 2244 0 FrameData[4]
rlabel metal2 43194 2975 43194 2975 0 FrameData[5]
rlabel metal3 942 2788 942 2788 0 FrameData[6]
rlabel via2 41722 3043 41722 3043 0 FrameData[7]
rlabel metal2 41538 3587 41538 3587 0 FrameData[8]
rlabel metal3 758 3604 758 3604 0 FrameData[9]
rlabel metal3 45380 1156 45380 1156 0 FrameData_O[0]
rlabel metal3 45449 3876 45449 3876 0 FrameData_O[10]
rlabel metal3 45196 4148 45196 4148 0 FrameData_O[11]
rlabel metal3 45012 4420 45012 4420 0 FrameData_O[12]
rlabel metal3 45196 4692 45196 4692 0 FrameData_O[13]
rlabel metal3 45449 4964 45449 4964 0 FrameData_O[14]
rlabel metal3 45196 5236 45196 5236 0 FrameData_O[15]
rlabel metal3 45564 5508 45564 5508 0 FrameData_O[16]
rlabel metal3 45196 5780 45196 5780 0 FrameData_O[17]
rlabel metal3 45449 6052 45449 6052 0 FrameData_O[18]
rlabel metal3 45196 6324 45196 6324 0 FrameData_O[19]
rlabel metal3 44644 1428 44644 1428 0 FrameData_O[1]
rlabel via2 44114 6613 44114 6613 0 FrameData_O[20]
rlabel metal2 44482 6749 44482 6749 0 FrameData_O[21]
rlabel metal3 45196 7140 45196 7140 0 FrameData_O[22]
rlabel metal3 45104 7412 45104 7412 0 FrameData_O[23]
rlabel metal3 45196 7684 45196 7684 0 FrameData_O[24]
rlabel metal3 45426 7956 45426 7956 0 FrameData_O[25]
rlabel metal3 45334 8228 45334 8228 0 FrameData_O[26]
rlabel metal3 44598 8500 44598 8500 0 FrameData_O[27]
rlabel metal2 43746 8415 43746 8415 0 FrameData_O[28]
rlabel metal1 43884 7514 43884 7514 0 FrameData_O[29]
rlabel metal3 44460 1700 44460 1700 0 FrameData_O[2]
rlabel metal2 43378 8653 43378 8653 0 FrameData_O[30]
rlabel metal1 43010 7922 43010 7922 0 FrameData_O[31]
rlabel metal1 44252 2822 44252 2822 0 FrameData_O[3]
rlabel metal3 45012 2244 45012 2244 0 FrameData_O[4]
rlabel metal3 45058 2516 45058 2516 0 FrameData_O[5]
rlabel metal3 45196 2788 45196 2788 0 FrameData_O[6]
rlabel metal3 45242 3060 45242 3060 0 FrameData_O[7]
rlabel metal3 45012 3332 45012 3332 0 FrameData_O[8]
rlabel metal3 45196 3604 45196 3604 0 FrameData_O[9]
rlabel metal1 37214 7378 37214 7378 0 FrameStrobe[0]
rlabel metal2 42412 3196 42412 3196 0 FrameStrobe[10]
rlabel metal2 42872 3332 42872 3332 0 FrameStrobe[11]
rlabel metal1 42274 7378 42274 7378 0 FrameStrobe[12]
rlabel metal3 39238 5236 39238 5236 0 FrameStrobe[13]
rlabel metal3 40572 5644 40572 5644 0 FrameStrobe[14]
rlabel metal2 36018 4556 36018 4556 0 FrameStrobe[15]
rlabel metal2 44712 3196 44712 3196 0 FrameStrobe[16]
rlabel metal1 42504 6970 42504 6970 0 FrameStrobe[17]
rlabel metal1 41722 7514 41722 7514 0 FrameStrobe[18]
rlabel metal1 44712 4522 44712 4522 0 FrameStrobe[19]
rlabel metal2 36662 7616 36662 7616 0 FrameStrobe[1]
rlabel metal2 39514 123 39514 123 0 FrameStrobe[2]
rlabel metal2 39882 140 39882 140 0 FrameStrobe[3]
rlabel metal2 14306 7684 14306 7684 0 FrameStrobe[4]
rlabel metal2 35098 3740 35098 3740 0 FrameStrobe[5]
rlabel metal1 39192 6086 39192 6086 0 FrameStrobe[6]
rlabel metal1 40434 6154 40434 6154 0 FrameStrobe[7]
rlabel metal2 41676 2924 41676 2924 0 FrameStrobe[8]
rlabel metal1 40848 6222 40848 6222 0 FrameStrobe[9]
rlabel metal1 4002 8602 4002 8602 0 FrameStrobe_O[0]
rlabel metal1 25162 8602 25162 8602 0 FrameStrobe_O[10]
rlabel metal2 27370 9863 27370 9863 0 FrameStrobe_O[11]
rlabel metal1 29486 8602 29486 8602 0 FrameStrobe_O[12]
rlabel metal1 31510 8602 31510 8602 0 FrameStrobe_O[13]
rlabel metal1 33626 8602 33626 8602 0 FrameStrobe_O[14]
rlabel metal1 35742 8602 35742 8602 0 FrameStrobe_O[15]
rlabel metal1 37858 8602 37858 8602 0 FrameStrobe_O[16]
rlabel metal1 40020 8602 40020 8602 0 FrameStrobe_O[17]
rlabel metal1 42320 8602 42320 8602 0 FrameStrobe_O[18]
rlabel metal1 44252 8602 44252 8602 0 FrameStrobe_O[19]
rlabel metal1 6256 8602 6256 8602 0 FrameStrobe_O[1]
rlabel metal1 8234 8602 8234 8602 0 FrameStrobe_O[2]
rlabel metal1 10350 8602 10350 8602 0 FrameStrobe_O[3]
rlabel metal2 12374 9856 12374 9856 0 FrameStrobe_O[4]
rlabel metal1 14582 8602 14582 8602 0 FrameStrobe_O[5]
rlabel metal1 16698 8602 16698 8602 0 FrameStrobe_O[6]
rlabel metal1 18814 8602 18814 8602 0 FrameStrobe_O[7]
rlabel metal1 20930 8602 20930 8602 0 FrameStrobe_O[8]
rlabel metal1 23046 8602 23046 8602 0 FrameStrobe_O[9]
rlabel metal2 138 1704 138 1704 0 N1END[0]
rlabel metal2 506 2350 506 2350 0 N1END[1]
rlabel metal2 874 2282 874 2282 0 N1END[2]
rlabel metal2 1242 55 1242 55 0 N1END[3]
rlabel metal1 8234 4794 8234 4794 0 N2END[0]
rlabel metal1 5796 4522 5796 4522 0 N2END[1]
rlabel metal1 6486 4114 6486 4114 0 N2END[2]
rlabel metal1 7774 4046 7774 4046 0 N2END[3]
rlabel metal2 6026 1401 6026 1401 0 N2END[4]
rlabel metal1 20470 5134 20470 5134 0 N2END[5]
rlabel metal2 19642 3774 19642 3774 0 N2END[6]
rlabel metal2 7130 2860 7130 2860 0 N2END[7]
rlabel metal2 1610 327 1610 327 0 N2MID[0]
rlabel metal2 1978 1075 1978 1075 0 N2MID[1]
rlabel metal2 2346 1075 2346 1075 0 N2MID[2]
rlabel metal2 2714 3676 2714 3676 0 N2MID[3]
rlabel metal2 3082 55 3082 55 0 N2MID[4]
rlabel metal2 3450 55 3450 55 0 N2MID[5]
rlabel metal1 13409 7378 13409 7378 0 N2MID[6]
rlabel metal2 18170 6460 18170 6460 0 N2MID[7]
rlabel metal1 9706 4522 9706 4522 0 N4END[0]
rlabel metal2 11178 191 11178 191 0 N4END[10]
rlabel metal2 11546 259 11546 259 0 N4END[11]
rlabel metal2 11914 803 11914 803 0 N4END[12]
rlabel metal2 12282 3132 12282 3132 0 N4END[13]
rlabel metal2 12650 3744 12650 3744 0 N4END[14]
rlabel metal2 13018 582 13018 582 0 N4END[15]
rlabel metal2 7866 1401 7866 1401 0 N4END[1]
rlabel metal2 8234 1194 8234 1194 0 N4END[2]
rlabel metal2 8602 1007 8602 1007 0 N4END[3]
rlabel metal2 8970 140 8970 140 0 N4END[4]
rlabel metal2 9338 956 9338 956 0 N4END[5]
rlabel metal2 16422 4386 16422 4386 0 N4END[6]
rlabel metal2 10074 1296 10074 1296 0 N4END[7]
rlabel metal2 10442 123 10442 123 0 N4END[8]
rlabel metal2 14766 2992 14766 2992 0 N4END[9]
rlabel metal1 41308 4590 41308 4590 0 NN4END[0]
rlabel metal1 43838 7310 43838 7310 0 NN4END[10]
rlabel metal2 17434 2095 17434 2095 0 NN4END[11]
rlabel metal2 17802 871 17802 871 0 NN4END[12]
rlabel metal2 18170 1401 18170 1401 0 NN4END[13]
rlabel metal2 18538 3200 18538 3200 0 NN4END[14]
rlabel metal2 18906 939 18906 939 0 NN4END[15]
rlabel metal2 13754 106 13754 106 0 NN4END[1]
rlabel metal1 39008 4590 39008 4590 0 NN4END[2]
rlabel metal1 15732 3434 15732 3434 0 NN4END[3]
rlabel metal1 16790 3162 16790 3162 0 NN4END[4]
rlabel metal1 34132 3366 34132 3366 0 NN4END[5]
rlabel metal1 34684 3502 34684 3502 0 NN4END[6]
rlabel metal2 15962 174 15962 174 0 NN4END[7]
rlabel metal2 16330 208 16330 208 0 NN4END[8]
rlabel metal1 18630 4998 18630 4998 0 NN4END[9]
rlabel metal1 19412 2822 19412 2822 0 S1BEG[0]
rlabel metal2 19642 1160 19642 1160 0 S1BEG[1]
rlabel metal2 20010 1160 20010 1160 0 S1BEG[2]
rlabel metal2 20378 1160 20378 1160 0 S1BEG[3]
rlabel metal2 20746 1160 20746 1160 0 S2BEG[0]
rlabel metal2 21114 55 21114 55 0 S2BEG[1]
rlabel metal2 21482 1160 21482 1160 0 S2BEG[2]
rlabel metal2 21850 1160 21850 1160 0 S2BEG[3]
rlabel metal2 22218 1160 22218 1160 0 S2BEG[4]
rlabel metal2 22586 1160 22586 1160 0 S2BEG[5]
rlabel metal2 22954 1296 22954 1296 0 S2BEG[6]
rlabel metal2 23322 1160 23322 1160 0 S2BEG[7]
rlabel metal2 23690 1160 23690 1160 0 S2BEGb[0]
rlabel metal2 24058 1160 24058 1160 0 S2BEGb[1]
rlabel metal2 24426 55 24426 55 0 S2BEGb[2]
rlabel metal2 24794 1296 24794 1296 0 S2BEGb[3]
rlabel metal2 25162 1160 25162 1160 0 S2BEGb[4]
rlabel metal2 25530 55 25530 55 0 S2BEGb[5]
rlabel metal2 25898 55 25898 55 0 S2BEGb[6]
rlabel metal2 26266 55 26266 55 0 S2BEGb[7]
rlabel metal2 26634 1296 26634 1296 0 S4BEG[0]
rlabel metal2 30314 1296 30314 1296 0 S4BEG[10]
rlabel metal2 30682 55 30682 55 0 S4BEG[11]
rlabel metal1 31188 2822 31188 2822 0 S4BEG[12]
rlabel metal2 31418 55 31418 55 0 S4BEG[13]
rlabel metal2 31786 1296 31786 1296 0 S4BEG[14]
rlabel metal2 32154 55 32154 55 0 S4BEG[15]
rlabel metal2 27002 55 27002 55 0 S4BEG[1]
rlabel metal2 27370 55 27370 55 0 S4BEG[2]
rlabel metal2 27738 1296 27738 1296 0 S4BEG[3]
rlabel metal2 28106 55 28106 55 0 S4BEG[4]
rlabel metal1 28566 2822 28566 2822 0 S4BEG[5]
rlabel metal2 28842 1296 28842 1296 0 S4BEG[6]
rlabel metal2 29210 1160 29210 1160 0 S4BEG[7]
rlabel metal2 29578 599 29578 599 0 S4BEG[8]
rlabel metal2 29946 599 29946 599 0 S4BEG[9]
rlabel metal2 32522 599 32522 599 0 SS4BEG[0]
rlabel metal1 36340 2822 36340 2822 0 SS4BEG[10]
rlabel metal2 36570 55 36570 55 0 SS4BEG[11]
rlabel metal2 36938 1296 36938 1296 0 SS4BEG[12]
rlabel metal2 37306 55 37306 55 0 SS4BEG[13]
rlabel metal2 37674 1330 37674 1330 0 SS4BEG[14]
rlabel metal2 38042 1296 38042 1296 0 SS4BEG[15]
rlabel metal2 32890 599 32890 599 0 SS4BEG[1]
rlabel metal2 33258 55 33258 55 0 SS4BEG[2]
rlabel metal1 33764 2822 33764 2822 0 SS4BEG[3]
rlabel metal2 33994 55 33994 55 0 SS4BEG[4]
rlabel metal2 34362 1296 34362 1296 0 SS4BEG[5]
rlabel metal2 34730 55 34730 55 0 SS4BEG[6]
rlabel metal2 35098 1194 35098 1194 0 SS4BEG[7]
rlabel metal2 35466 55 35466 55 0 SS4BEG[8]
rlabel metal2 35834 1330 35834 1330 0 SS4BEG[9]
rlabel metal1 37582 7786 37582 7786 0 UserCLK
rlabel metal1 1840 8602 1840 8602 0 UserCLKo
rlabel metal2 17250 4964 17250 4964 0 net1
rlabel via2 2346 4539 2346 4539 0 net10
rlabel metal2 42964 2924 42964 2924 0 net100
rlabel metal1 34684 2482 34684 2482 0 net101
rlabel metal1 32706 6630 32706 6630 0 net102
rlabel metal1 38456 7718 38456 7718 0 net103
rlabel metal1 35742 3706 35742 3706 0 net104
rlabel metal1 2070 8432 2070 8432 0 net105
rlabel metal2 43286 5780 43286 5780 0 net11
rlabel metal1 12420 2856 12420 2856 0 net12
rlabel metal2 41538 6256 41538 6256 0 net13
rlabel metal1 44298 6800 44298 6800 0 net14
rlabel metal1 43608 4726 43608 4726 0 net15
rlabel metal2 39790 8092 39790 8092 0 net16
rlabel metal1 43608 4998 43608 4998 0 net17
rlabel metal1 43470 6426 43470 6426 0 net18
rlabel metal1 43102 8058 43102 8058 0 net19
rlabel metal2 43470 3638 43470 3638 0 net2
rlabel metal1 42274 8058 42274 8058 0 net20
rlabel metal1 43562 7786 43562 7786 0 net21
rlabel metal2 36478 7684 36478 7684 0 net22
rlabel metal1 27025 1598 27025 1598 0 net23
rlabel via2 2714 7939 2714 7939 0 net24
rlabel metal1 42826 7888 42826 7888 0 net25
rlabel metal2 2346 3366 2346 3366 0 net26
rlabel metal1 4853 2346 4853 2346 0 net27
rlabel metal1 42872 2482 42872 2482 0 net28
rlabel metal1 44298 2992 44298 2992 0 net29
rlabel metal1 43194 3706 43194 3706 0 net3
rlabel metal1 43654 3094 43654 3094 0 net30
rlabel metal2 42274 3298 42274 3298 0 net31
rlabel metal1 44528 3502 44528 3502 0 net32
rlabel metal2 35466 8296 35466 8296 0 net33
rlabel metal2 40710 6663 40710 6663 0 net34
rlabel metal1 40572 6630 40572 6630 0 net35
rlabel metal1 39928 7174 39928 7174 0 net36
rlabel metal2 32430 8092 32430 8092 0 net37
rlabel metal2 34730 8092 34730 8092 0 net38
rlabel metal2 35834 8092 35834 8092 0 net39
rlabel metal1 43654 4250 43654 4250 0 net4
rlabel metal1 38226 8058 38226 8058 0 net40
rlabel metal1 39928 8058 39928 8058 0 net41
rlabel metal2 40894 8262 40894 8262 0 net42
rlabel metal1 43700 4794 43700 4794 0 net43
rlabel metal1 34960 7786 34960 7786 0 net44
rlabel metal2 9982 8262 9982 8262 0 net45
rlabel metal2 12006 8262 12006 8262 0 net46
rlabel metal1 13984 7718 13984 7718 0 net47
rlabel metal1 16606 5576 16606 5576 0 net48
rlabel metal1 36938 6358 36938 6358 0 net49
rlabel metal2 36846 6120 36846 6120 0 net5
rlabel metal1 36570 6120 36570 6120 0 net50
rlabel metal1 37996 6426 37996 6426 0 net51
rlabel metal1 38456 6154 38456 6154 0 net52
rlabel metal1 19366 2992 19366 2992 0 net53
rlabel metal2 19550 3774 19550 3774 0 net54
rlabel metal1 19826 2448 19826 2448 0 net55
rlabel metal1 17618 2346 17618 2346 0 net56
rlabel metal1 19504 6086 19504 6086 0 net57
rlabel metal1 20792 2482 20792 2482 0 net58
rlabel metal1 20286 2550 20286 2550 0 net59
rlabel metal2 37214 5610 37214 5610 0 net6
rlabel metal1 17204 7786 17204 7786 0 net60
rlabel metal2 19872 2516 19872 2516 0 net61
rlabel metal1 22678 2516 22678 2516 0 net62
rlabel metal1 5704 3910 5704 3910 0 net63
rlabel metal1 21804 2822 21804 2822 0 net64
rlabel metal2 21482 4046 21482 4046 0 net65
rlabel metal1 22126 3366 22126 3366 0 net66
rlabel metal1 24196 2482 24196 2482 0 net67
rlabel metal1 23874 5542 23874 5542 0 net68
rlabel metal1 15410 1802 15410 1802 0 net69
rlabel metal1 44298 5168 44298 5168 0 net7
rlabel metal1 15318 1734 15318 1734 0 net70
rlabel metal2 24150 1887 24150 1887 0 net71
rlabel metal1 25990 2482 25990 2482 0 net72
rlabel metal1 25300 6154 25300 6154 0 net73
rlabel metal2 16238 4896 16238 4896 0 net74
rlabel metal1 31004 2346 31004 2346 0 net75
rlabel metal1 31004 3026 31004 3026 0 net76
rlabel metal2 32154 2108 32154 2108 0 net77
rlabel via2 32522 2397 32522 2397 0 net78
rlabel metal2 32890 2465 32890 2465 0 net79
rlabel metal2 41446 5355 41446 5355 0 net8
rlabel metal1 27830 2414 27830 2414 0 net80
rlabel metal1 27462 2618 27462 2618 0 net81
rlabel metal1 27968 2482 27968 2482 0 net82
rlabel metal1 28796 2414 28796 2414 0 net83
rlabel metal1 28750 3026 28750 3026 0 net84
rlabel metal1 29394 3366 29394 3366 0 net85
rlabel metal1 29854 3366 29854 3366 0 net86
rlabel metal1 16928 3366 16928 3366 0 net87
rlabel metal1 17158 4454 17158 4454 0 net88
rlabel metal1 33120 2414 33120 2414 0 net89
rlabel metal1 44298 5644 44298 5644 0 net9
rlabel metal2 36294 3196 36294 3196 0 net90
rlabel metal1 36984 2414 36984 2414 0 net91
rlabel metal1 35098 2074 35098 2074 0 net92
rlabel metal1 39008 4454 39008 4454 0 net93
rlabel metal1 38456 3910 38456 3910 0 net94
rlabel metal1 40158 2414 40158 2414 0 net95
rlabel metal2 32798 4287 32798 4287 0 net96
rlabel metal2 33994 4964 33994 4964 0 net97
rlabel metal2 33718 5100 33718 5100 0 net98
rlabel metal1 33166 5542 33166 5542 0 net99
<< properties >>
string FIXED_BBOX 0 0 46000 11152
<< end >>
