module N_term_single (Ci,
    UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 input Ci;
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 sky130_fd_sc_hd__buf_1 _000_ (.A(FrameData[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 _001_ (.A(FrameData[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 _002_ (.A(FrameData[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 _003_ (.A(FrameData[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 _004_ (.A(FrameData[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 _005_ (.A(FrameData[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 _006_ (.A(FrameData[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 _007_ (.A(FrameData[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 _008_ (.A(FrameData[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 _009_ (.A(FrameData[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 _010_ (.A(FrameData[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 _011_ (.A(FrameData[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 _012_ (.A(FrameData[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 _013_ (.A(FrameData[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 _014_ (.A(FrameData[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 _015_ (.A(FrameData[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 _016_ (.A(FrameData[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 _017_ (.A(FrameData[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 _018_ (.A(FrameData[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 _019_ (.A(FrameData[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 _020_ (.A(FrameData[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 _021_ (.A(FrameData[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 _022_ (.A(FrameData[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 _023_ (.A(FrameData[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 _024_ (.A(FrameData[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 _025_ (.A(FrameData[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 _026_ (.A(FrameData[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 _027_ (.A(FrameData[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 _028_ (.A(FrameData[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 _029_ (.A(FrameData[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 _030_ (.A(FrameData[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 _031_ (.A(FrameData[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 _032_ (.A(FrameStrobe[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 _033_ (.A(FrameStrobe[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 _034_ (.A(FrameStrobe[2]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 _035_ (.A(FrameStrobe[3]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 _036_ (.A(FrameStrobe[4]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 _037_ (.A(FrameStrobe[5]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 _038_ (.A(FrameStrobe[6]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 _039_ (.A(FrameStrobe[7]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _040_ (.A(FrameStrobe[8]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _041_ (.A(FrameStrobe[9]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _042_ (.A(FrameStrobe[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 _043_ (.A(FrameStrobe[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 _044_ (.A(FrameStrobe[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 _045_ (.A(FrameStrobe[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 _046_ (.A(FrameStrobe[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 _047_ (.A(FrameStrobe[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 _048_ (.A(FrameStrobe[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 _049_ (.A(FrameStrobe[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 _050_ (.A(FrameStrobe[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _051_ (.A(FrameStrobe[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 _052_ (.A(N1END[3]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 _053_ (.A(N1END[2]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 _054_ (.A(N1END[1]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 _055_ (.A(N1END[0]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 _056_ (.A(N2MID[7]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 _057_ (.A(N2MID[6]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 _058_ (.A(N2MID[5]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 _059_ (.A(N2MID[4]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 _060_ (.A(N2MID[3]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 _061_ (.A(N2MID[2]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 _062_ (.A(N2MID[1]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 _063_ (.A(N2MID[0]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 _064_ (.A(N2END[7]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 _065_ (.A(N2END[6]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 _066_ (.A(N2END[5]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 _067_ (.A(N2END[4]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _068_ (.A(N2END[3]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 _069_ (.A(N2END[2]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 _070_ (.A(N2END[1]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 _071_ (.A(N2END[0]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _072_ (.A(N4END[15]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _073_ (.A(N4END[14]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _074_ (.A(N4END[13]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(N4END[12]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _076_ (.A(N4END[11]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _077_ (.A(N4END[10]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _078_ (.A(N4END[9]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(N4END[8]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _080_ (.A(N4END[7]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _081_ (.A(N4END[6]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _082_ (.A(N4END[5]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _083_ (.A(N4END[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _084_ (.A(N4END[3]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _085_ (.A(N4END[2]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _086_ (.A(N4END[1]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _087_ (.A(N4END[0]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(NN4END[15]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(NN4END[14]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _090_ (.A(NN4END[13]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _091_ (.A(NN4END[12]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _092_ (.A(NN4END[11]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _093_ (.A(NN4END[10]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _094_ (.A(NN4END[9]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _095_ (.A(NN4END[8]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(NN4END[7]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _097_ (.A(NN4END[6]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 _098_ (.A(NN4END[5]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _099_ (.A(NN4END[4]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _100_ (.A(NN4END[3]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _101_ (.A(NN4END[2]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _102_ (.A(NN4END[1]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _103_ (.A(NN4END[0]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 _104_ (.A(UserCLK),
    .X(net105));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_107 ();
 sky130_fd_sc_hd__buf_2 output1 (.A(net1),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(UserCLKo));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(FrameData[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameData[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(FrameData[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(FrameData[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(FrameData[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameData[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(FrameData[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(FrameData[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(FrameData[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(FrameData[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(FrameData[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(FrameData[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(FrameData[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(FrameData[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(FrameData[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(FrameData[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(FrameData[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(FrameData[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(FrameData[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(FrameData[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(FrameData[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(FrameData[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(FrameData[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(FrameStrobe[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(FrameStrobe[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(NN4END[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(NN4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(NN4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(NN4END[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(NN4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(NN4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(NN4END[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(FrameData[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(NN4END[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(UserCLK));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
endmodule
