* NGSPICE file created from LUT4AB.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt LUT4AB Ci Co E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2]
+ E1END[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7]
+ E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7]
+ E2END[0] E2END[1] E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0]
+ E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10]
+ E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8]
+ E6BEG[9] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5]
+ E6END[6] E6END[7] E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13]
+ EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6]
+ EE4BEG[7] EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13]
+ EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6]
+ EE4END[7] EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4]
+ N2END[5] N2END[6] N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5]
+ N2MID[6] N2MID[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3]
+ S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4]
+ S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5]
+ S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6]
+ S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1]
+ S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11]
+ SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4]
+ SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0]
+ W1BEG[1] W1BEG[2] W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1]
+ W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2]
+ W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3]
+ W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4]
+ W2MID[5] W2MID[6] W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3]
+ W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11]
+ W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9]
+ WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1]
+ WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9]
+ WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1]
+ WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
XFILLER_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2106_ net799 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2037_ net746 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_20_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1270_ net633 net628 net619 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_59_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0985_ _0115_ _0116_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q VGND VGND VPWR VPWR
+ _0117_ sky130_fd_sc_hd__mux2_1
X_1606_ net773 net711 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
X_1537_ net784 net700 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1468_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q _0527_ VGND VGND VPWR VPWR _0528_
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1399_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q _0638_ _0489_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__a211oi_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout650 net651 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__buf_2
Xfanout683 net686 VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__clkbuf_2
Xfanout661 net58 VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__buf_2
Xfanout694 FrameStrobe[2] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__clkbuf_2
Xfanout672 net673 VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0770_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _0618_ VGND VGND VPWR VPWR _0619_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1322_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q _0421_ _0423_ _0425_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q
+ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__o221a_1
X_1253_ net87 net89 net91 net115 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux4_1
XFILLER_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1184_ Inst_LH_LUT4c_frame_config_dffesr.LUT_flop _0574_ _0302_ VGND VGND VPWR VPWR
+ H sky130_fd_sc_hd__o21ba_4
XPHY_EDGE_ROW_20_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0968_ _0086_ _0099_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__or2_1
X_0899_ net86 net3 net9 net23 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux4_1
Xoutput231 net231 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput220 net220 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
Xoutput253 Inst_LUT4AB_switch_matrix.JN2BEG7 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__buf_6
Xoutput242 net242 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__buf_4
Xoutput286 net286 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput275 net275 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput264 net264 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput297 Inst_LUT4AB_switch_matrix.S1BEG3 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__buf_8
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1940_ net748 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1871_ net802 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0822_ net95 net123 net107 net139 Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
+ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__mux4_1
X_0753_ net26 net109 net126 Inst_LUT4AB_switch_matrix.E2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__mux4_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2354_ net129 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_2
X_1305_ net807 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__o21ba_1
X_2285_ Inst_LUT4AB_switch_matrix.NN4BEG2 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_67_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1236_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0349_ VGND VGND VPWR VPWR _0350_
+ sky130_fd_sc_hd__and2b_1
X_1167_ _0281_ _0282_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__nand2_1
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1098_ net77 net105 net20 Inst_LUT4AB_switch_matrix.JN2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__mux4_2
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2070_ net744 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1021_ net86 net97 net12 net125 Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q
+ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__mux4_1
XFILLER_46_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ net778 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1854_ net790 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1785_ net800 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0805_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0628_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__mux2_1
X_0736_ net462 net628 net619 net404 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__mux4_1
X_2337_ Inst_LUT4AB_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__buf_1
XFILLER_37_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1219_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q _0332_ _0334_ VGND VGND VPWR VPWR
+ _0335_ sky130_fd_sc_hd__a21oi_4
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2199_ net788 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1570_ net782 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_60_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2122_ net764 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2053_ net774 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1004_ _0132_ _0133_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VGND VGND VPWR VPWR
+ _0134_ sky130_fd_sc_hd__mux2_1
XFILLER_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1906_ net752 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer118 net513 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer129 net402 VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd1_1
X_1837_ net757 net664 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1768_ net768 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1699_ net778 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0719_ net131 VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__inv_1
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput120 W2END[1] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
Xinput131 W2MID[4] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_2
XFILLER_48_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ net745 net712 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1553_ net759 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_1484_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q _0529_ VGND VGND VPWR VPWR _0543_
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2105_ net801 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2036_ net748 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ net87 net89 net97 net660 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__mux4_1
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1605_ net775 net710 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_1536_ net787 net703 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_1467_ _0524_ _0525_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q VGND VGND VPWR VPWR
+ _0527_ sky130_fd_sc_hd__mux2_1
X_1398_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q net622 VGND VGND VPWR VPWR _0489_
+ sky130_fd_sc_hd__nor2_1
XFILLER_67_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2019_ net779 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout651 net652 VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkbuf_4
Xfanout640 net641 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__clkbuf_2
Xfanout684 net686 VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__buf_2
Xfanout673 FrameStrobe[7] VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__clkbuf_2
Xfanout662 net664 VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout695 net697 VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__buf_2
XFILLER_73_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1321_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q _0424_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q
+ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__a21bo_1
X_1252_ net59 net83 net2 net6 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux4_1
X_1183_ _0289_ _0301_ _0574_ _0294_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__o211a_1
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0967_ _0098_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ net94 net122 net110 net136 Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q
+ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux4_1
Xoutput210 net210 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput232 net232 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput221 net221 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
Xoutput243 Inst_LUT4AB_switch_matrix.N1BEG1 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__buf_4
Xoutput254 net254 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput276 net276 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput265 net265 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__buf_4
X_1519_ net803 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
Xoutput298 net298 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_8
Xoutput287 net287 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1870_ net754 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0821_ net61 net10 net67 net805 Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
+ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__mux4_1
X_0752_ _0599_ _0597_ _0602_ _0566_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG1
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2353_ net128 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_2
X_1304_ net660 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q VGND VGND VPWR VPWR _0409_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_67_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1235_ net655 net650 net625 net640 Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__mux4_1
XFILLER_64_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1166_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 _0283_ _0284_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__o22a_1
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1097_ _0220_ _0217_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.JN2BEG6 sky130_fd_sc_hd__mux2_4
XFILLER_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1999_ net802 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1020_ net9 net139 net114 Inst_LUT4AB_switch_matrix.JN2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_64_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ net782 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1853_ net792 net666 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0804_ _0639_ _0640_ _0649_ _0648_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q
+ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux4_2
X_1784_ net740 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0735_ net433 net648 net463 net643 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__mux4_2
X_2267_ Inst_LUT4AB_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_2
X_1218_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q _0333_ VGND VGND VPWR VPWR _0334_
+ sky130_fd_sc_hd__and2b_1
XFILLER_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2198_ net790 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_1
X_1149_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0250_ _0239_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__mux4_1
XFILLER_40_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2121_ net43 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2052_ net777 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1003_ net478 net630 net621 net618 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_49_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1905_ net759 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer119 net514 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1836_ net760 net664 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1767_ net771 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0718_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__inv_1
X_1698_ net782 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2319_ Inst_LUT4AB_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput110 S4END[3] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xinput121 W2END[2] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_2
Xinput132 W2MID[5] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1621_ net747 net712 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
X_1552_ net781 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
X_1483_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q _0538_ VGND VGND VPWR VPWR _0542_
+ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2104_ net740 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2035_ net750 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1819_ net796 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout800 net801 VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__buf_4
XFILLER_45_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer9 Inst_LUT4AB_switch_matrix.M_AH VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_59_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ net61 net69 net807 net12 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__mux4_1
X_1604_ net776 net709 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1535_ net788 net703 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_1466_ Inst_LUT4AB_switch_matrix.JN2BEG2 Inst_LUT4AB_switch_matrix.JS2BEG2 Inst_LUT4AB_switch_matrix.E2BEG2
+ Inst_LUT4AB_switch_matrix.JW2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q
+ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__mux4_2
X_1397_ net62 net806 net90 net656 Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux4_1
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2018_ net783 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold150 Inst_LC_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout630 net632 VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__buf_2
Xfanout641 net642 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__buf_2
Xfanout652 B VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__buf_8
Xfanout674 net677 VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__clkbuf_2
Xfanout663 net664 VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__clkbuf_1
Xfanout685 net686 VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__clkbuf_2
Xfanout696 net697 VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1320_ _0097_ net658 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q VGND VGND VPWR VPWR
+ _0424_ sky130_fd_sc_hd__mux2_1
X_1251_ _0361_ _0362_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VGND VGND VPWR VPWR
+ _0363_ sky130_fd_sc_hd__mux2_4
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1182_ _0297_ _0300_ _0280_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__mux2_1
XFILLER_64_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0966_ _0096_ _0097_ _0088_ _0087_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux4_2
X_0897_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q _0033_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q
+ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__a21bo_1
Xoutput200 net200 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
Xoutput222 net222 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput233 net233 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput211 net211 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput244 net244 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__buf_4
Xoutput255 net255 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput277 net277 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput266 Inst_LUT4AB_switch_matrix.N4BEG1 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_6
X_1518_ net755 net56 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
Xoutput299 net299 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__buf_6
Xoutput288 net288 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__buf_2
X_1449_ net415 _0068_ Inst_LUT4AB_switch_matrix.E2BEG0 _0084_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0820_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0664_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__a21bo_1
X_0751_ _0600_ _0601_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q VGND VGND VPWR VPWR
+ _0602_ sky130_fd_sc_hd__mux2_1
X_2352_ net127 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__buf_1
X_1303_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0407_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q
+ _0406_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__o211a_1
X_2283_ Inst_LUT4AB_switch_matrix.NN4BEG0 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_1
X_1234_ net646 net631 net477 net417 Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
+ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_67_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1165_ _0282_ _0281_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__nand2b_1
X_1096_ _0219_ _0218_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR VPWR
+ _0220_ sky130_fd_sc_hd__mux2_1
XFILLER_52_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1998_ net754 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0949_ net75 net131 net103 Inst_LUT4AB_switch_matrix.JS2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_7_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1921_ net784 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1852_ net794 net666 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0803_ net67 net95 net24 net123 Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q
+ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux4_2
X_1783_ net742 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0734_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__inv_1
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2335_ Inst_LUT4AB_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_1
X_2266_ N4END[15] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__buf_1
XFILLER_69_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1217_ Inst_LUT4AB_switch_matrix.JN2BEG5 Inst_LUT4AB_switch_matrix.E2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__mux2_4
X_2197_ net792 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_1
XFILLER_25_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1148_ _0267_ _0254_ _0227_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_4
XFILLER_52_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1079_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 _0193_ _0194_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__o22a_1
XFILLER_40_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2120_ net768 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2051_ net779 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1002_ net654 net650 net625 net641 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__mux4_1
Xrebuffer19 Inst_LUT4AB_switch_matrix.E2BEG6 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1904_ net781 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1835_ net762 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1766_ net772 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0717_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__inv_2
X_1697_ net784 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2318_ S4END[15] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_2
X_2249_ net73 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_1
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput100 S2MID[1] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_2
Xinput111 SS4END[0] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xinput122 W2END[3] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_2
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput133 W2MID[6] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1620_ net749 net712 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
X_1551_ net802 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
X_1482_ net548 Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0529_ _0540_ _0541_ VGND
+ VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a32o_1
XFILLER_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2103_ net743 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ net752 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1818_ net798 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1749_ net746 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout801 net29 VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__buf_4
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0982_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0113_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q
+ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_57_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1603_ net778 net710 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1534_ net790 net700 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_1465_ _0165_ _0119_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR
+ _0525_ sky130_fd_sc_hd__mux2_1
X_1396_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q _0487_ _0486_ VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.EE4BEG2 sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_66_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2017_ net785 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold151 Inst_LB_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout642 D VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__clkbuf_2
Xfanout620 net432 VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__buf_8
Xfanout631 net632 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__buf_6
Xfanout653 net657 VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__buf_8
Xfanout675 net677 VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__clkbuf_2
Xfanout664 net58 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout697 net699 VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__clkbuf_2
Xfanout686 FrameStrobe[4] VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1250_ net464 net630 net478 net480 Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q
+ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__mux4_2
X_1181_ _0298_ _0299_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__nand2_1
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0965_ net74 net17 net102 net130 Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q
+ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__mux4_2
X_0896_ net634 net629 net620 net483 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__mux4_2
Xoutput201 net201 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput223 net223 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput234 net234 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput212 net212 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__buf_8
Xoutput256 net256 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput267 Inst_LUT4AB_switch_matrix.N4BEG2 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__buf_6
X_1517_ net757 net56 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
Xoutput278 net278 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput289 net289 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__buf_2
X_1448_ net411 Inst_LUT4AB_switch_matrix.E2BEG1 net658 _0255_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1379_ _0595_ _0029_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q VGND VGND VPWR VPWR
+ _0473_ sky130_fd_sc_hd__mux2_1
XFILLER_70_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0750_ net22 net93 net121 net140 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_24_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2351_ Inst_LUT4AB_switch_matrix.JW2BEG7 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__buf_1
X_1302_ net628 net619 net523 net416 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux4_1
X_2282_ NN4END[15] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__buf_1
X_1233_ _0347_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG7 sky130_fd_sc_hd__inv_4
XFILLER_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1164_ _0281_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__nand2b_1
X_1095_ net62 net70 net5 net13 Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux4_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1997_ net756 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0948_ _0081_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG5 sky130_fd_sc_hd__inv_2
XFILLER_9_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0879_ _0017_ _0014_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.E2BEG2 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_7_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1920_ net787 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1851_ net796 net665 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0802_ net80 net804 net136 Inst_LUT4AB_switch_matrix.JS2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_12_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1782_ net744 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0733_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__inv_1
XFILLER_69_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2334_ SS4END[15] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2265_ N4END[14] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_1
X_1216_ Inst_LUT4AB_switch_matrix.JS2BEG5 Inst_LUT4AB_switch_matrix.JW2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux2_4
X_2196_ net794 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_1
XFILLER_25_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1147_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0250_ _0239_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__mux4_1
X_1078_ _0201_ _0202_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q VGND VGND VPWR VPWR
+ _0203_ sky130_fd_sc_hd__mux2_4
XFILLER_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2050_ net783 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1001_ _0131_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR E sky130_fd_sc_hd__mux2_4
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1903_ net802 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1834_ net764 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1765_ net774 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0716_ net18 VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__inv_1
X_1696_ net787 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2317_ S4END[14] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_2
X_2248_ net72 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_4
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2179_ Inst_LUT4AB_switch_matrix.EE4BEG0 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_11_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 S2MID[2] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
Xinput123 W2END[4] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_2
Xinput134 W2MID[7] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput112 SS4END[1] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
XFILLER_48_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1550_ net755 net702 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
X_1481_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0529_ _0539_ Inst_LH_LUT4c_frame_config_dffesr.c_reset_value
+ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2102_ net744 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2033_ net759 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1817_ net800 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1748_ net748 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1679_ net802 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout802 net803 VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ net646 net630 net621 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux4_1
X_1602_ net782 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
X_1533_ net792 net702 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
X_1464_ _0264_ _0670_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q VGND VGND VPWR VPWR
+ _0524_ sky130_fd_sc_hd__mux2_1
X_1395_ net59 net87 net2 net651 Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q
+ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux4_1
XFILLER_67_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2016_ net787 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold152 Inst_LA_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout632 G VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__buf_6
Xfanout621 net622 VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__buf_4
Xfanout643 net645 VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__buf_2
Xfanout676 net677 VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__buf_1
Xfanout654 net656 VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__buf_2
XFILLER_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout665 net666 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkbuf_2
Xfanout687 FrameStrobe[3] VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__buf_2
Xfanout698 net699 VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__buf_2
XFILLER_73_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1180_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0283_ _0287_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__o22a_1
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0964_ net73 net101 net16 Inst_LUT4AB_switch_matrix.E2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__mux4_1
X_0895_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q _0031_ VGND VGND VPWR VPWR _0032_
+ sky130_fd_sc_hd__and2b_1
Xoutput224 net224 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput235 net235 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput202 net202 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput213 net213 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
X_1516_ net760 net56 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
Xoutput257 net257 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput246 net246 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__buf_4
Xoutput268 net268 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput279 net279 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
X_1447_ net412 _0640_ Inst_LUT4AB_switch_matrix.E2BEG2 _0624_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_67_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1378_ net632 net622 net482 net408 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_2_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2350_ Inst_LUT4AB_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_6
X_1301_ _0405_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q VGND VGND VPWR VPWR _0406_
+ sky130_fd_sc_hd__nand2b_4
X_2281_ NN4END[14] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_1
X_1232_ _0342_ _0340_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q _0346_ VGND VGND VPWR
+ VPWR _0347_ sky130_fd_sc_hd__a31o_1
XFILLER_49_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1163_ _0246_ _0247_ _0249_ _0248_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux4_2
X_1094_ net90 net116 net98 net659 Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q
+ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux4_1
XFILLER_52_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1996_ net761 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0947_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q _0080_ _0075_ _0077_ VGND VGND VPWR
+ VPWR _0081_ sky130_fd_sc_hd__a2bb2o_4
X_0878_ _0015_ _0016_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VGND VGND VPWR VPWR
+ _0017_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1850_ net798 net665 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1781_ net747 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_12_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0801_ _0644_ _0642_ _0647_ _0573_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG1
+ sky130_fd_sc_hd__a22o_4
X_0732_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__inv_1
X_2333_ SS4END[14] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_2
X_2264_ N4END[13] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_1
X_1215_ _0331_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop Inst_LD_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR D sky130_fd_sc_hd__mux2_4
X_2195_ net796 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_1
X_1146_ _0264_ _0265_ _0256_ _0255_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux4_2
XFILLER_25_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1077_ _0121_ _0120_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q VGND VGND VPWR VPWR
+ _0202_ sky130_fd_sc_hd__mux2_4
X_1979_ net797 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_48_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1000_ _0124_ _0110_ _0107_ _0127_ _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a32o_1
XFILLER_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1902_ net754 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1833_ net767 net663 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1764_ net777 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0715_ net75 VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__inv_1
X_1695_ net788 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2316_ S4END[13] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_2
X_2247_ net71 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2178_ EE4END[15] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1129_ _0246_ _0247_ _0249_ _0248_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q
+ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux4_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput102 S2MID[3] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
Xinput124 W2END[5] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xinput135 W6END[0] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_2
Xinput113 SS4END[2] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ _0289_ _0301_ _0539_ _0294_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__o211ai_1
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2101_ net746 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2032_ net780 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1816_ net54 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1747_ net750 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1678_ net755 net717 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout803 net28 VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0111_ VGND VGND VPWR VPWR _0112_
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1601_ net784 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
X_1532_ net794 net702 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1463_ _0287_ _0276_ _0286_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__a21bo_4
X_1394_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q _0485_ _0483_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q
+ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__o211a_1
XFILLER_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2015_ net35 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold153 Inst_LF_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout633 net634 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__buf_8
Xfanout622 H VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__clkbuf_4
Xfanout644 net645 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__buf_8
Xfanout666 net667 VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__clkbuf_2
Xfanout655 net656 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout677 net678 VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout688 FrameStrobe[3] VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout699 FrameStrobe[1] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0963_ _0090_ _0092_ _0095_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG5 sky130_fd_sc_hd__o22a_4
X_0894_ net653 net649 net639 net645 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__mux4_2
Xoutput225 net225 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput203 net203 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
Xoutput214 net214 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput236 net236 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
X_1515_ net762 net56 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
Xoutput258 net258 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput247 net247 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_6
Xoutput269 net269 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__buf_2
X_1446_ net804 net108 net93 net433 Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG0 sky130_fd_sc_hd__mux4_1
X_1377_ _0469_ _0470_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q VGND VGND VPWR VPWR
+ _0471_ sky130_fd_sc_hd__mux2_1
XFILLER_55_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1300_ _0639_ _0046_ _0082_ _0235_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux4_2
X_2280_ NN4END[13] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__buf_1
X_1231_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q _0345_ VGND VGND VPWR VPWR _0346_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_67_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1162_ _0235_ _0236_ _0238_ _0237_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux4_2
X_1093_ _0215_ _0216_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR VPWR
+ _0217_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_15_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ net763 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0946_ _0078_ _0079_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VGND VGND VPWR VPWR
+ _0080_ sky130_fd_sc_hd__mux2_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0877_ net804 net94 net122 net136 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_7_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1429_ net525 _0088_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q VGND VGND VPWR VPWR
+ _0516_ sky130_fd_sc_hd__mux2_1
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1780_ net748 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_12_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0800_ _0645_ _0646_ _0572_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__mux2_1
X_0731_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__inv_1
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2332_ SS4END[13] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2263_ N4END[12] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_1
X_1214_ _0324_ _0330_ _0320_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__mux2_4
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2194_ net798 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_1
X_1145_ net72 net15 net100 net128 Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q
+ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__mux4_1
XFILLER_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1076_ _0118_ _0119_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q VGND VGND VPWR VPWR
+ _0201_ sky130_fd_sc_hd__mux2_1
XFILLER_52_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1978_ net799 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0929_ net61 net69 net807 net12 Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux4_1
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1901_ net757 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1832_ net42 net663 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1763_ net779 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0714_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__inv_1
X_1694_ net790 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2315_ S4END[12] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_2
XFILLER_57_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2177_ EE4END[14] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1128_ net66 net111 net9 net122 Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q
+ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux4_2
XFILLER_15_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1059_ _0152_ _0184_ _0181_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__a21oi_1
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput125 W2END[6] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput136 W6END[1] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput103 S2MID[4] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput114 SS4END[3] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2100_ net748 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2031_ net802 net692 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1815_ net743 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1746_ net752 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1677_ net757 net717 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout804 net23 VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__buf_2
X_2229_ net719 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1600_ net787 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_1531_ net796 net702 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_26_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1462_ net463 Inst_LUT4AB_switch_matrix.JW2BEG3 _0165_ _0018_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG0
+ sky130_fd_sc_hd__mux4_2
X_1393_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__inv_1
XFILLER_67_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2014_ net791 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1729_ net784 net725 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xhold154 Inst_LH_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout623 net624 VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__buf_8
Xfanout634 net637 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__buf_8
Xfanout645 E VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__buf_8
Xfanout667 FrameStrobe[8] VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__buf_2
XFILLER_58_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout656 net657 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__buf_2
Xfanout678 FrameStrobe[6] VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__clkbuf_2
Xfanout689 FrameStrobe[3] VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__buf_2
XFILLER_73_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0962_ _0093_ _0094_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q VGND VGND VPWR VPWR
+ _0095_ sky130_fd_sc_hd__mux2_1
X_0893_ _0028_ _0029_ _0019_ _0018_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q
+ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__mux4_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput226 net226 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput215 net215 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
Xoutput204 net204 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput237 net237 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
X_1514_ net764 net56 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
Xoutput259 net259 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput248 net248 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__buf_8
XFILLER_4_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1445_ net805 net109 net94 net649 Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG1 sky130_fd_sc_hd__mux4_1
X_1376_ net627 net642 net647 net636 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux4_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1230_ _0343_ _0344_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q VGND VGND VPWR VPWR
+ _0345_ sky130_fd_sc_hd__mux2_1
X_1161_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux _0276_ _0279_ VGND VGND VPWR VPWR
+ _0280_ sky130_fd_sc_hd__a21oi_4
X_1092_ net646 net621 net477 net405 Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q
+ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_50_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1994_ net765 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0945_ net89 net115 net97 net660 Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__mux4_1
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0876_ net60 net82 net66 net9 Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q
+ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_7_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1428_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q _0638_ _0514_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__a211oi_1
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1359_ net62 net806 net659 net434 Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__mux4_1
XFILLER_55_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0730_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__inv_2
XFILLER_69_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2331_ SS4END[12] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_2
X_2262_ N4END[11] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_1
X_1213_ _0329_ _0326_ _0315_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__mux2_1
X_2193_ net800 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_1
X_1144_ net71 net14 net127 Inst_LUT4AB_switch_matrix.JW2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux4_1
XFILLER_25_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1075_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0198_ _0199_ _0195_
+ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_63_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1977_ net801 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0928_ _0061_ _0062_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VGND VGND VPWR VPWR
+ _0063_ sky130_fd_sc_hd__mux2_4
X_0859_ _0701_ _0700_ _0697_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__mux2_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1900_ net760 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1831_ net770 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1762_ net783 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0713_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__inv_1
X_1693_ net792 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2314_ S4END[11] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_2
X_2245_ Inst_LUT4AB_switch_matrix.JN2BEG6 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_1
X_2176_ EE4END[13] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_1
X_1127_ net81 net121 net113 Inst_LUT4AB_switch_matrix.E2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux4_2
XFILLER_65_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1058_ _0182_ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__nand2_1
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput126 W2END[7] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xinput115 W1END[0] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
Xinput104 S2MID[5] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
Xinput137 WW4END[0] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2030_ net754 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1814_ net53 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1745_ net759 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_15_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1676_ net761 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout805 net22 VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2228_ FrameStrobe[13] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2159_ E6END[6] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_1
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1530_ net798 net700 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
X_1461_ net641 _0068_ Inst_LUT4AB_switch_matrix.JW2BEG0 _0084_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG1
+ sky130_fd_sc_hd__mux4_1
X_1392_ net627 _0097_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q VGND VGND VPWR VPWR
+ _0484_ sky130_fd_sc_hd__mux2_1
XFILLER_67_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2013_ net793 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1728_ net786 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1659_ net796 net719 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
Xfanout624 C VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__buf_8
Xfanout657 A VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__buf_12
Xfanout635 net636 VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__buf_8
Xfanout646 net647 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__buf_2
Xfanout679 net681 VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__clkbuf_2
Xfanout668 FrameStrobe[8] VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__buf_2
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0961_ net87 net89 net97 net660 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__mux4_1
X_0892_ net74 net17 net102 net130 Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__mux4_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput216 net216 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
Xoutput205 net205 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput227 net227 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput238 net238 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
X_1513_ net766 net56 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
Xoutput249 net249 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__buf_6
X_1444_ net91 net136 net110 net414 Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1375_ net806 net659 net656 net651 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_53_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1160_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__inv_2
XFILLER_49_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1091_ net655 net650 net626 net641 Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_50_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1993_ net767 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0944_ net61 net69 net807 net12 Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux4_1
X_0875_ _0012_ _0013_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VGND VGND VPWR VPWR
+ _0014_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_7_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1427_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q net622 VGND VGND VPWR VPWR _0514_
+ sky130_fd_sc_hd__nor2_1
X_1358_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q _0452_ _0454_ VGND VGND VPWR VPWR
+ _0455_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1289_ net62 net64 net80 net25 Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux4_1
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2330_ SS4END[11] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
X_2261_ N4END[10] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_1
X_1212_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0050_ _0327_ _0328_
+ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__o211a_1
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2192_ net740 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_1
X_1143_ _0260_ _0258_ _0263_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JW2BEG6 sky130_fd_sc_hd__o22a_4
XFILLER_18_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1074_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 _0193_ _0196_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_63_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1976_ net741 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0927_ net646 net631 net621 net524 Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux4_2
X_0858_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ _0695_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux2_4
X_0789_ _0633_ _0632_ _0636_ _0570_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG3
+ sky130_fd_sc_hd__a22o_4
XFILLER_56_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1830_ net773 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1761_ net785 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0712_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__inv_1
X_1692_ net795 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2313_ S4END[10] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_2
X_2244_ Inst_LUT4AB_switch_matrix.JN2BEG5 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_2
X_2175_ EE4END[12] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
X_1126_ net74 net17 net102 net130 Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q
+ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__mux4_2
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1057_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0055_ _0153_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_23_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1959_ net771 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput116 W1END[1] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_4
Xinput127 W2MID[0] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xinput105 S2MID[6] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput138 WW4END[1] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XFILLER_71_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1813_ net747 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1744_ net780 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1675_ net763 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout806 net5 VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__clkbuf_4
X_2227_ FrameStrobe[12] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2158_ E6END[5] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2089_ net767 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ net62 net70 net806 net13 Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1460_ net464 Inst_LUT4AB_switch_matrix.JW2BEG1 net658 _0255_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_4_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1391_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q _0482_ VGND VGND VPWR VPWR _0483_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ net795 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1727_ net789 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1658_ net798 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
Xfanout658 _0247_ VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__buf_4
X_1589_ net747 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
Xfanout647 E VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__buf_2
Xfanout636 net637 VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__buf_8
XFILLER_58_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout625 net627 VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__buf_2
Xfanout669 net671 VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__buf_2
XFILLER_37_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0960_ net61 net69 net807 net12 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__mux4_1
XFILLER_40_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0891_ net73 net129 net16 Inst_LUT4AB_switch_matrix.E2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux4_1
Xoutput217 net217 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
Xoutput206 net206 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput228 net228 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput239 net239 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
X_1512_ net769 net56 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
X_1443_ net92 net107 net135 net445 Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1374_ _0465_ _0468_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.E6BEG1 sky130_fd_sc_hd__mux2_4
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1090_ _0050_ _0060_ _0105_ _0102_ _0197_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a311o_1
XFILLER_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1992_ net768 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_13_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0943_ _0076_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__a21boi_2
XFILLER_9_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0874_ net636 net630 net622 net402 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__mux4_1
X_1426_ net62 net806 net659 net656 Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__mux4_1
X_1357_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q _0638_ _0453_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_66_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1288_ net804 net120 net92 net136 Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
+ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux4_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2260_ N4END[9] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_1
X_1211_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0316_ _0317_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__o22a_1
X_2191_ net743 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_1
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1142_ _0261_ _0262_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VGND VGND VPWR VPWR
+ _0263_ sky130_fd_sc_hd__mux2_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1073_ _0190_ _0191_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_63_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1975_ net742 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0926_ net655 net650 net625 net640 Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__mux4_1
X_0857_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0695_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__mux2_4
X_0788_ _0634_ _0635_ _0569_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1409_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q _0498_ VGND VGND VPWR VPWR _0499_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1760_ net786 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0711_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__inv_2
X_1691_ net797 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2312_ S4END[9] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_2
X_2174_ EE4END[11] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
X_1125_ net73 net129 net101 net413 Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q
+ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_48_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1056_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0057_ _0155_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__o22a_1
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1958_ net772 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0909_ _0043_ _0044_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q VGND VGND VPWR VPWR
+ _0045_ sky130_fd_sc_hd__mux2_1
X_1889_ net784 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput117 W1END[2] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_2
Xinput106 S2MID[7] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
Xinput139 WW4END[2] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_2
Xinput128 W2MID[1] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1812_ net748 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1743_ net802 net730 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1674_ net765 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout807 net4 VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__buf_4
X_2226_ net731 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_36_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2157_ E6END[4] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_1
X_2088_ net768 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1108_ _0230_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a21bo_1
X_1039_ net653 net648 net444 net644 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux4_2
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1390_ net658 _0149_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q VGND VGND VPWR VPWR
+ _0482_ sky130_fd_sc_hd__mux2_1
XFILLER_67_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2011_ net797 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1726_ net791 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1657_ net800 net719 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_1588_ net749 net709 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
Xfanout648 net649 VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__buf_8
Xfanout637 F VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__buf_8
Xfanout626 net627 VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout659 net118 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2209_ net766 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_56_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0890_ net474 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG4 sky130_fd_sc_hd__inv_6
Xoutput207 net207 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput229 net229 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
X_1511_ net770 net56 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
Xoutput218 net218 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
X_1442_ net462 Inst_LUT4AB_switch_matrix.JS2BEG3 _0165_ _0018_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1373_ _0467_ _0466_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q VGND VGND VPWR VPWR
+ _0468_ sky130_fd_sc_hd__mux2_4
XFILLER_67_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1709_ net48 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_69_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1991_ net771 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0942_ net646 net631 net621 Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__mux4_2
XFILLER_9_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0873_ net656 net649 net639 net644 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__mux4_2
XFILLER_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1425_ _0510_ _0512_ _0508_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.NN4BEG2
+ sky130_fd_sc_hd__a21oi_1
X_1356_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q net412 VGND VGND VPWR VPWR _0453_
+ sky130_fd_sc_hd__nor2_1
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1287_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q _0393_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q
+ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_66_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1210_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0051_ VGND VGND
+ VPWR VPWR _0327_ sky130_fd_sc_hd__or2_1
X_2190_ net745 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_1
X_1141_ net88 net90 net98 net659 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__mux4_1
X_1072_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__inv_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1974_ net744 net686 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0925_ _0048_ _0030_ _0055_ _0058_ _0056_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a221o_1
X_0856_ _0696_ _0697_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__nor2_1
X_0787_ net67 net807 net10 net805 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__mux4_1
X_1408_ net61 net807 Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q VGND VGND VPWR VPWR
+ _0498_ sky130_fd_sc_hd__mux2_1
XFILLER_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1339_ net630 _0595_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _0439_ sky130_fd_sc_hd__mux2_1
XFILLER_71_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput390 net390 VGND VGND VPWR VPWR WW4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_59_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1690_ net799 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2311_ S4END[8] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_2
X_2242_ Inst_LUT4AB_switch_matrix.JN2BEG3 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__buf_1
X_2173_ EE4END[10] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1124_ _0245_ _0242_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.E2BEG6 sky130_fd_sc_hd__mux2_4
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1055_ _0179_ _0180_ _0152_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1957_ net774 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1888_ net786 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0908_ net88 net96 net116 net659 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux4_1
X_0839_ _0678_ _0679_ _0605_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__mux2_1
Xinput118 W1END[3] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
Xinput107 S4END[0] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
Xinput129 W2MID[2] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1811_ net750 net58 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1742_ net754 net725 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1673_ net767 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2225_ net734 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2156_ E6END[3] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2087_ net771 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ net646 net427 net635 net430 Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__mux4_2
X_1038_ net72 net15 net100 net128 Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q
+ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux4_2
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2010_ net799 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1725_ net793 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xhold147 Inst_LE_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ net740 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
X_1587_ net751 net710 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
Xfanout627 C VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__buf_8
Xfanout638 net639 VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__buf_8
Xfanout649 net652 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__buf_8
XFILLER_58_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2208_ net769 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_1
X_2139_ Inst_LUT4AB_switch_matrix.E2BEG0 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_6
XFILLER_66_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone70 net645 VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__buf_6
Xoutput208 net208 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput219 net219 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
X_1510_ net543 _0562_ _0560_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__mux2_1
X_1441_ net628 _0068_ Inst_LUT4AB_switch_matrix.JS2BEG0 _0084_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1372_ net630 net622 Inst_LUT4AB_switch_matrix.M_AD net416 Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux4_2
XFILLER_67_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1708_ net46 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1639_ net770 net714 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1990_ net772 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_15_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0941_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q _0074_ VGND VGND VPWR VPWR _0075_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_9_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0872_ _0011_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR B sky130_fd_sc_hd__mux2_4
XFILLER_9_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1424_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q _0511_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q
+ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__a21oi_1
X_1355_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q _0451_ VGND VGND VPWR VPWR _0452_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_50_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1286_ net446 net444 net463 net643 Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q
+ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_66_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1140_ net62 net70 net806 net13 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__mux4_1
XFILLER_37_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1071_ _0190_ _0191_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__nand2_1
XFILLER_18_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1973_ net746 net686 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0924_ _0058_ _0055_ _0056_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a21o_1
X_0855_ _0696_ _0697_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__nand2_1
X_0786_ net95 net123 net107 net139 Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q
+ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__mux4_1
X_1407_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q _0496_ _0494_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q
+ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__o211a_1
X_1338_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q _0437_ VGND VGND VPWR VPWR _0438_
+ sky130_fd_sc_hd__nand2_1
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1269_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q _0377_ VGND VGND VPWR VPWR _0378_
+ sky130_fd_sc_hd__or2_1
XFILLER_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput380 net380 VGND VGND VPWR VPWR WW4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput391 net391 VGND VGND VPWR VPWR WW4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2310_ S4END[7] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_2
X_2241_ Inst_LUT4AB_switch_matrix.JN2BEG2 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_6
X_2172_ EE4END[9] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1123_ _0244_ _0243_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VGND VGND VPWR VPWR
+ _0245_ sky130_fd_sc_hd__mux2_1
X_1054_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0057_ _0155_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__o22a_1
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1956_ net777 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0907_ net60 net68 net3 net11 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux4_1
X_1887_ net789 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0838_ _0681_ _0680_ _0605_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__mux2_1
X_0769_ net434 net638 net624 net644 Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__mux4_1
Xinput108 S4END[1] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
Xinput119 W2END[0] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_39_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1810_ net752 net58 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_70_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1741_ net756 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1672_ net768 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2224_ net664 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__buf_1
X_2155_ E6END[2] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_1
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1106_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q _0228_ VGND VGND VPWR VPWR _0229_
+ sky130_fd_sc_hd__and2b_1
X_2086_ net772 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1037_ net71 net99 net127 net479 Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q
+ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux4_1
XFILLER_53_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_1_0__leaf_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1939_ net750 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput90 S1END[3] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1724_ net795 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold148 Inst_LD_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ net743 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
X_1586_ net752 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
Xfanout628 net629 VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__buf_6
Xfanout639 D VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_8
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout617 net431 VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__buf_8
XFILLER_58_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2207_ net770 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_1
XFILLER_73_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2069_ net746 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput209 net209 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
X_1440_ net619 Inst_LUT4AB_switch_matrix.JS2BEG1 net658 _0255_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1371_ _0639_ _0046_ _0082_ _0235_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux4_1
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1707_ net762 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1638_ net773 net714 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_1569_ net784 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_69_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0940_ net654 net650 net626 net640 Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux4_1
X_0871_ _0706_ _0010_ _0688_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__mux2_4
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1423_ net115 net651 Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q VGND VGND VPWR VPWR
+ _0511_ sky130_fd_sc_hd__mux2_1
X_1354_ net525 _0121_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q VGND VGND VPWR VPWR
+ _0451_ sky130_fd_sc_hd__mux2_1
X_1285_ _0580_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__or2_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1070_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0194_ VGND VGND
+ VPWR VPWR _0195_ sky130_fd_sc_hd__or2_1
XFILLER_18_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1972_ net749 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0923_ _0692_ _0693_ _0698_ _0699_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a31oi_4
X_0854_ _0594_ _0595_ _0604_ _0603_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q
+ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux4_2
X_0785_ _0630_ _0569_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0633_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2386_ Inst_LUT4AB_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__buf_1
X_1406_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__inv_1
X_1337_ _0029_ _0238_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _0437_ sky130_fd_sc_hd__mux2_1
XFILLER_68_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1268_ net648 net638 net623 net643 Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1199_ _0030_ _0049_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nand2_1
XFILLER_36_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput370 net370 VGND VGND VPWR VPWR W6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput392 net392 VGND VGND VPWR VPWR WW4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput381 net381 VGND VGND VPWR VPWR WW4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_59_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2240_ Inst_LUT4AB_switch_matrix.JN2BEG1 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__buf_2
X_2171_ EE4END[8] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1122_ net62 net70 net806 net13 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux4_1
X_1053_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0055_ _0153_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__o22a_1
XFILLER_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1955_ net779 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0906_ _0040_ _0041_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q VGND VGND VPWR VPWR
+ _0042_ sky130_fd_sc_hd__mux2_4
X_1886_ net791 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0837_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ _0628_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__mux2_1
X_0768_ net634 net629 net620 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__mux4_2
Xinput109 S4END[2] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
X_2369_ W6END[11] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_39_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1740_ net761 net725 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1671_ net771 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2223_ net665 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2154_ net21 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1105_ net657 net651 net626 net640 Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__mux4_1
X_2085_ net774 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1036_ _0163_ _0160_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.JW2BEG4 sky130_fd_sc_hd__mux2_4
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1938_ net752 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1869_ net756 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput80 N4END[1] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
Xinput91 S2END[0] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_10_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1723_ net797 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
Xhold149 Inst_LG_LUT4c_frame_config_dffesr.LUT_flop VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ net745 net719 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
X_1585_ net758 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
Xfanout618 net480 VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__buf_12
Xfanout629 G VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_8
X_2206_ net773 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_1
X_2068_ net748 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1019_ _0144_ _0142_ _0147_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JN2BEG2 sky130_fd_sc_hd__o22a_4
XFILLER_53_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone50 net639 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__buf_6
Xclone83 net637 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1370_ _0464_ _0463_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q VGND VGND VPWR VPWR
+ _0465_ sky130_fd_sc_hd__mux2_1
XFILLER_67_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1706_ net765 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1637_ net775 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
X_1568_ net787 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1499_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q _0529_ VGND VGND VPWR VPWR _0554_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0870_ _0009_ _0709_ _0696_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__mux2_1
XFILLER_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1422_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q _0509_ VGND VGND VPWR VPWR _0510_
+ sky130_fd_sc_hd__nand2b_1
X_1353_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q _0450_ _0449_ VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.SS4BEG2 sky130_fd_sc_hd__o21ba_1
X_1284_ net634 net629 net619 net416 Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__mux4_2
XFILLER_51_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0999_ _0073_ _0129_ _0124_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_6_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout790 net791 VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1971_ net751 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0922_ _0052_ _0053_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__nand2_1
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0853_ _0639_ _0640_ _0649_ _0648_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q
+ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__mux4_2
X_0784_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q _0631_ VGND VGND VPWR VPWR _0632_
+ sky130_fd_sc_hd__or2_4
X_1405_ net632 _0595_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q VGND VGND VPWR VPWR
+ _0495_ sky130_fd_sc_hd__mux2_1
X_1336_ _0435_ _0436_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.WW4BEG1 sky130_fd_sc_hd__mux2_4
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput1 Ci VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_12
XFILLER_28_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1267_ net650 net654 net520 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.M_AB sky130_fd_sc_hd__mux2_4
X_1198_ _0314_ _0059_ Inst_LD_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0315_ sky130_fd_sc_hd__mux2_4
XFILLER_24_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput360 net360 VGND VGND VPWR VPWR W2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput371 net371 VGND VGND VPWR VPWR W6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput393 net393 VGND VGND VPWR VPWR WW4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput382 Inst_LUT4AB_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR WW4BEG[12] sky130_fd_sc_hd__buf_6
XFILLER_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_29_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2170_ EE4END[7] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
X_1121_ net88 net90 net98 net659 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__mux4_1
X_1052_ _0177_ _0157_ _0152_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
XFILLER_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1954_ net783 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0905_ net635 net630 net621 net403 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__mux4_2
X_1885_ net793 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0836_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ _0628_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__mux2_1
X_0767_ _0613_ _0614_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q VGND VGND VPWR VPWR
+ _0616_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_47_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2368_ W6END[10] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__buf_4
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2299_ net99 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_39_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1319_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q _0422_ VGND VGND VPWR VPWR _0423_
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_56_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput190 net190 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK VGND VGND VPWR VPWR clknet_1_0__leaf_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1670_ net772 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2222_ net672 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_1
XFILLER_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2153_ net20 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_1
X_1104_ _0214_ _0198_ Inst_LG_LUT4c_frame_config_dffesr.c_I0mux _0226_ VGND VGND VPWR
+ VPWR _0227_ sky130_fd_sc_hd__a31o_1
XFILLER_53_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2084_ net777 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1035_ _0161_ _0162_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VGND VGND VPWR VPWR
+ _0163_ sky130_fd_sc_hd__mux2_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1937_ net758 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1868_ net760 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput81 N4END[2] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
Xinput70 N2END[7] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
X_0819_ net462 net628 net619 net618 Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__mux4_1
X_1799_ net41 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput92 S2END[1] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1722_ net799 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1653_ net747 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1584_ net781 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
Xfanout619 net620 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__buf_6
X_2205_ net775 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2136_ Inst_LUT4AB_switch_matrix.E1BEG1 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__buf_4
X_2067_ net750 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1018_ _0145_ _0146_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q VGND VGND VPWR VPWR
+ _0147_ sky130_fd_sc_hd__mux2_1
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone40 A VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_1
Xclone51 D VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_1
Xclone84 net636 VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_6
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1705_ net767 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1636_ net776 net714 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
X_1567_ net788 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_1498_ net542 _0553_ _0551_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__mux2_1
XFILLER_39_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ net771 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1421_ net59 net2 Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q VGND VGND VPWR VPWR _0509_
+ sky130_fd_sc_hd__mux2_1
X_1352_ net59 net115 net2 net649 Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
+ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__mux4_1
X_1283_ _0386_ _0387_ _0390_ _0579_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0998_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0104_ _0105_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0128_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__o221a_1
X_1619_ net751 net712 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout780 net781 VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__buf_2
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout791 net34 VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__buf_4
XFILLER_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1970_ net753 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0921_ _0052_ _0053_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__and2_1
X_0852_ _0691_ _0694_ Inst_LB_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0695_ sky130_fd_sc_hd__mux2_4
X_0783_ net653 net648 net623 net643 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__mux4_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1404_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q _0493_ VGND VGND VPWR VPWR _0494_
+ sky130_fd_sc_hd__nand2_1
X_1335_ net621 _0639_ _0046_ _0085_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__mux4_2
Xinput2 E1END[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1266_ _0375_ _0376_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.M_AH sky130_fd_sc_hd__mux2_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1197_ _0313_ _0312_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q VGND VGND VPWR VPWR
+ _0314_ sky130_fd_sc_hd__mux2_1
XFILLER_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput361 net361 VGND VGND VPWR VPWR W2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput350 net350 VGND VGND VPWR VPWR W1BEG[3] sky130_fd_sc_hd__buf_8
Xoutput394 net394 VGND VGND VPWR VPWR WW4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput383 Inst_LUT4AB_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR WW4BEG[13] sky130_fd_sc_hd__buf_8
Xoutput372 net372 VGND VGND VPWR VPWR W6BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1120_ _0240_ _0241_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VGND VGND VPWR VPWR
+ _0242_ sky130_fd_sc_hd__mux2_4
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1051_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0055_ _0175_ _0176_
+ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__o211a_1
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1953_ net785 net57 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0904_ net654 net650 net625 net641 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__mux4_1
X_1884_ net32 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0835_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0628_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0766_ _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__inv_1
X_2367_ W6END[9] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_39_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2298_ Inst_LUT4AB_switch_matrix.JS2BEG7 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__buf_6
X_1318_ _0595_ _0029_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q VGND VGND VPWR VPWR
+ _0422_ sky130_fd_sc_hd__mux2_1
X_1249_ net654 net649 net624 net638 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__mux4_2
XFILLER_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput180 Inst_LUT4AB_switch_matrix.EE4BEG3 VGND VGND VPWR VPWR EE4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput191 net191 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2221_ net676 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_2
X_2152_ net19 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_1
X_1103_ Inst_LG_LUT4c_frame_config_dffesr.c_I0mux _0225_ VGND VGND VPWR VPWR _0226_
+ sky130_fd_sc_hd__and2b_1
X_2083_ net779 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1034_ net88 net96 net90 net116 Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
+ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__mux4_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1936_ net780 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1867_ net762 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput82 N4END[3] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
Xinput60 N1END[1] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_4
Xinput71 N2MID[0] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlymetal6s2s_1
X_0818_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0662_ VGND VGND VPWR VPWR _0663_
+ sky130_fd_sc_hd__and2b_1
X_1798_ net773 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput93 S2END[2] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
X_0749_ net59 net65 net81 net8 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__mux4_1
XFILLER_69_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ net801 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1652_ net749 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
X_1583_ net803 net709 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2204_ net776 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_1
X_2135_ Inst_LUT4AB_switch_matrix.E1BEG0 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_1
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2066_ net752 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1017_ net804 net94 net122 net138 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux4_1
X_1919_ net788 net677 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone52 net649 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1704_ net768 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1635_ net778 net714 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
X_1566_ net790 net705 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1497_ Inst_LD_LUT4c_frame_config_dffesr.c_reset_value _0331_ _0552_ VGND VGND VPWR
+ VPWR _0553_ sky130_fd_sc_hd__mux2_2
XFILLER_39_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2118_ net772 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ net785 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1420_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q _0507_ _0505_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q
+ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__o211a_1
X_1351_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q _0448_ _0446_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q
+ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__o211a_1
X_1282_ _0388_ _0389_ _0578_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
XFILLER_48_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0997_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0100_ _0101_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__o22a_1
X_1618_ net753 net712 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
X_1549_ net757 net703 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_regs_0_UserCLK UserCLK VGND VGND VPWR VPWR UserCLK_regs sky130_fd_sc_hd__clkbuf_16
Xfanout770 net41 VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__buf_4
Xfanout781 net38 VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__buf_4
Xfanout792 net793 VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ _0052_ _0053_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__or2_2
XFILLER_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0851_ _0693_ _0692_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__nand2_2
X_0782_ net633 net628 net619 net523 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__mux4_2
XFILLER_5_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2383_ WW4END[15] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1403_ _0029_ _0224_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q VGND VGND VPWR VPWR
+ _0493_ sky130_fd_sc_hd__mux2_1
X_1334_ net62 net90 net118 net654 Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__mux4_1
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1265_ _0374_ _0338_ _0370_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux2_1
Xinput3 E1END[1] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1196_ _0138_ _0139_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q VGND VGND VPWR VPWR
+ _0313_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput362 net362 VGND VGND VPWR VPWR W2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput351 net351 VGND VGND VPWR VPWR W2BEG[0] sky130_fd_sc_hd__buf_4
Xoutput340 net340 VGND VGND VPWR VPWR SS4BEG[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput384 net384 VGND VGND VPWR VPWR WW4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput373 net373 VGND VGND VPWR VPWR W6BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0155_ VGND VGND
+ VPWR VPWR _0176_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1952_ net786 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0903_ net67 net10 net113 net123 Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q
+ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux4_2
X_1883_ net31 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0834_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0628_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0765_ net78 net21 net106 net134 Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q
+ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__mux4_2
X_2366_ W6END[8] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_2
X_1317_ net631 net622 net482 net406 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux4_2
X_1248_ _0360_ _0357_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.JS2BEG7 sky130_fd_sc_hd__mux2_4
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1179_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0284_ _0286_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__o22a_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput170 net170 VGND VGND VPWR VPWR E6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput181 net181 VGND VGND VPWR VPWR EE4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput192 net192 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2220_ net682 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_2
X_2151_ net18 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_1
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1102_ _0221_ _0222_ _0224_ _0223_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__mux4_2
X_2082_ net783 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1033_ net60 net68 net3 net11 Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__mux4_1
XFILLER_53_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1935_ net803 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1866_ net764 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput61 N1END[2] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_4
X_0817_ net433 net648 net463 net643 Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__mux4_2
Xinput72 N2MID[1] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
X_1797_ net775 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput50 FrameData[3] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
X_0748_ _0565_ _0598_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _0599_ sky130_fd_sc_hd__o21a_1
Xinput83 NN4END[0] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 S2END[3] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
X_2349_ Inst_LUT4AB_switch_matrix.JW2BEG5 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__buf_1
XFILLER_69_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1720_ net741 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1651_ net751 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
X_1582_ net49 net707 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
X_2203_ net778 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2134_ clknet_1_1__leaf_UserCLK_regs _0007_ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2065_ net759 net696 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1016_ net66 net82 net3 net9 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_14_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1918_ net790 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1849_ net29 net665 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone20 C VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1703_ net770 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1634_ net782 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
X_1565_ net792 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1496_ _0538_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q VGND VGND VPWR VPWR _0552_
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2117_ net774 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2048_ net786 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1350_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__inv_1
X_1281_ net84 net7 net806 net804 Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__mux4_1
XFILLER_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0996_ _0125_ _0126_ _0073_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1617_ net47 net712 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
X_1548_ net760 net700 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1479_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q _0538_ VGND VGND VPWR VPWR _0539_
+ sky130_fd_sc_hd__nand2_2
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_UserCLK_regs UserCLK_regs VGND VGND VPWR VPWR clknet_0_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_17_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout760 net761 VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__clkbuf_4
Xfanout793 net33 VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__buf_4
Xfanout771 net41 VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__buf_4
Xfanout782 net783 VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__buf_4
XFILLER_18_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0850_ _0605_ net1 VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__nand2_8
X_0781_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__mux2_1
XFILLER_5_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1402_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q _0488_ _0490_ _0492_ VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.EE4BEG1 sky130_fd_sc_hd__o22a_4
X_2382_ WW4END[14] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_2
X_1333_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q _0434_ _0433_ VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.WW4BEG2 sky130_fd_sc_hd__o21ba_1
X_1264_ _0373_ _0374_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ _0375_ sky130_fd_sc_hd__mux2_4
XFILLER_68_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 E1END[2] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1195_ _0149_ _0148_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q VGND VGND VPWR VPWR
+ _0312_ sky130_fd_sc_hd__mux2_1
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0979_ net654 net650 net625 net640 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux4_1
Xoutput352 net352 VGND VGND VPWR VPWR W2BEG[1] sky130_fd_sc_hd__buf_8
Xoutput330 net330 VGND VGND VPWR VPWR SS4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput341 net341 VGND VGND VPWR VPWR SS4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput363 net363 VGND VGND VPWR VPWR W2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput385 Inst_LUT4AB_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR WW4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput374 net374 VGND VGND VPWR VPWR W6BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_59_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1951_ net789 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0902_ net84 net25 net108 Inst_LUT4AB_switch_matrix.JS2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__mux4_2
X_1882_ net799 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0833_ _0676_ _0652_ _0650_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__mux2_4
X_0764_ net77 net105 net133 Inst_LUT4AB_switch_matrix.JN2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__mux4_1
X_2365_ W6END[7] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_2
X_1316_ _0418_ _0419_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q VGND VGND VPWR VPWR
+ _0420_ sky130_fd_sc_hd__mux2_1
X_2296_ Inst_LUT4AB_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_2
X_1247_ _0358_ _0359_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VGND VGND VPWR VPWR
+ _0360_ sky130_fd_sc_hd__mux2_1
X_1178_ _0295_ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__nand2_1
XFILLER_64_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput160 net160 VGND VGND VPWR VPWR E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput182 net182 VGND VGND VPWR VPWR EE4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput171 net171 VGND VGND VPWR VPWR E6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput193 net193 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2150_ net17 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_1
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1101_ net70 net13 net98 net137 Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q
+ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__mux4_2
X_2081_ net785 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1032_ _0158_ _0159_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VGND VGND VPWR VPWR
+ _0160_ sky130_fd_sc_hd__mux2_4
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1934_ net754 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1865_ net766 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput40 FrameData[21] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
X_1796_ net776 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput62 N1END[3] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_4
Xinput73 N2MID[2] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
X_0816_ net63 net91 net6 net140 Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q
+ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__mux4_2
Xinput51 FrameData[4] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
X_0747_ net415 net629 net620 net618 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__mux4_1
Xinput84 NN4END[1] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
Xinput95 S2END[4] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
X_2348_ net479 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__buf_6
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2279_ NN4END[12] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1650_ net753 net719 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_1581_ net48 net707 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_2202_ net782 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_1
X_2133_ clknet_1_1__leaf_UserCLK_regs _0006_ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
X_2064_ net780 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_34_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1015_ _0143_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q
+ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1917_ net33 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1848_ net740 net665 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1779_ net750 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_4_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone21 net637 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1702_ net773 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1633_ net784 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
X_1564_ net794 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
X_1495_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q _0529_ VGND VGND VPWR VPWR _0551_
+ sky130_fd_sc_hd__nand2_1
X_2116_ net777 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2047_ net789 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1280_ net92 net120 net108 net136 Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux4_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0995_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0104_ _0105_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__o22a_1
X_1616_ net38 net712 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1547_ net762 net702 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1478_ _0537_ _0535_ _0533_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__o21a_4
XFILLER_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout750 net751 VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__clkbuf_4
Xfanout794 net795 VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__clkbuf_4
Xfanout772 FrameData[23] VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__clkbuf_4
Xfanout783 net37 VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__clkbuf_4
Xfanout761 net46 VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__clkbuf_8
XFILLER_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0780_ _0627_ net1 Inst_LA_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0628_ sky130_fd_sc_hd__mux2_4
XFILLER_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1401_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q _0491_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q
+ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a21bo_1
X_2381_ WW4END[13] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1332_ net59 net115 net87 net446 Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
+ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__mux4_1
X_1263_ _0373_ net617 _0371_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux2_4
Xinput5 E1END[3] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1194_ net484 net646 _0311_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.M_EF sky130_fd_sc_hd__mux2_4
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0978_ _0108_ _0109_ _0073_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__a21o_1
Xoutput353 net353 VGND VGND VPWR VPWR W2BEG[2] sky130_fd_sc_hd__buf_4
Xoutput320 net320 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR SS4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput342 net342 VGND VGND VPWR VPWR SS4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput364 net364 VGND VGND VPWR VPWR W2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput386 net386 VGND VGND VPWR VPWR WW4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput375 net375 VGND VGND VPWR VPWR W6BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1950_ net791 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0901_ _0034_ _0032_ _0037_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JS2BEG2 sky130_fd_sc_hd__o22a_4
X_1881_ net801 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0832_ _0674_ _0675_ _0605_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__mux2_1
X_0763_ _0608_ _0609_ _0612_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JN2BEG3 sky130_fd_sc_hd__o22a_4
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2364_ W6END[6] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_2
X_1315_ net626 net640 net646 net636 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux4_1
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2295_ net526 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__buf_6
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1246_ net87 net115 net91 net117 Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q
+ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux4_1
X_1177_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0283_ _0287_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_22_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput150 net150 VGND VGND VPWR VPWR E2BEG[4] sky130_fd_sc_hd__buf_8
Xoutput161 net161 VGND VGND VPWR VPWR E2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput183 net183 VGND VGND VPWR VPWR EE4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput172 net172 VGND VGND VPWR VPWR E6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput194 net194 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1100_ net82 net24 net110 Inst_LUT4AB_switch_matrix.JN2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__mux4_1
X_2080_ net786 net699 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_36_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1031_ net478 net630 net621 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux4_2
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1933_ net756 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput30 FrameData[11] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
X_1864_ net768 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1795_ net778 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0815_ net79 net22 net107 Inst_LUT4AB_switch_matrix.JW2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__mux4_1
Xinput63 N2END[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xinput52 FrameData[5] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
Xinput41 FrameData[24] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
X_0746_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q _0596_ VGND VGND VPWR VPWR _0597_
+ sky130_fd_sc_hd__or2_1
Xinput74 N2MID[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
Xinput85 NN4END[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput96 S2END[5] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
X_2347_ Inst_LUT4AB_switch_matrix.JW2BEG3 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__buf_6
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2278_ NN4END[11] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_1
X_1229_ net87 net89 net111 net137 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__mux4_1
XFILLER_52_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1580_ net761 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2201_ net784 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
X_2132_ clknet_1_1__leaf_UserCLK_regs _0005_ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_53_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2063_ net802 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1014_ net637 net630 net622 net407 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__mux4_2
X_1916_ net794 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_62_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1847_ net743 net665 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1778_ net752 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0729_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_71_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1701_ net775 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1632_ net787 net715 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
X_1563_ net796 net705 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
X_1494_ net544 _0550_ _0548_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__mux2_1
XFILLER_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2115_ net779 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2046_ net791 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0100_ _0101_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__o22a_1
X_1615_ net803 net712 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
X_1546_ net764 net700 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1477_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q _0536_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q
+ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__a21bo_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2029_ net756 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout740 net741 VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__clkbuf_4
Xfanout751 net51 VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__buf_4
Xfanout762 net763 VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__clkbuf_4
Xfanout773 FrameData[23] VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__clkbuf_4
Xfanout784 net785 VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__buf_4
XFILLER_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout795 net32 VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1400_ net525 _0070_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q VGND VGND VPWR VPWR
+ _0491_ sky130_fd_sc_hd__mux2_1
X_2380_ WW4END[12] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_2
X_1331_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q _0432_ _0430_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q
+ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__o211a_1
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1262_ net622 net631 _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__mux2_1
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 E2END[0] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
X_1193_ _0306_ net475 Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VGND VGND VPWR VPWR
+ _0311_ sky130_fd_sc_hd__mux2_4
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0977_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 _0100_ _0105_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__o22a_1
Xoutput310 net310 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__buf_2
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 net321 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput343 net343 VGND VGND VPWR VPWR SS4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput332 net332 VGND VGND VPWR VPWR SS4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput387 net387 VGND VGND VPWR VPWR WW4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput365 net365 VGND VGND VPWR VPWR W2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput354 net354 VGND VGND VPWR VPWR W2BEG[3] sky130_fd_sc_hd__buf_8
Xoutput376 net376 VGND VGND VPWR VPWR W6BEG[7] sky130_fd_sc_hd__buf_2
X_1529_ net800 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0036_ _0035_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q VGND VGND VPWR VPWR
+ _0037_ sky130_fd_sc_hd__mux2_1
X_1880_ net741 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0831_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ _0628_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__mux2_1
X_0762_ _0610_ _0611_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q VGND VGND VPWR VPWR
+ _0612_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2363_ W6END[5] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_2
X_1314_ net806 net659 net654 net651 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux4_1
X_2294_ Inst_LUT4AB_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1245_ net59 net63 net2 net6 Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux4_1
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1176_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0284_ _0286_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__o22a_1
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_1_1__leaf_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput151 net151 VGND VGND VPWR VPWR E2BEG[5] sky130_fd_sc_hd__buf_6
Xoutput184 net184 VGND VGND VPWR VPWR EE4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput162 net162 VGND VGND VPWR VPWR E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput173 net173 VGND VGND VPWR VPWR E6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput195 net195 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ net654 net650 net625 net641 Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux4_1
XFILLER_61_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1932_ net761 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_61_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1863_ net771 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0814_ _0656_ _0654_ _0659_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JW2BEG1 sky130_fd_sc_hd__o22a_4
Xinput20 E2MID[6] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
Xinput31 FrameData[12] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
X_1794_ net782 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput64 N2END[1] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 FrameData[7] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
Xinput42 FrameData[25] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xinput86 NN4END[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput75 N2MID[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
X_0745_ net433 net639 net624 net645 Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__mux4_1
Xinput97 S2END[6] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2346_ Inst_LUT4AB_switch_matrix.JW2BEG2 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_1
XFILLER_69_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2277_ NN4END[10] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1228_ net59 net63 net2 net6 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__mux4_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1159_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux _0277_ VGND VGND VPWR VPWR _0278_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2200_ net787 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
X_2131_ clknet_1_0__leaf_UserCLK_regs _0004_ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2062_ net754 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1013_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q _0141_ VGND VGND VPWR VPWR _0142_
+ sky130_fd_sc_hd__and2b_1
XFILLER_19_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1915_ net796 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1846_ net745 net666 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1777_ net759 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0728_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2329_ SS4END[10] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_2
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1700_ net776 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1631_ net788 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_1562_ net798 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_1493_ Inst_LC_LUT4c_frame_config_dffesr.c_reset_value _0186_ _0549_ VGND VGND VPWR
+ VPWR _0550_ sky130_fd_sc_hd__mux2_2
XFILLER_39_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2114_ net783 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2045_ net793 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1829_ net775 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0993_ _0122_ _0123_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q VGND VGND VPWR VPWR
+ _0124_ sky130_fd_sc_hd__mux2_4
XFILLER_8_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1614_ net49 net710 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
X_1545_ net766 net700 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1476_ Inst_LUT4AB_switch_matrix.JS2BEG1 Inst_LUT4AB_switch_matrix.JW2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__mux2_1
XFILLER_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2028_ net761 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout741 net54 VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__buf_4
Xfanout730 net731 VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkbuf_2
Xfanout752 net753 VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__clkbuf_4
Xfanout785 net36 VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__clkbuf_4
Xfanout774 FrameData[22] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__clkbuf_4
Xfanout763 net45 VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__clkbuf_8
Xfanout796 net797 VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__clkbuf_4
XFILLER_65_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1330_ _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__inv_1
X_1261_ _0371_ _0311_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ _0372_ sky130_fd_sc_hd__mux2_1
Xinput7 E2END[1] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
X_1192_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q _0309_ _0308_ VGND VGND VPWR VPWR
+ _0310_ sky130_fd_sc_hd__a21oi_4
XFILLER_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0976_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0101_ _0104_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__o22a_1
Xoutput300 net300 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__buf_8
Xoutput311 net311 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput322 net322 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput333 net333 VGND VGND VPWR VPWR SS4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput344 net344 VGND VGND VPWR VPWR SS4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput366 net366 VGND VGND VPWR VPWR W2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput355 net355 VGND VGND VPWR VPWR W2BEG[4] sky130_fd_sc_hd__buf_8
Xoutput377 net377 VGND VGND VPWR VPWR W6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput388 net388 VGND VGND VPWR VPWR WW4BEG[3] sky130_fd_sc_hd__buf_2
X_1528_ net740 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1459_ net637 _0640_ Inst_LUT4AB_switch_matrix.JW2BEG2 _0624_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0830_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0628_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__mux2_1
X_0761_ net805 net95 net123 net135 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__mux4_1
X_2362_ W6END[4] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_2
X_2293_ Inst_LUT4AB_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_6
X_1313_ _0584_ _0412_ _0417_ _0408_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W6BEG1
+ sky130_fd_sc_hd__a31o_1
X_1244_ _0355_ _0356_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VGND VGND VPWR VPWR
+ _0357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1175_ _0280_ _0288_ _0289_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__o211ai_2
XFILLER_64_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0959_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0091_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__a21bo_1
Xoutput152 net152 VGND VGND VPWR VPWR E2BEG[6] sky130_fd_sc_hd__buf_6
Xoutput141 net141 VGND VGND VPWR VPWR Co sky130_fd_sc_hd__buf_8
Xoutput174 net174 VGND VGND VPWR VPWR EE4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput185 net185 VGND VGND VPWR VPWR EE4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput163 Inst_LUT4AB_switch_matrix.E6BEG0 VGND VGND VPWR VPWR E6BEG[10] sky130_fd_sc_hd__buf_6
Xoutput196 net196 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1931_ net763 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1862_ net772 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0813_ _0657_ _0658_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q VGND VGND VPWR VPWR
+ _0659_ sky130_fd_sc_hd__mux2_1
Xinput21 E2MID[7] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput10 E2END[4] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
X_1793_ net785 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput54 FrameData[9] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
Xinput32 FrameData[13] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 FrameData[26] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
X_0744_ net74 net17 net102 net130 Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q
+ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__mux4_2
Xinput76 N2MID[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput65 N2END[2] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput87 S1END[0] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xinput98 S2END[7] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
X_2345_ Inst_LUT4AB_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__buf_6
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2276_ NN4END[9] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_1
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1227_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0341_ VGND VGND VPWR VPWR _0342_
+ sky130_fd_sc_hd__nand2_1
XFILLER_52_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1158_ _0221_ _0222_ _0224_ _0223_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__mux4_1
X_1089_ _0213_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop Inst_LF_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR F sky130_fd_sc_hd__mux2_4
XFILLER_4_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2130_ clknet_1_0__leaf_UserCLK_regs _0003_ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2061_ net756 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1012_ net656 net651 net642 net647 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__mux4_1
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1914_ net798 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1845_ net747 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1776_ net780 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0727_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__inv_1
X_2328_ SS4END[9] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_2
XFILLER_57_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2259_ N4END[8] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone68 net634 VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1630_ net790 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_1561_ net800 net705 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
X_1492_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q _0538_ VGND VGND VPWR VPWR _0549_
+ sky130_fd_sc_hd__nand2_2
XFILLER_66_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2113_ net36 net739 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2044_ net795 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1828_ net776 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_9_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1759_ net789 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0992_ _0121_ _0120_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q VGND VGND VPWR VPWR
+ _0123_ sky130_fd_sc_hd__mux2_4
X_1613_ net757 net710 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
X_1544_ net769 net700 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
X_1475_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q _0534_ VGND VGND VPWR VPWR _0535_
+ sky130_fd_sc_hd__and2b_1
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2027_ net763 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout720 net721 VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__buf_2
Xfanout742 FrameData[8] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__buf_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout731 FrameStrobe[11] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__buf_2
Xfanout764 net765 VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__clkbuf_4
Xfanout753 net50 VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__buf_4
Xfanout775 FrameData[22] VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__buf_4
Xfanout797 net31 VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__clkbuf_4
Xfanout786 FrameData[17] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__clkbuf_4
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1260_ _0370_ _0335_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VGND VGND VPWR VPWR
+ _0371_ sky130_fd_sc_hd__mux2_4
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 E2END[2] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
X_1191_ Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q
+ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_4
XFILLER_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0975_ _0103_ _0106_ _0073_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__a21bo_1
Xoutput301 net301 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__buf_6
Xoutput334 Inst_LUT4AB_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR SS4BEG[13] sky130_fd_sc_hd__buf_6
Xoutput312 net312 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput323 net323 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput356 net356 VGND VGND VPWR VPWR W2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput345 net345 VGND VGND VPWR VPWR SS4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput367 net367 VGND VGND VPWR VPWR W6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput378 net378 VGND VGND VPWR VPWR W6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput389 net389 VGND VGND VPWR VPWR WW4BEG[4] sky130_fd_sc_hd__buf_2
X_1527_ net743 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1458_ net65 net80 net804 net464 Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG0 sky130_fd_sc_hd__mux4_1
X_1389_ _0478_ _0481_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.EE4BEG3 sky130_fd_sc_hd__mux2_4
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0760_ net67 net807 net79 net10 Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q
+ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__mux4_1
X_2361_ W6END[3] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_2
X_2292_ Inst_LUT4AB_switch_matrix.JS2BEG1 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_1
X_1312_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q _0415_ _0416_ VGND VGND VPWR VPWR
+ _0417_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_22_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1243_ net646 net631 net636 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_39_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1174_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux _0276_ _0291_ _0292_ _0279_ VGND
+ VGND VPWR VPWR _0293_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_47_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0958_ net647 net632 net622 net618 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux4_1
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0889_ _0023_ _0021_ _0026_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR
+ VPWR _0027_ sky130_fd_sc_hd__o22ai_4
Xoutput142 net142 VGND VGND VPWR VPWR E1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput153 Inst_LUT4AB_switch_matrix.E2BEG7 VGND VGND VPWR VPWR E2BEG[7] sky130_fd_sc_hd__buf_6
Xoutput175 net175 VGND VGND VPWR VPWR EE4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput186 net186 VGND VGND VPWR VPWR EE4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput164 Inst_LUT4AB_switch_matrix.E6BEG1 VGND VGND VPWR VPWR E6BEG[11] sky130_fd_sc_hd__buf_8
Xoutput197 net197 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
XFILLER_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1930_ net44 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1861_ net774 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0812_ net93 net121 net109 net135 Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux4_1
Xinput11 E2END[5] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
Xinput22 E6END[0] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
X_1792_ net786 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput55 FrameStrobe[15] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xinput33 FrameData[14] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
Xinput44 FrameData[27] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
X_0743_ net16 net101 net129 Inst_LUT4AB_switch_matrix.E2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__mux4_2
Xinput77 N2MID[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput66 N2END[3] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
Xinput88 S1END[1] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xinput99 S2MID[0] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
X_2344_ Inst_LUT4AB_switch_matrix.JW2BEG0 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2275_ NN4END[8] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_1
X_1226_ net647 net632 net637 net408 Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q
+ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux4_1
XFILLER_25_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1157_ _0251_ _0214_ _0198_ _0252_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a31o_4
XFILLER_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1088_ _0212_ _0206_ _0203_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_4
XFILLER_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ net761 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1011_ _0138_ _0139_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q VGND VGND VPWR VPWR
+ _0140_ sky130_fd_sc_hd__mux2_1
XFILLER_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1913_ net800 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1844_ net748 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1775_ net28 net735 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0726_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_31_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2327_ SS4END[8] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_2
X_2258_ N4END[7] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
X_1209_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0050_ _0051_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o221a_1
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2189_ net747 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_1
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone36 net521 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_8
Xclone69 net624 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1560_ net740 net705 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
X_1491_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q _0529_ VGND VGND VPWR VPWR _0548_
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2112_ net786 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2043_ net797 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1827_ net778 net664 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_9_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1758_ net791 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1689_ net801 net723 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0991_ _0118_ _0119_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q VGND VGND VPWR VPWR
+ _0122_ sky130_fd_sc_hd__mux2_1
X_1612_ net760 net710 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_1543_ net770 net702 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
X_1474_ Inst_LUT4AB_switch_matrix.JN2BEG1 Inst_LUT4AB_switch_matrix.E2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_65_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2026_ net765 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_24_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout732 net733 VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout721 FrameStrobe[13] VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__clkbuf_2
Xfanout710 FrameStrobe[16] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__clkbuf_2
Xfanout754 net755 VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__clkbuf_4
Xfanout743 FrameData[8] VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__buf_4
Xfanout765 net44 VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__buf_4
Xfanout776 net777 VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__buf_4
Xfanout798 net799 VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__clkbuf_4
Xfanout787 FrameData[17] VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__buf_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1190_ _0027_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q _0307_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q
+ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a211oi_4
XFILLER_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 E2END[3] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_17_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0974_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 _0104_ _0105_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__o22a_1
Xoutput302 net302 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__buf_8
Xoutput324 net324 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput335 net335 VGND VGND VPWR VPWR SS4BEG[14] sky130_fd_sc_hd__buf_4
Xoutput313 net313 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput346 net346 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
X_1526_ net745 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
Xoutput357 net357 VGND VGND VPWR VPWR W2BEG[6] sky130_fd_sc_hd__buf_8
Xoutput368 Inst_LUT4AB_switch_matrix.W6BEG0 VGND VGND VPWR VPWR W6BEG[10] sky130_fd_sc_hd__buf_6
Xoutput379 net379 VGND VGND VPWR VPWR WW4BEG[0] sky130_fd_sc_hd__buf_2
X_1457_ net66 net81 net805 net478 Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG1 sky130_fd_sc_hd__mux4_2
X_1388_ _0479_ _0480_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q VGND VGND VPWR VPWR
+ _0481_ sky130_fd_sc_hd__mux2_4
XFILLER_67_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2009_ net801 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2360_ W6END[2] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_2
X_2291_ Inst_LUT4AB_switch_matrix.JS2BEG0 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_6
X_1311_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q _0414_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1242_ net655 net651 net626 net640 Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux4_1
XFILLER_64_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0283_ _0287_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ _0290_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__o221a_1
XFILLER_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0957_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0089_ VGND VGND VPWR VPWR _0090_
+ sky130_fd_sc_hd__and2b_1
X_0888_ _0025_ _0024_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VGND VGND VPWR VPWR
+ _0026_ sky130_fd_sc_hd__mux2_1
Xoutput143 net143 VGND VGND VPWR VPWR E1BEG[1] sky130_fd_sc_hd__buf_4
Xoutput154 net154 VGND VGND VPWR VPWR E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput176 net176 VGND VGND VPWR VPWR EE4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput165 net165 VGND VGND VPWR VPWR E6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput187 net187 VGND VGND VPWR VPWR EE4BEG[7] sky130_fd_sc_hd__buf_2
X_1509_ Inst_LG_LUT4c_frame_config_dffesr.c_reset_value _0275_ _0561_ VGND VGND VPWR
+ VPWR _0562_ sky130_fd_sc_hd__mux2_2
Xoutput198 net198 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
XFILLER_55_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ net777 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1791_ net788 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0811_ net59 net8 net65 net805 Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__mux4_1
Xinput12 E2END[6] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0742_ _0590_ _0589_ _0593_ _0564_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG3
+ sky130_fd_sc_hd__a22o_4
Xinput23 E6END[1] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 FrameData[15] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput45 FrameData[28] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput78 N2MID[7] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_2
Xinput67 N2END[4] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput56 FrameStrobe[19] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xinput89 S1END[2] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2343_ Inst_LUT4AB_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_6
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2274_ NN4END[7] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1225_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0339_ VGND VGND VPWR VPWR _0340_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1156_ _0275_ Inst_LG_LUT4c_frame_config_dffesr.LUT_flop Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR G sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_35_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1087_ _0211_ _0208_ _0189_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
XFILLER_52_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1989_ net774 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ net78 net21 net106 net134 Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q
+ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__mux4_1
XFILLER_19_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1912_ net740 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1843_ net51 net666 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1774_ net754 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0725_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__inv_1
XFILLER_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2326_ SS4END[7] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_2
X_2257_ N4END[6] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
XFILLER_72_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1208_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 _0316_ _0317_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__o22a_1
X_2188_ net749 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_1
XFILLER_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1139_ _0259_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__a21bo_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1490_ net545 _0547_ _0545_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__mux2_1
X_2111_ net789 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2042_ net799 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_47_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1826_ net782 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1757_ net793 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1688_ net741 net723 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ S4END[6] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0990_ net85 net7 net92 net120 Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q
+ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__mux4_2
X_1611_ net763 net710 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_1542_ net773 net702 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1473_ _0530_ _0531_ _0532_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q
+ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__a221o_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2025_ net767 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_47_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1809_ net758 net663 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout700 net703 VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__clkbuf_2
Xfanout733 net734 VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__clkbuf_2
Xfanout711 FrameStrobe[16] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout722 FrameStrobe[13] VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__clkbuf_2
Xfanout755 net49 VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__buf_4
Xfanout744 net745 VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__clkbuf_4
Xfanout766 net767 VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__buf_4
Xfanout799 net30 VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__buf_4
Xfanout777 net40 VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__clkbuf_4
Xfanout788 net789 VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__buf_4
XFILLER_65_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0973_ _0086_ _0098_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__or2_2
Xoutput314 net314 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput303 net303 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__buf_6
Xoutput325 net325 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput358 net358 VGND VGND VPWR VPWR W2BEG[7] sky130_fd_sc_hd__buf_6
X_1525_ net747 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ sky130_fd_sc_hd__dlxtp_1
Xoutput336 net336 VGND VGND VPWR VPWR SS4BEG[15] sky130_fd_sc_hd__buf_4
Xoutput347 net347 VGND VGND VPWR VPWR W1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput369 Inst_LUT4AB_switch_matrix.W6BEG1 VGND VGND VPWR VPWR W6BEG[11] sky130_fd_sc_hd__buf_6
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1456_ net63 net82 net136 net631 Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG2 sky130_fd_sc_hd__mux4_2
X_1387_ _0235_ _0625_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q VGND VGND VPWR VPWR
+ _0480_ sky130_fd_sc_hd__mux2_4
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2008_ net741 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer90 net635 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1310_ net464 net415 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q VGND VGND VPWR VPWR
+ _0415_ sky130_fd_sc_hd__mux2_1
X_1241_ _0351_ _0350_ _0354_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JN2BEG7 sky130_fd_sc_hd__o22a_1
XFILLER_49_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1172_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0286_ VGND VGND
+ VPWR VPWR _0291_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_47_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0956_ net657 net652 net627 net642 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__mux4_1
X_0887_ net60 net68 net3 net11 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__mux4_1
Xoutput144 Inst_LUT4AB_switch_matrix.E1BEG2 VGND VGND VPWR VPWR E1BEG[2] sky130_fd_sc_hd__buf_8
Xoutput155 net155 VGND VGND VPWR VPWR E2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput166 net166 VGND VGND VPWR VPWR E6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput177 net177 VGND VGND VPWR VPWR EE4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput188 net188 VGND VGND VPWR VPWR EE4BEG[8] sky130_fd_sc_hd__buf_2
X_1508_ _0538_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q VGND VGND VPWR VPWR _0561_
+ sky130_fd_sc_hd__nand2_4
Xoutput199 net199 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
X_1439_ net434 _0640_ Inst_LUT4AB_switch_matrix.JS2BEG2 _0624_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1790_ net790 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0810_ _0655_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__a21bo_1
Xinput13 E2END[7] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
X_0741_ _0591_ _0592_ _0563_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__mux2_1
Xinput24 EE4END[0] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput35 FrameData[16] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
Xinput46 FrameData[29] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput68 N2END[5] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
Xinput57 FrameStrobe[5] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
Xinput79 N4END[0] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2273_ NN4END[6] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_1
X_1224_ net656 net652 net627 net642 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__mux4_1
X_1155_ _0274_ _0268_ _0266_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_35_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1086_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0196_ _0209_ _0210_
+ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__o211a_1
XFILLER_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1988_ net777 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0939_ _0072_ Inst_LE_LUT4c_frame_config_dffesr.c_I0mux _0071_ VGND VGND VPWR VPWR
+ _0073_ sky130_fd_sc_hd__o21ai_4
XFILLER_68_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1911_ net743 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1842_ net50 net666 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1773_ net756 net728 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0724_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__inv_1
XFILLER_69_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2325_ SS4END[6] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2256_ N4END[5] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
X_1207_ _0319_ _0323_ _0315_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_4
X_2187_ net751 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__buf_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1138_ net646 net621 net635 net417 Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q
+ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__mux4_2
XFILLER_43_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1069_ _0190_ _0192_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__or2_1
XFILLER_68_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2110_ net791 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2041_ net801 net694 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_17_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1825_ net784 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1756_ net795 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1687_ net742 net723 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2308_ S4END[5] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_68_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ Inst_LUT4AB_switch_matrix.JN2BEG0 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__buf_4
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1610_ net764 net711 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_1541_ net775 net702 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
X_1472_ _0139_ _0068_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR
+ _0532_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2024_ net768 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1808_ net781 net663 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1739_ net762 net725 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout701 net703 VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout723 FrameStrobe[13] VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__buf_1
Xfanout712 net55 VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__clkbuf_2
Xfanout756 net757 VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__clkbuf_4
Xfanout734 net735 VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__clkbuf_2
Xfanout745 net53 VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__buf_4
Xfanout767 net43 VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_37_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout778 net779 VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__buf_4
Xfanout789 net35 VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__buf_4
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0972_ _0086_ _0099_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__nand2_1
Xoutput304 net443 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__buf_6
Xoutput326 net326 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput315 net315 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__buf_2
X_1524_ net749 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ sky130_fd_sc_hd__dlxtp_1
Xoutput359 net359 VGND VGND VPWR VPWR W2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput348 Inst_LUT4AB_switch_matrix.W1BEG1 VGND VGND VPWR VPWR W1BEG[1] sky130_fd_sc_hd__buf_4
Xoutput337 net337 VGND VGND VPWR VPWR SS4BEG[1] sky130_fd_sc_hd__buf_2
X_1455_ net64 net135 net79 net412 Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG3 sky130_fd_sc_hd__mux4_1
X_1386_ net647 _0082_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q VGND VGND VPWR VPWR
+ _0479_ sky130_fd_sc_hd__mux2_4
X_2007_ net742 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer80 _0027_ VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__buf_6
Xrebuffer91 H VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1240_ _0352_ _0353_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q VGND VGND VPWR VPWR
+ _0354_ sky130_fd_sc_hd__mux2_1
X_1171_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 _0284_ VGND VGND
+ VPWR VPWR _0290_ sky130_fd_sc_hd__or2_1
XFILLER_66_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0955_ net66 net94 net9 net138 Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q
+ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_30_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0886_ net88 net96 net90 net116 Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q
+ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__mux4_1
Xoutput145 Inst_LUT4AB_switch_matrix.E1BEG3 VGND VGND VPWR VPWR E1BEG[3] sky130_fd_sc_hd__buf_4
Xoutput156 net156 VGND VGND VPWR VPWR E2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput167 net167 VGND VGND VPWR VPWR E6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput189 net189 VGND VGND VPWR VPWR EE4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput178 Inst_LUT4AB_switch_matrix.EE4BEG1 VGND VGND VPWR VPWR EE4BEG[13] sky130_fd_sc_hd__buf_6
X_1507_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q _0529_ VGND VGND VPWR VPWR _0560_
+ sky130_fd_sc_hd__nand2_1
X_1438_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q _0523_ _0522_ VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.NN4BEG0 sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_38_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1369_ net4 net660 net656 net651 Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__mux4_1
XFILLER_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0740_ net61 net67 net79 net10 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__mux4_1
Xinput14 E2MID[0] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
Xinput25 EE4END[1] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput36 FrameData[18] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput69 N2END[6] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
Xinput58 FrameStrobe[9] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
Xinput47 FrameData[2] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2272_ NN4END[5] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_1
X_1223_ _0337_ _0338_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.M_AD sky130_fd_sc_hd__mux2_4
XFILLER_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1154_ _0269_ _0273_ _0227_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1085_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0193_ _0198_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__o22a_1
XFILLER_52_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1987_ net779 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0938_ _0067_ _0068_ _0070_ _0069_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux4_2
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0869_ _0710_ _0008_ _0697_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__mux2_1
XFILLER_28_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ net745 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_42_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1841_ net758 net665 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1772_ net761 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0723_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__inv_1
X_2324_ SS4END[5] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2255_ N4END[4] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_1
X_2186_ net753 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_1
X_1206_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0050_ _0321_ _0322_
+ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__o211a_1
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1137_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q _0257_ VGND VGND VPWR VPWR _0258_
+ sky130_fd_sc_hd__and2b_1
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1068_ _0190_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone17 G VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__buf_6
Xclone39 net657 VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__buf_8
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2040_ net741 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1824_ net787 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1755_ net797 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1686_ net744 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_13_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2307_ S4END[4] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_2
X_2238_ Inst_LUT4AB_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_68_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ EE4END[6] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ net776 net702 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
X_1471_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _0615_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
+ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2023_ net771 net690 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1807_ net803 net661 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1738_ net764 net724 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1669_ net774 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout724 net726 VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__buf_2
Xfanout702 net703 VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__clkbuf_2
Xfanout713 net714 VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__clkbuf_2
Xfanout746 FrameData[6] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__buf_4
Xfanout735 FrameStrobe[10] VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__clkbuf_2
Xfanout757 net48 VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__buf_4
Xfanout768 net769 VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__clkbuf_4
Xfanout779 net39 VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__clkbuf_4
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0971_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0100_ _0101_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_70_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput305 net305 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__buf_6
Xoutput316 net316 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__buf_2
X_1523_ net751 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
Xoutput349 Inst_LUT4AB_switch_matrix.W1BEG2 VGND VGND VPWR VPWR W1BEG[2] sky130_fd_sc_hd__buf_8
Xoutput327 net327 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput338 net338 VGND VGND VPWR VPWR SS4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1454_ net445 Inst_LUT4AB_switch_matrix.JN2BEG3 _0165_ _0018_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG0
+ sky130_fd_sc_hd__mux4_1
X_1385_ net60 net3 net88 net642 Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux4_1
XFILLER_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2006_ net744 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer81 net476 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__buf_6
XFILLER_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer92 H VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__buf_6
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1170_ _0264_ _0265_ _0256_ _0255_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__mux4_2
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0954_ net85 net109 net8 Inst_LUT4AB_switch_matrix.E2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_30_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0885_ _0022_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_65_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput146 net146 VGND VGND VPWR VPWR E2BEG[0] sky130_fd_sc_hd__buf_8
Xoutput157 net157 VGND VGND VPWR VPWR E2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput168 net168 VGND VGND VPWR VPWR E6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput179 net179 VGND VGND VPWR VPWR EE4BEG[14] sky130_fd_sc_hd__buf_6
X_1506_ net547 _0559_ _0557_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__mux2_2
X_1437_ net61 net660 net807 net477 Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
+ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__mux4_1
X_1368_ net625 net641 net647 net477 Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__mux4_1
XFILLER_46_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1299_ _0401_ _0399_ _0404_ _0583_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG0
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput15 E2MID[1] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
Xinput26 EE4END[2] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput37 FrameData[19] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput59 N1END[0] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
Xinput48 FrameData[30] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
XFILLER_42_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2340_ Inst_LUT4AB_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__buf_1
XFILLER_69_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2271_ NN4END[4] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_1
X_1222_ _0337_ net483 net522 VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__mux2_4
X_1153_ _0270_ _0271_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1084_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0194_ VGND VGND
+ VPWR VPWR _0209_ sky130_fd_sc_hd__or2_1
X_1986_ net783 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0937_ _0060_ _0050_ Inst_LE_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0071_ sky130_fd_sc_hd__a21bo_1
X_0868_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ _0695_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__mux2_1
X_0799_ net85 net26 net2 net805 Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__mux4_1
XFILLER_57_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1840_ net781 net665 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1771_ net763 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0722_ Inst_LH_LUT4c_frame_config_dffesr.c_out_mux VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__inv_2
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2323_ SS4END[4] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_2
X_2254_ net78 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_2
X_2185_ net758 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__buf_1
X_1205_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0316_ _0317_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__o22a_1
X_1136_ net655 net651 net625 net640 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux4_1
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1067_ _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone18 net428 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__buf_8
X_1969_ net758 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1823_ net788 net663 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1754_ net799 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1685_ net746 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2306_ net106 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__buf_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2237_ Inst_LUT4AB_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ EE4END[5] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2099_ net750 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1119_ net647 net485 net637 net402 Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q
+ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_51_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1470_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _0221_ VGND VGND VPWR VPWR _0530_
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2022_ net772 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_65_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1806_ net755 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1737_ net766 net725 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1668_ net777 net717 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout703 FrameStrobe[18] VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout714 net715 VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout725 net726 VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__clkbuf_2
Xfanout747 FrameData[6] VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__clkbuf_4
Xfanout736 net738 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__buf_2
Xfanout758 net759 VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__clkbuf_4
X_1599_ net788 net710 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ sky130_fd_sc_hd__dlxtp_1
Xfanout769 net42 VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__buf_4
XFILLER_73_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0970_ _0101_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput306 net306 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput317 net317 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__buf_6
X_1522_ net753 net700 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
Xoutput328 net328 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput339 net339 VGND VGND VPWR VPWR SS4BEG[3] sky130_fd_sc_hd__buf_2
X_1453_ net645 _0068_ Inst_LUT4AB_switch_matrix.JN2BEG0 _0084_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG1
+ sky130_fd_sc_hd__mux4_1
X_1384_ _0586_ _0471_ _0477_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E6BEG0
+ sky130_fd_sc_hd__a21o_1
XFILLER_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2005_ net746 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer82 net487 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkbuf_2
Xrebuffer60 net455 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer93 net512 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_41_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0953_ _0082_ _0083_ _0085_ _0084_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q
+ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_30_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0884_ net635 net630 net621 net617 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__mux4_2
Xoutput147 net147 VGND VGND VPWR VPWR E2BEG[1] sky130_fd_sc_hd__buf_4
Xoutput158 net158 VGND VGND VPWR VPWR E2BEGb[4] sky130_fd_sc_hd__buf_2
X_1505_ Inst_LF_LUT4c_frame_config_dffesr.c_reset_value _0213_ _0558_ VGND VGND VPWR
+ VPWR _0559_ sky130_fd_sc_hd__mux2_2
Xoutput169 net169 VGND VGND VPWR VPWR E6BEG[5] sky130_fd_sc_hd__buf_2
X_1436_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q _0521_ _0519_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q
+ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__o211a_1
X_1367_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q _0462_ _0461_ VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.SS4BEG0 sky130_fd_sc_hd__o21ba_1
X_1298_ _0402_ _0403_ _0582_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput16 E2MID[2] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 EE4END[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput38 FrameData[1] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
Xinput49 FrameData[31] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2270_ Inst_LUT4AB_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__buf_6
X_1221_ net640 net625 _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__mux2_4
XFILLER_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1152_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0251_ _0253_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_35_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1083_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0196_ _0198_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__o221a_1
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1985_ net785 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0936_ net70 net98 net26 net126 Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q
+ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux4_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0867_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ _0695_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__mux2_1
X_0798_ net109 net113 net121 net135 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__mux4_1
X_1419_ _0506_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__inv_1
XFILLER_68_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1770_ net765 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0721_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__inv_1
X_2322_ Inst_LUT4AB_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2253_ net77 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_1
X_1204_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0051_ VGND VGND
+ VPWR VPWR _0321_ sky130_fd_sc_hd__or2_1
X_2184_ net781 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_1
X_1135_ net64 net92 net27 net120 Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q
+ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux4_2
XFILLER_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1066_ _0096_ _0097_ _0088_ _0087_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q
+ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux4_2
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1968_ net780 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1899_ net762 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0919_ _0053_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__inv_2
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1822_ net34 net663 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_60_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1753_ net801 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1684_ net749 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2305_ net105 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_68_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ EE4END[4] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ net753 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1118_ net656 net652 net627 net640 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux4_1
X_1049_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0057_ _0153_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_51_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2021_ net774 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1805_ net757 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1736_ net42 net725 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1667_ net779 net717 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout704 FrameStrobe[17] VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__clkbuf_2
X_1598_ net790 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
Xfanout715 net55 VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout748 net749 VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__clkbuf_4
Xfanout737 net738 VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__buf_2
Xfanout726 FrameStrobe[12] VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__clkbuf_2
Xfanout759 net47 VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__clkbuf_4
X_2219_ net686 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput307 net307 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__buf_2
X_1521_ net759 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
Xoutput329 net329 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput318 net318 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__buf_2
XFILLER_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1452_ net415 Inst_LUT4AB_switch_matrix.JN2BEG1 net658 _0255_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG2
+ sky130_fd_sc_hd__mux4_2
X_1383_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q _0472_ _0474_ _0476_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q
+ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__o221a_1
X_2004_ net52 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1719_ net742 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer61 net456 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer94 Inst_LUT4AB_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0952_ net68 net11 net112 net124 Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q
+ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__mux4_2
XFILLER_13_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0883_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q _0020_ VGND VGND VPWR VPWR _0021_
+ sky130_fd_sc_hd__and2b_1
Xoutput148 net148 VGND VGND VPWR VPWR E2BEG[2] sky130_fd_sc_hd__buf_6
Xoutput159 net159 VGND VGND VPWR VPWR E2BEGb[5] sky130_fd_sc_hd__buf_2
X_1504_ _0538_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q VGND VGND VPWR VPWR _0558_
+ sky130_fd_sc_hd__nand2_4
X_1435_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__inv_1
X_1366_ net61 net660 net807 net415 Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q
+ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__mux4_1
X_1297_ net64 net806 net80 net7 Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_38_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput17 E2MID[3] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
Xinput28 FrameData[0] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput39 FrameData[20] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_1
X_1220_ _0335_ net475 Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ _0336_ sky130_fd_sc_hd__mux2_4
XFILLER_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1151_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0250_ _0239_ VGND
+ VGND VPWR VPWR _0271_ sky130_fd_sc_hd__or3b_1
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1082_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0193_ _0194_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_35_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1984_ net786 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0935_ net82 net122 net9 Inst_LUT4AB_switch_matrix.JN2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux4_2
X_0866_ _0708_ _0707_ _0697_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__mux2_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0797_ _0572_ _0643_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0644_ sky130_fd_sc_hd__o21a_1
X_1418_ net627 _0097_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q VGND VGND VPWR VPWR
+ _0506_ sky130_fd_sc_hd__mux2_1
XFILLER_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1349_ net414 _0097_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q VGND VGND VPWR VPWR
+ _0447_ sky130_fd_sc_hd__mux2_1
XFILLER_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0720_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__inv_2
X_2321_ Inst_LUT4AB_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_2
X_2252_ net76 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_2
X_1203_ _0164_ _0165_ _0173_ _0172_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q
+ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__mux4_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2183_ net803 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
X_1134_ net83 net119 net805 net479 Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux4_2
XFILLER_65_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1065_ _0082_ _0083_ _0085_ _0084_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux4_2
XFILLER_18_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1967_ net802 net683 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0918_ net525 _0047_ _0039_ _0038_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q
+ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux4_2
X_1898_ net764 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0849_ net1 _0605_ _0650_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__o21ai_4
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1821_ net792 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1752_ net741 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1683_ net751 net723 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2304_ net104 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_1
X_2235_ Inst_LUT4AB_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_68_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ _0235_ _0236_ _0238_ _0237_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q
+ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__mux4_2
XFILLER_53_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2097_ net759 net738 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1048_ _0164_ _0165_ _0173_ _0172_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q
+ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_51_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2020_ net777 net689 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1804_ net760 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1735_ net770 net725 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1666_ net783 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout705 FrameStrobe[17] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__dlymetal6s2s_1
X_1597_ net792 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
Xfanout738 net739 VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkbuf_2
Xfanout749 net52 VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__buf_4
Xfanout727 FrameStrobe[12] VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__buf_2
Xfanout716 FrameStrobe[14] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__buf_2
XFILLER_65_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2218_ net690 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__buf_1
X_2149_ net16 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_1
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput308 net308 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__buf_2
X_1520_ net781 net701 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
Xoutput319 net319 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__buf_4
X_1451_ net411 _0640_ Inst_LUT4AB_switch_matrix.JN2BEG2 _0624_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1382_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q _0475_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q
+ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__a21bo_1
XFILLER_67_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2003_ net750 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1718_ net744 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1649_ net758 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer62 net457 VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer95 net488 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer130 net402 VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0951_ net80 net112 net123 Inst_LUT4AB_switch_matrix.JS2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux4_2
XFILLER_9_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0882_ net654 net650 net625 net641 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__mux4_1
Xoutput149 net149 VGND VGND VPWR VPWR E2BEG[3] sky130_fd_sc_hd__buf_2
X_1503_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q _0529_ VGND VGND VPWR VPWR _0557_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_34_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1434_ net632 _0595_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q VGND VGND VPWR VPWR
+ _0520_ sky130_fd_sc_hd__mux2_1
X_1365_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q _0460_ _0458_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q
+ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__o211a_1
X_1296_ net804 net112 net120 net136 Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_38_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 E2MID[4] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 FrameData[10] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_70_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1150_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0239_ _0250_ VGND
+ VGND VPWR VPWR _0270_ sky130_fd_sc_hd__or3b_1
X_1081_ _0200_ _0205_ _0189_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_35_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ net789 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0934_ net78 net21 net106 net134 Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q
+ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux4_2
X_0865_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0695_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__mux2_1
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0796_ net462 net411 net619 net416 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__mux4_2
X_1417_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q _0504_ VGND VGND VPWR VPWR _0505_
+ sky130_fd_sc_hd__nand2_1
XFILLER_68_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1348_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q _0445_ VGND VGND VPWR VPWR _0446_
+ sky130_fd_sc_hd__nand2_1
X_1279_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0384_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o21a_1
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2320_ Inst_LUT4AB_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__buf_1
X_2251_ net75 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
X_1202_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 _0050_ _0051_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__o221a_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1133_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0250_ _0239_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux4_1
XFILLER_65_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1064_ _0187_ _0188_ Inst_LF_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0189_ sky130_fd_sc_hd__mux2_4
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1966_ net754 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0917_ _0028_ _0029_ _0019_ _0018_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q
+ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__mux4_2
X_1897_ net766 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0848_ _0689_ _0690_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q VGND VGND VPWR VPWR
+ _0691_ sky130_fd_sc_hd__mux2_1
X_0779_ _0616_ _0626_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q VGND VGND VPWR VPWR
+ _0627_ sky130_fd_sc_hd__mux2_1
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1820_ net794 net662 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1751_ net742 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1682_ net753 net722 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2303_ net103 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_2
XFILLER_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2234_ net56 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_68_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1116_ net84 net96 net11 net124 Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q
+ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux4_2
X_2096_ net780 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1047_ net63 net91 net25 net119 Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q
+ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_51_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1949_ net793 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_8_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1803_ net762 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1734_ net773 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1665_ net785 net716 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xfanout706 FrameStrobe[17] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__clkbuf_2
X_1596_ net794 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
Xfanout728 net729 VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__clkbuf_2
Xfanout739 FrameStrobe[0] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__clkbuf_2
Xfanout717 FrameStrobe[14] VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2217_ FrameStrobe[2] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2148_ net15 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_1
XFILLER_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2079_ net789 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput309 net309 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__buf_2
X_1450_ net643 Inst_LUT4AB_switch_matrix.E2BEG3 _0165_ _0018_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_4_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1381_ _0097_ net658 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q VGND VGND VPWR VPWR
+ _0475_ sky130_fd_sc_hd__mux2_1
X_2002_ net752 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1717_ net746 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1648_ net781 net719 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_1579_ net763 net707 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer41 net436 VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_2
Xrebuffer63 net458 VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer85 Inst_LUT4AB_switch_matrix.JW2BEG4 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_24_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer131 _0046_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__buf_6
Xrebuffer120 net515 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0950_ net76 net19 net104 net132 Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q
+ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__mux4_1
XFILLER_9_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0881_ net65 net8 net93 net139 Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q
+ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__mux4_2
XFILLER_40_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1502_ net541 _0556_ _0554_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__mux2_1
X_1433_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q _0518_ VGND VGND VPWR VPWR _0519_
+ sky130_fd_sc_hd__nand2_1
X_1364_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__inv_1
X_1295_ _0582_ _0400_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q VGND VGND VPWR VPWR
+ _0401_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_38_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput19 E2MID[5] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1080_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0196_ _0198_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ _0204_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__o221a_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ net791 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0933_ net77 net133 net20 Inst_LUT4AB_switch_matrix.JN2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux4_1
X_0864_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0695_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__mux2_1
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0795_ _0641_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q VGND VGND VPWR VPWR _0642_
+ sky130_fd_sc_hd__or2_4
X_1416_ net658 _0019_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q VGND VGND VPWR VPWR
+ _0504_ sky130_fd_sc_hd__mux2_1
X_1347_ net658 _0173_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q VGND VGND VPWR VPWR
+ _0445_ sky130_fd_sc_hd__mux2_1
XFILLER_68_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1278_ _0578_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__or2_4
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2250_ net74 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_2
X_1201_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0316_ _0317_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o22a_1
X_2181_ Inst_LUT4AB_switch_matrix.EE4BEG2 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
X_1132_ _0252_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__inv_1
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1063_ _0105_ _0060_ _0050_ _0102_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a31o_1
XFILLER_21_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1965_ net756 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0916_ _0030_ _0048_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__nand2_1
X_1896_ net768 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0847_ _0625_ _0624_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q VGND VGND VPWR VPWR
+ _0690_ sky130_fd_sc_hd__mux2_1
X_0778_ _0625_ _0624_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q VGND VGND VPWR VPWR
+ _0626_ sky130_fd_sc_hd__mux2_1
X_2379_ WW4END[11] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1750_ net744 net729 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1681_ net758 net723 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2302_ net102 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_1
X_2233_ net702 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_1
X_2164_ E6END[11] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
X_1115_ net23 net108 net140 net489 Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q
+ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__mux4_2
X_2095_ net802 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1046_ net79 net135 net111 Inst_LUT4AB_switch_matrix.JW2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_51_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1948_ net795 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1879_ net742 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_8_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1802_ net764 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1733_ net775 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1664_ net786 net717 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1595_ net796 net710 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
Xfanout729 net730 VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__clkbuf_4
Xfanout707 FrameStrobe[17] VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout718 FrameStrobe[14] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__clkbuf_2
X_2216_ net699 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__buf_1
X_2147_ net14 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
X_2078_ net791 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1029_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 _0055_ _0154_ _0156_
+ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__o211a_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1380_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q _0473_ VGND VGND VPWR VPWR _0474_
+ sky130_fd_sc_hd__and2b_1
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2001_ net759 net688 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_67_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1716_ net749 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1647_ net803 net719 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
X_1578_ net765 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer42 net437 VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkbuf_2
Xrebuffer64 net459 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer53 net448 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer86 Inst_LUT4AB_switch_matrix.M_AB VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer121 net516 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer132 Inst_LUT4AB_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0880_ net81 net8 net126 Inst_LUT4AB_switch_matrix.E2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__mux4_2
X_1501_ Inst_LE_LUT4c_frame_config_dffesr.c_reset_value _0131_ _0555_ VGND VGND VPWR
+ VPWR _0556_ sky130_fd_sc_hd__mux2_2
X_1432_ _0029_ _0249_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q VGND VGND VPWR VPWR
+ _0518_ sky130_fd_sc_hd__mux2_1
X_1363_ net411 _0595_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR
+ _0459_ sky130_fd_sc_hd__mux2_1
X_1294_ net633 net628 net619 net618 Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_38_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1981_ net793 net685 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0932_ _0066_ _0063_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.JN2BEG5 sky130_fd_sc_hd__mux2_4
X_0863_ _0705_ _0702_ _0696_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__mux2_4
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0794_ net653 net444 net623 net643 Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux4_2
X_1415_ _0502_ _0503_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.NN4BEG3 sky130_fd_sc_hd__mux2_4
X_1346_ _0443_ _0444_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.SS4BEG3 sky130_fd_sc_hd__mux2_1
XFILLER_68_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1277_ net633 net628 net619 net404 Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
+ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__mux4_2
XFILLER_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1200_ _0030_ _0049_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__or2_1
X_1131_ _0239_ _0250_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__and2_1
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1062_ _0067_ _0068_ _0070_ _0069_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux4_2
XFILLER_65_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1964_ net761 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0915_ _0030_ _0048_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__or2_4
X_1895_ net771 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0846_ _0613_ _0614_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q VGND VGND VPWR VPWR
+ _0689_ sky130_fd_sc_hd__mux2_1
X_0777_ net69 net114 net12 net125 Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q
+ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__mux4_2
X_2378_ WW4END[10] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1329_ net414 _0097_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _0431_ sky130_fd_sc_hd__mux2_1
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput290 net290 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_47_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1680_ net780 net720 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2301_ net101 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__buf_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2232_ net707 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_1
X_2163_ E6END[10] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
X_1114_ net76 net19 net104 net132 Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q
+ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__mux4_1
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2094_ net754 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1045_ _0171_ _0168_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.JW2BEG2 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_51_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1947_ net797 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1878_ net745 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0829_ _0671_ _0672_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q VGND VGND VPWR VPWR
+ _0673_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1801_ net766 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_13_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1732_ net776 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1663_ net789 net717 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1594_ net798 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
Xfanout708 net709 VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__clkbuf_2
Xfanout719 FrameStrobe[14] VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2215_ net739 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2077_ net793 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1028_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0155_ VGND VGND
+ VPWR VPWR _0156_ sky130_fd_sc_hd__or2_1
XFILLER_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2000_ net780 net687 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1715_ net751 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1646_ net755 net715 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
X_1577_ net43 net707 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer10 net403 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2129_ clknet_1_0__leaf_UserCLK_regs _0002_ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer43 net438 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkbuf_2
Xrebuffer54 net449 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_2
Xrebuffer65 net460 VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer87 Inst_LUT4AB_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer122 net517 VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1500_ _0538_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR _0555_
+ sky130_fd_sc_hd__nand2_4
X_1431_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q _0513_ _0515_ _0517_ VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.NN4BEG1 sky130_fd_sc_hd__o22a_1
X_1362_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q _0457_ VGND VGND VPWR VPWR _0458_
+ sky130_fd_sc_hd__nand2_1
X_1293_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q _0398_ VGND VGND VPWR VPWR _0399_
+ sky130_fd_sc_hd__or2_1
XFILLER_23_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1629_ net792 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1980_ net795 net684 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0931_ _0064_ _0065_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VGND VGND VPWR VPWR
+ _0066_ sky130_fd_sc_hd__mux2_1
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0862_ _0704_ _0703_ _0697_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__mux2_1
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0793_ net76 net19 net104 net132 Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q
+ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux4_2
X_1414_ net647 _0082_ _0235_ _0604_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q
+ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux4_2
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1345_ net645 _0082_ _0235_ _0661_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__mux4_1
XFILLER_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1276_ net446 net444 net463 net643 Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__mux4_1
XFILLER_24_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1130_ _0239_ _0250_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__or2_1
X_1061_ _0186_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR C sky130_fd_sc_hd__mux2_4
XFILLER_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1963_ net763 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0914_ _0048_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_2
X_1894_ net772 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0845_ _0686_ _0687_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q VGND VGND VPWR VPWR
+ _0688_ sky130_fd_sc_hd__mux2_1
X_0776_ net86 net137 net110 Inst_LUT4AB_switch_matrix.JN2BEG1 Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__mux4_2
X_2377_ WW4END[9] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1328_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q _0429_ VGND VGND VPWR VPWR _0430_
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1259_ _0575_ _0369_ _0368_ _0367_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a2bb2o_4
XTAP_TAPCELL_ROW_19_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput280 net280 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput291 net291 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2300_ net100 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_1
X_2231_ net711 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_1
X_2162_ E6END[9] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_1
XFILLER_38_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2093_ net756 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1113_ net18 net131 net103 net429 Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q
+ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__mux4_2
X_1044_ _0170_ _0169_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VGND VGND VPWR VPWR
+ _0171_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1946_ net30 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1877_ net746 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0828_ _0661_ _0660_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q VGND VGND VPWR VPWR
+ _0672_ sky130_fd_sc_hd__mux2_1
X_0759_ _0606_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q
+ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__a21bo_1
XFILLER_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1800_ net769 net734 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1731_ net778 net726 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1662_ net790 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_1593_ net800 net709 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
Xfanout709 FrameStrobe[16] VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__clkbuf_2
X_2214_ net755 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_1
X_2145_ net413 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_4
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2076_ net795 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1027_ _0052_ _0054_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__or2_1
X_1929_ net766 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1714_ net753 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1645_ net757 net715 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
X_1576_ net769 net707 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer11 Inst_LUT4AB_switch_matrix.M_AH VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__buf_6
X_2128_ clknet_1_0__leaf_UserCLK_regs _0001_ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer22 net617 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_8
Xrebuffer44 net439 VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkbuf_2
Xrebuffer55 net450 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_2
Xrebuffer33 net486 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__buf_6
X_2059_ net763 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer66 net461 VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer88 net430 VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_24_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer123 net518 VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q _0516_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q
+ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a21bo_1
X_1361_ _0029_ _0256_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR
+ _0457_ sky130_fd_sc_hd__mux2_1
X_1292_ net446 net638 net623 net643 Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux4_1
XFILLER_48_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1628_ net794 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
X_1559_ net743 net705 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0930_ net89 net115 net97 net660 Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q
+ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux4_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0861_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0695_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__mux2_1
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0792_ net75 net18 net131 Inst_LUT4AB_switch_matrix.JS2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__mux4_2
XFILLER_5_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1413_ net60 net3 net116 net642 Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q
+ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__mux4_1
XFILLER_68_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1344_ net60 net3 net116 net445 Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__mux4_1
X_1275_ _0378_ _0380_ _0383_ _0577_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1060_ _0178_ _0185_ _0174_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_25_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ net765 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0913_ net525 _0047_ _0039_ _0038_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q
+ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__mux4_2
X_1893_ net774 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0844_ _0661_ _0660_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q VGND VGND VPWR VPWR
+ _0687_ sky130_fd_sc_hd__mux2_1
X_0775_ _0619_ _0620_ _0623_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JN2BEG1 sky130_fd_sc_hd__o2bb2a_4
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2376_ WW4END[8] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_2
X_1327_ net658 _0039_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _0429_ sky130_fd_sc_hd__mux2_1
XFILLER_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1258_ Inst_LUT4AB_switch_matrix.JS2BEG7 Inst_LUT4AB_switch_matrix.JW2BEG7 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux2_4
XFILLER_71_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1189_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q Inst_LUT4AB_switch_matrix.JN2BEG4
+ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_19_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput270 net270 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput281 net281 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput292 net292 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2230_ net714 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
X_2161_ E6END[8] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_1
X_2092_ net760 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1112_ _0231_ _0229_ _0234_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JS2BEG6 sky130_fd_sc_hd__o22a_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1043_ net60 net66 net27 net804 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_16_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1945_ net800 net682 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1876_ net749 net671 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0827_ _0669_ _0670_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q VGND VGND VPWR VPWR
+ _0671_ sky130_fd_sc_hd__mux2_1
X_0758_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q _0607_ VGND VGND VPWR VPWR _0608_
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2359_ net134 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_67_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1730_ net782 net725 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1661_ net792 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1592_ net740 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_2213_ net757 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__buf_1
X_2144_ Inst_LUT4AB_switch_matrix.E2BEG5 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_4
X_2075_ net797 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1026_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0057_ _0153_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__o22a_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1928_ net769 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_12_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1859_ net779 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1713_ net758 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1644_ net46 net715 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
X_1575_ net770 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer12 net405 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer23 net617 VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_6
Xrebuffer45 net440 VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__clkbuf_2
X_2127_ clknet_1_1__leaf_UserCLK_regs _0000_ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.LUT_flop
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer34 net427 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__buf_6
XFILLER_66_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2058_ net765 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer67 Inst_LUT4AB_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_2
Xrebuffer56 net451 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ net20 net133 net105 Inst_LUT4AB_switch_matrix.JN2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__mux4_1
Xrebuffer89 net430 VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_24_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer124 net519 VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1360_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q _0456_ _0455_ VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.SS4BEG1 sky130_fd_sc_hd__o21ba_4
X_1291_ _0392_ _0394_ _0397_ _0581_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1627_ net796 net714 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
X_1558_ net745 net705 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
X_1489_ Inst_LB_LUT4c_frame_config_dffesr.c_reset_value _0011_ _0546_ VGND VGND VPWR
+ VPWR _0547_ sky130_fd_sc_hd__mux2_2
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0860_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ _0695_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__mux2_1
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0791_ _0567_ _0568_ _0571_ _0637_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q
+ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__mux4_2
X_1412_ _0499_ _0501_ _0497_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.EE4BEG0
+ sky130_fd_sc_hd__a21oi_1
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1343_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q _0442_ _0441_ VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.WW4BEG0 sky130_fd_sc_hd__o21ba_1
XFILLER_68_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1274_ _0381_ _0382_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VGND VGND VPWR VPWR
+ _0383_ sky130_fd_sc_hd__mux2_1
XFILLER_68_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0989_ net27 net138 net107 Inst_LUT4AB_switch_matrix.JW2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__mux4_2
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 FrameStrobe[3] VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1961_ net767 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0912_ net76 net19 net104 net132 Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q
+ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__mux4_1
X_1892_ net40 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0843_ _0669_ _0670_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q VGND VGND VPWR VPWR
+ _0686_ sky130_fd_sc_hd__mux2_1
X_0774_ _0621_ _0622_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q VGND VGND VPWR VPWR
+ _0623_ sky130_fd_sc_hd__mux2_1
X_2375_ WW4END[7] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_2
X_1326_ _0427_ _0428_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.WW4BEG3 sky130_fd_sc_hd__mux2_4
Xclone8 _0337_ _0338_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VGND VGND VPWR VPWR
+ net402 sky130_fd_sc_hd__mux2_4
X_1257_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q Inst_LUT4AB_switch_matrix.E2BEG7
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__a21oi_1
X_1188_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__inv_2
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput260 net260 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput271 net271 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput282 Inst_LUT4AB_switch_matrix.NN4BEG1 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__buf_6
Xoutput293 net293 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_59_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2160_ E6END[7] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_1
X_2091_ net762 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1111_ _0232_ _0233_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q VGND VGND VPWR VPWR
+ _0234_ sky130_fd_sc_hd__mux2_1
X_1042_ net110 net122 net114 net136 Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q
+ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux4_1
X_1944_ net741 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1875_ net750 net670 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0826_ net72 net15 net100 net128 Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q
+ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__mux4_1
X_0757_ net653 net649 net624 net644 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__mux4_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2358_ net133 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1309_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__inv_1
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1660_ net794 net718 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
X_1591_ net743 net710 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_2212_ net760 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
X_2143_ Inst_LUT4AB_switch_matrix.E2BEG4 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_8
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2074_ net799 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1025_ _0052_ _0054_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__nand2_1
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1927_ net770 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1858_ net783 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0809_ net633 net628 net620 net404 Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
+ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux4_2
X_1789_ net792 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1712_ net781 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1643_ net45 net715 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1574_ net773 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_2126_ net755 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer35 net435 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkbuf_2
Xrebuffer13 Inst_LUT4AB_switch_matrix.M_AH VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer46 net441 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkbuf_2
X_2057_ net767 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer57 net452 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ _0137_ _0134_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.JN2BEG4 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_24_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer125 _0310_ VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1290_ _0395_ _0396_ _0580_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux2_1
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1626_ net798 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
X_1557_ net747 net705 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
X_1488_ _0538_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q VGND VGND VPWR VPWR _0546_
+ sky130_fd_sc_hd__nand2_4
X_2109_ net793 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0790_ Inst_LUT4AB_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__inv_1
XFILLER_5_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1411_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q _0500_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q
+ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1342_ net61 net89 net660 net478 Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux4_2
X_1273_ net92 net120 net108 net136 Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux4_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0988_ net72 net15 net100 net128 Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q
+ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__mux4_1
X_1609_ net766 net711 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout691 net692 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkbuf_2
Xfanout680 net681 VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1960_ net768 net679 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0911_ net75 net18 net103 net488 Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q
+ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__mux4_2
X_1891_ net39 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0842_ _0685_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop Inst_LA_LUT4c_frame_config_dffesr.c_out_mux
+ VGND VGND VPWR VPWR A sky130_fd_sc_hd__mux2_4
X_0773_ net805 net93 net121 net135 Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
+ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__mux4_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2374_ WW4END[6] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1325_ net644 _0082_ _0235_ _0649_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux4_2
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1256_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q Inst_LUT4AB_switch_matrix.JN2BEG7
+ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__nand2b_1
X_1187_ _0304_ _0303_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q VGND VGND VPWR VPWR
+ _0305_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_19_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput261 net261 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput250 Inst_LUT4AB_switch_matrix.JN2BEG4 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_8
Xoutput294 Inst_LUT4AB_switch_matrix.S1BEG0 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__buf_8
Xoutput272 net272 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput283 net283 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__buf_8
XFILLER_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1110_ net90 net116 net98 net659 Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__mux4_1
X_2090_ net765 net697 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_38_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1041_ _0166_ _0167_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VGND VGND VPWR VPWR
+ _0168_ sky130_fd_sc_hd__mux2_4
XFILLER_9_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1943_ net742 net681 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1874_ net753 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0825_ net71 net14 net99 Inst_LUT4AB_switch_matrix.JW2BEG3 Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__mux4_1
X_0756_ net634 net411 net412 net416 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__mux4_2
Xclkbuf_0_UserCLK UserCLK VGND VGND VPWR VPWR clknet_0_UserCLK sky130_fd_sc_hd__clkbuf_16
X_2357_ net132 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1308_ net414 net444 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q VGND VGND VPWR VPWR
+ _0413_ sky130_fd_sc_hd__mux2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1239_ net87 net115 net91 net660 Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
+ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__mux4_1
XFILLER_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1590_ net745 net708 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2211_ net45 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
X_2142_ Inst_LUT4AB_switch_matrix.E2BEG3 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_1
XFILLER_38_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2073_ net801 net698 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1024_ _0151_ _0058_ Inst_LC_LUT4c_frame_config_dffesr.c_I0mux VGND VGND VPWR VPWR
+ _0152_ sky130_fd_sc_hd__mux2_1
X_1926_ net773 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1857_ net785 net667 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0808_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0653_ VGND VGND VPWR VPWR _0654_
+ sky130_fd_sc_hd__and2b_1
X_1788_ net794 net733 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0739_ net805 net95 net123 net135 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_55_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1711_ net803 net727 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1642_ net44 net712 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1573_ net775 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2125_ net756 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer14 net407 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd1_1
X_2056_ net769 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer47 net442 VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_2
Xrebuffer58 net453 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_2
X_1007_ _0136_ _0135_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VGND VGND VPWR VPWR
+ _0137_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1909_ net747 net676 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_32_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer126 _0310_ VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__buf_6
XFILLER_57_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1625_ net800 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ sky130_fd_sc_hd__dlxtp_1
X_1556_ net748 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ sky130_fd_sc_hd__dlxtp_1
X_1487_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q _0529_ VGND VGND VPWR VPWR _0545_
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2108_ net795 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2039_ net742 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1410_ net89 net477 Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q VGND VGND VPWR VPWR
+ _0500_ sky130_fd_sc_hd__mux2_1
X_1341_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q _0440_ _0438_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__o211a_1
X_1272_ net62 net7 net64 net804 Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__mux4_1
XFILLER_36_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0987_ net14 net99 net127 Inst_LUT4AB_switch_matrix.JW2BEG5 Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__mux4_2
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1608_ net769 net711 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ sky130_fd_sc_hd__dlxtp_1
X_1539_ net778 net700 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout670 net671 VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__clkbuf_2
Xfanout692 FrameStrobe[2] VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__buf_2
Xfanout681 net57 VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0910_ _0045_ _0042_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.JS2BEG4 sky130_fd_sc_hd__mux2_4
X_1890_ net37 net672 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0841_ _0677_ _0684_ _0673_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__mux2_4
X_0772_ net65 net2 net81 net8 Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2373_ WW4END[5] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_2
X_1324_ net60 net88 net116 net445 Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux4_1
XFILLER_56_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1255_ _0366_ _0363_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR
+ Inst_LUT4AB_switch_matrix.JW2BEG7 sky130_fd_sc_hd__mux2_4
X_1186_ Inst_LUT4AB_switch_matrix.JN2BEG6 Inst_LUT4AB_switch_matrix.E2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q
+ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_4
XFILLER_64_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput240 net240 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput262 net262 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput251 net251 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__buf_6
Xoutput295 Inst_LUT4AB_switch_matrix.S1BEG1 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__buf_4
Xoutput284 Inst_LUT4AB_switch_matrix.NN4BEG3 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput273 net273 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1040_ net462 net628 net412 net416 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux4_1
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1942_ net744 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1873_ net758 net673 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0824_ _0665_ _0663_ _0668_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JW2BEG3 sky130_fd_sc_hd__o22a_4
X_0755_ _0594_ _0595_ _0604_ _0603_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q
+ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__mux4_2
X_2356_ net131 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__buf_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1307_ _0409_ _0410_ _0411_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q
+ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__a221o_1
X_1238_ net59 net63 net2 net24 Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__mux4_1
XFILLER_44_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1169_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 _0286_ _0287_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ _0285_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__o221a_1
XFILLER_12_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2210_ net764 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
X_2141_ Inst_LUT4AB_switch_matrix.E2BEG2 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_4
X_2072_ net741 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1023_ _0140_ _0150_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q VGND VGND VPWR VPWR
+ _0151_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1925_ net775 net675 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1856_ net787 net665 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1787_ net796 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0807_ net434 net638 net623 net643 Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__mux4_1
X_0738_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q _0587_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__o21a_1
XFILLER_57_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2339_ clknet_1_0__leaf_UserCLK VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__buf_2
XFILLER_69_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1710_ net755 net721 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1641_ net766 net715 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1572_ net776 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sky130_fd_sc_hd__dlxtp_1
X_2124_ net760 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2055_ net771 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer48 net447 VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__clkbuf_2
Xrebuffer37 Inst_LUT4AB_switch_matrix.M_EF VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__buf_6
Xrebuffer59 net454 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1006_ net60 net68 net3 net11 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__mux4_1
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1908_ net748 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_32_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer127 Inst_LUT4AB_switch_matrix.M_AB VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__buf_6
X_1839_ net803 net665 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput140 WW4END[3] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1624_ net740 net712 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.c_reset_value
+ sky130_fd_sc_hd__dlxtp_1
X_1555_ net751 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ sky130_fd_sc_hd__dlxtp_1
X_1486_ net546 _0544_ _0543_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__mux2_1
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2107_ net797 net736 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2038_ net744 net691 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1340_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__inv_1
XFILLER_68_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1271_ _0576_ _0379_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q VGND VGND VPWR VPWR
+ _0380_ sky130_fd_sc_hd__o21a_1
X_0986_ _0112_ _0114_ _0117_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.JW2BEG5 sky130_fd_sc_hd__o22a_2
X_1607_ net770 net711 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ sky130_fd_sc_hd__dlxtp_1
X_1538_ net782 net700 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ sky130_fd_sc_hd__dlxtp_1
X_1469_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q _0526_ _0528_ VGND VGND VPWR VPWR
+ _0529_ sky130_fd_sc_hd__a21oi_4
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout660 net117 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__buf_4
Xfanout671 net673 VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__clkbuf_2
Xfanout693 net694 VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__clkbuf_2
Xfanout682 net57 VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__buf_2
XFILLER_65_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0840_ _0682_ _0683_ _0650_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__mux2_1
X_0771_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _0617_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q
+ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__a21boi_2
X_2372_ WW4END[4] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_2
X_1323_ _0585_ _0420_ _0426_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W6BEG0
+ sky130_fd_sc_hd__a21o_1
X_1254_ _0364_ _0365_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VGND VGND VPWR VPWR
+ _0366_ sky130_fd_sc_hd__mux2_1
XFILLER_49_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1185_ net481 Inst_LUT4AB_switch_matrix.JW2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q
+ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_4
XFILLER_64_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0969_ _0098_ _0086_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__nand2_4
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput230 net230 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput241 net241 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput252 net252 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_4
Xoutput285 net285 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput274 net274 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput263 net263 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput296 Inst_LUT4AB_switch_matrix.S1BEG2 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__buf_8
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1941_ net746 net680 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1872_ net780 net669 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0823_ _0666_ _0667_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q VGND VGND VPWR VPWR
+ _0668_ sky130_fd_sc_hd__mux2_1
X_0754_ net83 net93 net8 net121 Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q
+ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__mux4_2
X_2355_ net130 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__buf_1
XFILLER_29_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1306_ net433 net446 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q VGND VGND VPWR VPWR
+ _0411_ sky130_fd_sc_hd__mux2_1
X_1237_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0348_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a21bo_1
X_1168_ _0282_ _0281_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__or2_4
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1099_ net78 net21 net106 net134 Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q
+ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__mux4_1
XFILLER_52_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2140_ Inst_LUT4AB_switch_matrix.E2BEG1 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_6
X_2071_ net742 net695 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ _0149_ _0148_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q VGND VGND VPWR VPWR
+ _0150_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1924_ net776 net674 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1855_ net788 net668 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1786_ net798 net732 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_0806_ _0629_ _0651_ _0605_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__mux2_4
X_0737_ _0563_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__or2_1
X_2338_ Inst_LUT4AB_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__buf_1
XFILLER_69_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1640_ net769 net713 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1571_ net778 net706 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2123_ net762 net737 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2054_ net772 net693 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer49 net481 VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__buf_6
Xrebuffer38 H VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__buf_6
X_1005_ net88 net96 net116 net659 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__mux4_1
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1907_ net750 net678 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer128 _0335_ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd1_1
X_1838_ net755 net664 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1769_ net767 net731 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput130 W2MID[3] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1623_ net743 net55 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.c_I0mux
+ sky130_fd_sc_hd__dlxtp_1
X_1554_ net752 net704 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ sky130_fd_sc_hd__dlxtp_1
X_1485_ Inst_LA_LUT4c_frame_config_dffesr.c_reset_value _0685_ _0542_ VGND VGND VPWR
+ VPWR _0544_ sky130_fd_sc_hd__mux2_2
.ends

