module S_term_single2 (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 sky130_fd_sc_hd__clkbuf_2 _000_ (.A(FrameData[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 _001_ (.A(FrameData[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 _002_ (.A(FrameData[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 _003_ (.A(FrameData[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 _004_ (.A(FrameData[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 _005_ (.A(FrameData[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 _006_ (.A(FrameData[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 _007_ (.A(FrameData[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 _008_ (.A(FrameData[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 _009_ (.A(FrameData[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 _010_ (.A(FrameData[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 _011_ (.A(FrameData[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 _012_ (.A(FrameData[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 _013_ (.A(FrameData[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 _014_ (.A(FrameData[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 _015_ (.A(FrameData[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 _016_ (.A(FrameData[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 _017_ (.A(FrameData[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 _018_ (.A(FrameData[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 _019_ (.A(FrameData[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 _020_ (.A(FrameData[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 _021_ (.A(FrameData[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 _022_ (.A(FrameData[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 _023_ (.A(FrameData[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 _024_ (.A(FrameData[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 _025_ (.A(FrameData[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 _026_ (.A(FrameData[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 _027_ (.A(FrameData[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 _028_ (.A(FrameData[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 _029_ (.A(FrameData[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 _030_ (.A(FrameData[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 _031_ (.A(FrameData[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 _032_ (.A(FrameStrobe[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 _033_ (.A(FrameStrobe[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 _034_ (.A(FrameStrobe[2]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 _035_ (.A(FrameStrobe[3]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 _036_ (.A(FrameStrobe[4]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 _037_ (.A(FrameStrobe[5]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 _038_ (.A(FrameStrobe[6]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 _039_ (.A(FrameStrobe[7]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _040_ (.A(FrameStrobe[8]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 _041_ (.A(FrameStrobe[9]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 _042_ (.A(FrameStrobe[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 _043_ (.A(FrameStrobe[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 _044_ (.A(FrameStrobe[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 _045_ (.A(FrameStrobe[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 _046_ (.A(FrameStrobe[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 _047_ (.A(FrameStrobe[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 _048_ (.A(FrameStrobe[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 _049_ (.A(FrameStrobe[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 _050_ (.A(FrameStrobe[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _051_ (.A(FrameStrobe[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 _052_ (.A(S1END[3]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 _053_ (.A(S1END[2]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 _054_ (.A(S1END[1]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 _055_ (.A(S1END[0]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 _056_ (.A(S2MID[7]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 _057_ (.A(S2MID[6]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 _058_ (.A(S2MID[5]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 _059_ (.A(S2MID[4]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 _060_ (.A(S2MID[3]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 _061_ (.A(S2MID[2]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 _062_ (.A(S2MID[1]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 _063_ (.A(S2MID[0]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 _064_ (.A(S2END[7]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 _065_ (.A(S2END[6]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 _066_ (.A(S2END[5]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 _067_ (.A(S2END[4]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _068_ (.A(S2END[3]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 _069_ (.A(S2END[2]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 _070_ (.A(S2END[1]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 _071_ (.A(S2END[0]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 _072_ (.A(S4END[15]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 _073_ (.A(S4END[14]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 _074_ (.A(S4END[13]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 _075_ (.A(S4END[12]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 _076_ (.A(S4END[11]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 _077_ (.A(S4END[10]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 _078_ (.A(S4END[9]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 _079_ (.A(S4END[8]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 _080_ (.A(S4END[7]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 _081_ (.A(S4END[6]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 _082_ (.A(S4END[5]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 _083_ (.A(S4END[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _084_ (.A(S4END[3]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _085_ (.A(S4END[2]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _086_ (.A(S4END[1]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 _087_ (.A(S4END[0]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(SS4END[15]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(SS4END[14]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _090_ (.A(SS4END[13]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _091_ (.A(SS4END[12]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _092_ (.A(SS4END[11]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _093_ (.A(SS4END[10]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _094_ (.A(SS4END[9]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _095_ (.A(SS4END[8]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(SS4END[7]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _097_ (.A(SS4END[6]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 _098_ (.A(SS4END[5]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _099_ (.A(SS4END[4]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 _100_ (.A(SS4END[3]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 _101_ (.A(SS4END[2]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 _102_ (.A(SS4END[1]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 _103_ (.A(SS4END[0]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 _104_ (.A(UserCLK),
    .X(net105));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_135 ();
 sky130_fd_sc_hd__buf_2 output1 (.A(net1),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(UserCLKo));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(FrameData[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameData[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(FrameData[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(FrameData[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(FrameData[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameData[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(FrameData[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(FrameData[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(FrameData[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(FrameData[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(FrameData[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(FrameData[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(FrameData[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(FrameData[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(FrameData[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(FrameData[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(FrameData[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(FrameData[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(FrameData[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(FrameData[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(FrameData[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(FrameData[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(FrameData[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(FrameData[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(FrameData[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(S4END[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(S4END[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(SS4END[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(SS4END[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(SS4END[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(SS4END[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(SS4END[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(SS4END[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(SS4END[15]));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
endmodule
