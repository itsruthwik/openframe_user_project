magic
tech sky130A
magscale 1 2
timestamp 1746536547
<< viali >>
rect 1501 42313 1535 42347
rect 1961 42313 1995 42347
rect 2421 42313 2455 42347
rect 2789 42313 2823 42347
rect 3065 42313 3099 42347
rect 3433 42313 3467 42347
rect 4261 42313 4295 42347
rect 4629 42313 4663 42347
rect 5181 42313 5215 42347
rect 5549 42313 5583 42347
rect 6101 42313 6135 42347
rect 6561 42313 6595 42347
rect 7021 42313 7055 42347
rect 7481 42313 7515 42347
rect 7941 42313 7975 42347
rect 8309 42313 8343 42347
rect 1685 42177 1719 42211
rect 1777 42177 1811 42211
rect 2237 42177 2271 42211
rect 2605 42177 2639 42211
rect 3249 42177 3283 42211
rect 3617 42177 3651 42211
rect 4077 42177 4111 42211
rect 4813 42177 4847 42211
rect 4997 42177 5031 42211
rect 5733 42177 5767 42211
rect 5917 42177 5951 42211
rect 6377 42177 6411 42211
rect 6837 42177 6871 42211
rect 7297 42177 7331 42211
rect 7757 42177 7791 42211
rect 8125 42177 8159 42211
rect 1777 41769 1811 41803
rect 8309 41769 8343 41803
rect 1501 41701 1535 41735
rect 7941 41701 7975 41735
rect 1685 41565 1719 41599
rect 1961 41565 1995 41599
rect 7481 41565 7515 41599
rect 7757 41565 7791 41599
rect 8125 41565 8159 41599
rect 7665 41429 7699 41463
rect 8309 41225 8343 41259
rect 7941 41089 7975 41123
rect 8125 41089 8159 41123
rect 7757 40885 7791 40919
rect 2053 40477 2087 40511
rect 7665 40477 7699 40511
rect 2237 40341 2271 40375
rect 7849 40341 7883 40375
rect 7757 40001 7791 40035
rect 8125 40001 8159 40035
rect 7941 39865 7975 39899
rect 8309 39797 8343 39831
rect 2789 39389 2823 39423
rect 7481 39389 7515 39423
rect 7757 39389 7791 39423
rect 8125 39389 8159 39423
rect 2973 39253 3007 39287
rect 7665 39253 7699 39287
rect 7941 39253 7975 39287
rect 8309 39253 8343 39287
rect 7757 38913 7791 38947
rect 8125 38913 8159 38947
rect 7941 38777 7975 38811
rect 8309 38709 8343 38743
rect 7665 38505 7699 38539
rect 2697 38301 2731 38335
rect 7481 38301 7515 38335
rect 7757 38301 7791 38335
rect 8125 38301 8159 38335
rect 2881 38165 2915 38199
rect 7941 38165 7975 38199
rect 8309 38165 8343 38199
rect 7665 37961 7699 37995
rect 7481 37825 7515 37859
rect 7757 37825 7791 37859
rect 8125 37825 8159 37859
rect 7941 37689 7975 37723
rect 8309 37621 8343 37655
rect 7665 37417 7699 37451
rect 7481 37213 7515 37247
rect 7757 37213 7791 37247
rect 8125 37213 8159 37247
rect 7941 37077 7975 37111
rect 8309 37077 8343 37111
rect 2605 36873 2639 36907
rect 2421 36737 2455 36771
rect 7757 36737 7791 36771
rect 8125 36737 8159 36771
rect 7941 36601 7975 36635
rect 8309 36533 8343 36567
rect 2237 36261 2271 36295
rect 2053 36125 2087 36159
rect 7757 36125 7791 36159
rect 8125 36125 8159 36159
rect 7941 35989 7975 36023
rect 8309 35989 8343 36023
rect 7757 35649 7791 35683
rect 8125 35649 8159 35683
rect 7941 35513 7975 35547
rect 8309 35445 8343 35479
rect 1777 35241 1811 35275
rect 7665 35241 7699 35275
rect 1593 35037 1627 35071
rect 7481 35037 7515 35071
rect 7757 35037 7791 35071
rect 8125 35037 8159 35071
rect 7941 34901 7975 34935
rect 8309 34901 8343 34935
rect 7941 34697 7975 34731
rect 7757 34561 7791 34595
rect 8125 34561 8159 34595
rect 8309 34357 8343 34391
rect 2053 33949 2087 33983
rect 7757 33949 7791 33983
rect 8125 33949 8159 33983
rect 2237 33813 2271 33847
rect 7941 33813 7975 33847
rect 8309 33813 8343 33847
rect 1869 33609 1903 33643
rect 1685 33473 1719 33507
rect 7757 33473 7791 33507
rect 8125 33473 8159 33507
rect 7941 33337 7975 33371
rect 8309 33269 8343 33303
rect 2605 33065 2639 33099
rect 2421 32861 2455 32895
rect 7481 32861 7515 32895
rect 7757 32861 7791 32895
rect 8125 32861 8159 32895
rect 7665 32725 7699 32759
rect 7941 32725 7975 32759
rect 8309 32725 8343 32759
rect 2789 32521 2823 32555
rect 2605 32385 2639 32419
rect 7757 32385 7791 32419
rect 8125 32385 8159 32419
rect 7941 32249 7975 32283
rect 8309 32181 8343 32215
rect 2973 31977 3007 32011
rect 7941 31909 7975 31943
rect 2789 31773 2823 31807
rect 7205 31773 7239 31807
rect 7757 31773 7791 31807
rect 8125 31773 8159 31807
rect 7389 31637 7423 31671
rect 8309 31637 8343 31671
rect 2237 31433 2271 31467
rect 2053 31297 2087 31331
rect 7757 31297 7791 31331
rect 8125 31297 8159 31331
rect 7941 31161 7975 31195
rect 2789 31093 2823 31127
rect 8309 31093 8343 31127
rect 7021 30685 7055 30719
rect 7757 30685 7791 30719
rect 8125 30685 8159 30719
rect 7205 30549 7239 30583
rect 7941 30549 7975 30583
rect 8309 30549 8343 30583
rect 1593 30209 1627 30243
rect 2605 30209 2639 30243
rect 7113 30209 7147 30243
rect 7757 30209 7791 30243
rect 8125 30209 8159 30243
rect 1777 30073 1811 30107
rect 7941 30073 7975 30107
rect 2789 30005 2823 30039
rect 7297 30005 7331 30039
rect 8309 30005 8343 30039
rect 7297 29597 7331 29631
rect 7757 29597 7791 29631
rect 8125 29597 8159 29631
rect 7481 29461 7515 29495
rect 7941 29461 7975 29495
rect 8309 29461 8343 29495
rect 2697 29257 2731 29291
rect 7297 29257 7331 29291
rect 2513 29121 2547 29155
rect 7113 29121 7147 29155
rect 7757 29121 7791 29155
rect 8125 29121 8159 29155
rect 7941 28985 7975 29019
rect 8309 28917 8343 28951
rect 7665 28713 7699 28747
rect 7481 28509 7515 28543
rect 7757 28509 7791 28543
rect 8125 28509 8159 28543
rect 7941 28373 7975 28407
rect 8309 28373 8343 28407
rect 7665 28169 7699 28203
rect 7481 28033 7515 28067
rect 7757 28033 7791 28067
rect 8125 28033 8159 28067
rect 7941 27897 7975 27931
rect 8309 27829 8343 27863
rect 7665 27625 7699 27659
rect 2605 27557 2639 27591
rect 2421 27421 2455 27455
rect 7481 27421 7515 27455
rect 7757 27421 7791 27455
rect 8125 27421 8159 27455
rect 7941 27285 7975 27319
rect 8309 27285 8343 27319
rect 7481 27081 7515 27115
rect 7297 26945 7331 26979
rect 7757 26945 7791 26979
rect 8125 26945 8159 26979
rect 7941 26809 7975 26843
rect 8309 26741 8343 26775
rect 7205 26537 7239 26571
rect 7389 26469 7423 26503
rect 7849 26469 7883 26503
rect 7021 26333 7055 26367
rect 8033 26333 8067 26367
rect 8125 26333 8159 26367
rect 7297 26265 7331 26299
rect 8309 26197 8343 26231
rect 2145 25993 2179 26027
rect 3157 25993 3191 26027
rect 7205 25993 7239 26027
rect 1961 25857 1995 25891
rect 2973 25857 3007 25891
rect 7021 25857 7055 25891
rect 7757 25857 7791 25891
rect 8125 25857 8159 25891
rect 7941 25721 7975 25755
rect 8309 25653 8343 25687
rect 1869 25449 1903 25483
rect 7389 25449 7423 25483
rect 1685 25245 1719 25279
rect 7205 25245 7239 25279
rect 7757 25245 7791 25279
rect 8125 25245 8159 25279
rect 3065 25177 3099 25211
rect 7941 25109 7975 25143
rect 8309 25109 8343 25143
rect 7021 24769 7055 24803
rect 7297 24769 7331 24803
rect 7757 24769 7791 24803
rect 8125 24769 8159 24803
rect 7205 24633 7239 24667
rect 7481 24633 7515 24667
rect 7941 24565 7975 24599
rect 8309 24565 8343 24599
rect 3433 24361 3467 24395
rect 5089 24361 5123 24395
rect 7665 24361 7699 24395
rect 3617 24157 3651 24191
rect 4905 24157 4939 24191
rect 7481 24157 7515 24191
rect 7757 24157 7791 24191
rect 8125 24157 8159 24191
rect 7021 24089 7055 24123
rect 7941 24021 7975 24055
rect 8309 24021 8343 24055
rect 1777 23817 1811 23851
rect 1961 23681 1995 23715
rect 7757 23681 7791 23715
rect 8125 23681 8159 23715
rect 7941 23545 7975 23579
rect 4997 23477 5031 23511
rect 8309 23477 8343 23511
rect 7665 23273 7699 23307
rect 7481 23069 7515 23103
rect 7757 23069 7791 23103
rect 8125 23069 8159 23103
rect 7941 22933 7975 22967
rect 8309 22933 8343 22967
rect 3801 22729 3835 22763
rect 7205 22729 7239 22763
rect 7573 22729 7607 22763
rect 1869 22593 1903 22627
rect 3617 22593 3651 22627
rect 7021 22593 7055 22627
rect 7757 22593 7791 22627
rect 8125 22593 8159 22627
rect 2053 22457 2087 22491
rect 7941 22389 7975 22423
rect 8309 22389 8343 22423
rect 7113 22117 7147 22151
rect 4537 21981 4571 22015
rect 6745 21981 6779 22015
rect 7297 21981 7331 22015
rect 7757 21981 7791 22015
rect 8125 21981 8159 22015
rect 4721 21845 4755 21879
rect 6929 21845 6963 21879
rect 7481 21845 7515 21879
rect 7941 21845 7975 21879
rect 8309 21845 8343 21879
rect 1777 21641 1811 21675
rect 7389 21641 7423 21675
rect 1593 21505 1627 21539
rect 7757 21505 7791 21539
rect 8125 21505 8159 21539
rect 3709 21301 3743 21335
rect 7297 21301 7331 21335
rect 7941 21301 7975 21335
rect 8309 21301 8343 21335
rect 6929 21097 6963 21131
rect 7941 21029 7975 21063
rect 6745 20893 6779 20927
rect 7757 20893 7791 20927
rect 8125 20893 8159 20927
rect 8309 20757 8343 20791
rect 5273 20553 5307 20587
rect 5549 20553 5583 20587
rect 5089 20417 5123 20451
rect 5365 20417 5399 20451
rect 7757 20417 7791 20451
rect 8125 20417 8159 20451
rect 7941 20213 7975 20247
rect 8309 20213 8343 20247
rect 2605 20009 2639 20043
rect 4905 20009 4939 20043
rect 2421 19805 2455 19839
rect 4721 19805 4755 19839
rect 7757 19805 7791 19839
rect 8125 19805 8159 19839
rect 7941 19669 7975 19703
rect 8309 19669 8343 19703
rect 1869 19465 1903 19499
rect 3525 19465 3559 19499
rect 3617 19465 3651 19499
rect 6653 19465 6687 19499
rect 7665 19465 7699 19499
rect 7849 19465 7883 19499
rect 8309 19465 8343 19499
rect 1685 19329 1719 19363
rect 3341 19329 3375 19363
rect 3801 19329 3835 19363
rect 6469 19329 6503 19363
rect 7481 19329 7515 19363
rect 8033 19329 8067 19363
rect 8125 19329 8159 19363
rect 7297 18921 7331 18955
rect 7665 18921 7699 18955
rect 7113 18717 7147 18751
rect 7481 18717 7515 18751
rect 7757 18717 7791 18751
rect 8125 18717 8159 18751
rect 7941 18581 7975 18615
rect 8309 18581 8343 18615
rect 4813 18377 4847 18411
rect 7389 18377 7423 18411
rect 4629 18241 4663 18275
rect 7205 18241 7239 18275
rect 1777 17833 1811 17867
rect 6837 17833 6871 17867
rect 1593 17629 1627 17663
rect 6653 17629 6687 17663
rect 7113 17289 7147 17323
rect 6929 17153 6963 17187
rect 1869 16201 1903 16235
rect 4905 16201 4939 16235
rect 6561 16201 6595 16235
rect 7573 16201 7607 16235
rect 2053 16065 2087 16099
rect 4721 16065 4755 16099
rect 6377 16065 6411 16099
rect 7389 16065 7423 16099
rect 2237 15657 2271 15691
rect 2053 15453 2087 15487
rect 6561 15113 6595 15147
rect 6377 14977 6411 15011
rect 2145 14569 2179 14603
rect 6929 14569 6963 14603
rect 8125 14569 8159 14603
rect 1961 14365 1995 14399
rect 6745 14365 6779 14399
rect 7941 14365 7975 14399
rect 1869 13481 1903 13515
rect 8033 13481 8067 13515
rect 1685 13277 1719 13311
rect 7849 13277 7883 13311
rect 5917 12393 5951 12427
rect 7665 12393 7699 12427
rect 5733 12189 5767 12223
rect 7481 12189 7515 12223
rect 7849 11849 7883 11883
rect 8033 11713 8067 11747
rect 1869 11305 1903 11339
rect 5825 11305 5859 11339
rect 2053 11101 2087 11135
rect 5641 11101 5675 11135
rect 6929 10761 6963 10795
rect 6745 10625 6779 10659
rect 6929 9537 6963 9571
rect 7113 9401 7147 9435
rect 7297 9129 7331 9163
rect 7113 8925 7147 8959
rect 6561 8585 6595 8619
rect 6377 8449 6411 8483
rect 7205 8041 7239 8075
rect 7021 7837 7055 7871
rect 7941 6749 7975 6783
rect 7757 6613 7791 6647
rect 7389 6409 7423 6443
rect 7205 6273 7239 6307
rect 6009 5865 6043 5899
rect 5825 5661 5859 5695
rect 6193 4777 6227 4811
rect 6009 4573 6043 4607
rect 7297 4097 7331 4131
rect 7481 3961 7515 3995
rect 7941 3689 7975 3723
rect 8125 3485 8159 3519
rect 6101 3145 6135 3179
rect 6561 3145 6595 3179
rect 5917 3009 5951 3043
rect 6377 3009 6411 3043
rect 7849 3009 7883 3043
rect 8033 2873 8067 2907
<< metal1 >>
rect 1104 42458 8740 42480
rect 1104 42406 3010 42458
rect 3062 42406 3074 42458
rect 3126 42406 3138 42458
rect 3190 42406 3202 42458
rect 3254 42406 3266 42458
rect 3318 42406 8740 42458
rect 1104 42384 8740 42406
rect 1210 42304 1216 42356
rect 1268 42344 1274 42356
rect 1489 42347 1547 42353
rect 1489 42344 1501 42347
rect 1268 42316 1501 42344
rect 1268 42304 1274 42316
rect 1489 42313 1501 42316
rect 1535 42313 1547 42347
rect 1489 42307 1547 42313
rect 1670 42304 1676 42356
rect 1728 42344 1734 42356
rect 1949 42347 2007 42353
rect 1949 42344 1961 42347
rect 1728 42316 1961 42344
rect 1728 42304 1734 42316
rect 1949 42313 1961 42316
rect 1995 42313 2007 42347
rect 1949 42307 2007 42313
rect 2130 42304 2136 42356
rect 2188 42344 2194 42356
rect 2409 42347 2467 42353
rect 2409 42344 2421 42347
rect 2188 42316 2421 42344
rect 2188 42304 2194 42316
rect 2409 42313 2421 42316
rect 2455 42313 2467 42347
rect 2409 42307 2467 42313
rect 2590 42304 2596 42356
rect 2648 42344 2654 42356
rect 2777 42347 2835 42353
rect 2777 42344 2789 42347
rect 2648 42316 2789 42344
rect 2648 42304 2654 42316
rect 2777 42313 2789 42316
rect 2823 42313 2835 42347
rect 2777 42307 2835 42313
rect 2866 42304 2872 42356
rect 2924 42344 2930 42356
rect 3053 42347 3111 42353
rect 3053 42344 3065 42347
rect 2924 42316 3065 42344
rect 2924 42304 2930 42316
rect 3053 42313 3065 42316
rect 3099 42313 3111 42347
rect 3053 42307 3111 42313
rect 3421 42347 3479 42353
rect 3421 42313 3433 42347
rect 3467 42344 3479 42347
rect 3510 42344 3516 42356
rect 3467 42316 3516 42344
rect 3467 42313 3479 42316
rect 3421 42307 3479 42313
rect 3510 42304 3516 42316
rect 3568 42304 3574 42356
rect 3970 42304 3976 42356
rect 4028 42344 4034 42356
rect 4249 42347 4307 42353
rect 4249 42344 4261 42347
rect 4028 42316 4261 42344
rect 4028 42304 4034 42316
rect 4249 42313 4261 42316
rect 4295 42313 4307 42347
rect 4249 42307 4307 42313
rect 4430 42304 4436 42356
rect 4488 42344 4494 42356
rect 4617 42347 4675 42353
rect 4617 42344 4629 42347
rect 4488 42316 4629 42344
rect 4488 42304 4494 42316
rect 4617 42313 4629 42316
rect 4663 42313 4675 42347
rect 4617 42307 4675 42313
rect 4890 42304 4896 42356
rect 4948 42344 4954 42356
rect 5169 42347 5227 42353
rect 5169 42344 5181 42347
rect 4948 42316 5181 42344
rect 4948 42304 4954 42316
rect 5169 42313 5181 42316
rect 5215 42313 5227 42347
rect 5169 42307 5227 42313
rect 5350 42304 5356 42356
rect 5408 42344 5414 42356
rect 5537 42347 5595 42353
rect 5537 42344 5549 42347
rect 5408 42316 5549 42344
rect 5408 42304 5414 42316
rect 5537 42313 5549 42316
rect 5583 42313 5595 42347
rect 5537 42307 5595 42313
rect 5810 42304 5816 42356
rect 5868 42344 5874 42356
rect 6089 42347 6147 42353
rect 6089 42344 6101 42347
rect 5868 42316 6101 42344
rect 5868 42304 5874 42316
rect 6089 42313 6101 42316
rect 6135 42313 6147 42347
rect 6089 42307 6147 42313
rect 6270 42304 6276 42356
rect 6328 42344 6334 42356
rect 6549 42347 6607 42353
rect 6549 42344 6561 42347
rect 6328 42316 6561 42344
rect 6328 42304 6334 42316
rect 6549 42313 6561 42316
rect 6595 42313 6607 42347
rect 6549 42307 6607 42313
rect 6730 42304 6736 42356
rect 6788 42344 6794 42356
rect 7009 42347 7067 42353
rect 7009 42344 7021 42347
rect 6788 42316 7021 42344
rect 6788 42304 6794 42316
rect 7009 42313 7021 42316
rect 7055 42313 7067 42347
rect 7009 42307 7067 42313
rect 7190 42304 7196 42356
rect 7248 42344 7254 42356
rect 7469 42347 7527 42353
rect 7469 42344 7481 42347
rect 7248 42316 7481 42344
rect 7248 42304 7254 42316
rect 7469 42313 7481 42316
rect 7515 42313 7527 42347
rect 7469 42307 7527 42313
rect 7650 42304 7656 42356
rect 7708 42344 7714 42356
rect 7929 42347 7987 42353
rect 7929 42344 7941 42347
rect 7708 42316 7941 42344
rect 7708 42304 7714 42316
rect 7929 42313 7941 42316
rect 7975 42313 7987 42347
rect 7929 42307 7987 42313
rect 8110 42304 8116 42356
rect 8168 42344 8174 42356
rect 8297 42347 8355 42353
rect 8297 42344 8309 42347
rect 8168 42316 8309 42344
rect 8168 42304 8174 42316
rect 8297 42313 8309 42316
rect 8343 42313 8355 42347
rect 8297 42307 8355 42313
rect 4522 42236 4528 42288
rect 4580 42276 4586 42288
rect 4580 42248 6868 42276
rect 4580 42236 4586 42248
rect 1670 42168 1676 42220
rect 1728 42168 1734 42220
rect 1765 42211 1823 42217
rect 1765 42177 1777 42211
rect 1811 42177 1823 42211
rect 1765 42171 1823 42177
rect 2225 42211 2283 42217
rect 2225 42177 2237 42211
rect 2271 42177 2283 42211
rect 2225 42171 2283 42177
rect 1578 42100 1584 42152
rect 1636 42140 1642 42152
rect 1780 42140 1808 42171
rect 1636 42112 1808 42140
rect 2240 42140 2268 42171
rect 2590 42168 2596 42220
rect 2648 42168 2654 42220
rect 3237 42211 3295 42217
rect 3237 42177 3249 42211
rect 3283 42208 3295 42211
rect 3418 42208 3424 42220
rect 3283 42180 3424 42208
rect 3283 42177 3295 42180
rect 3237 42171 3295 42177
rect 3418 42168 3424 42180
rect 3476 42168 3482 42220
rect 3602 42168 3608 42220
rect 3660 42168 3666 42220
rect 3786 42168 3792 42220
rect 3844 42208 3850 42220
rect 4065 42211 4123 42217
rect 4065 42208 4077 42211
rect 3844 42180 4077 42208
rect 3844 42168 3850 42180
rect 4065 42177 4077 42180
rect 4111 42177 4123 42211
rect 4065 42171 4123 42177
rect 4801 42211 4859 42217
rect 4801 42177 4813 42211
rect 4847 42208 4859 42211
rect 4890 42208 4896 42220
rect 4847 42180 4896 42208
rect 4847 42177 4859 42180
rect 4801 42171 4859 42177
rect 4890 42168 4896 42180
rect 4948 42168 4954 42220
rect 4982 42168 4988 42220
rect 5040 42168 5046 42220
rect 5626 42168 5632 42220
rect 5684 42208 5690 42220
rect 5721 42211 5779 42217
rect 5721 42208 5733 42211
rect 5684 42180 5733 42208
rect 5684 42168 5690 42180
rect 5721 42177 5733 42180
rect 5767 42177 5779 42211
rect 5721 42171 5779 42177
rect 5902 42168 5908 42220
rect 5960 42168 5966 42220
rect 6840 42217 6868 42248
rect 7024 42248 8156 42276
rect 7024 42220 7052 42248
rect 6365 42211 6423 42217
rect 6365 42177 6377 42211
rect 6411 42177 6423 42211
rect 6365 42171 6423 42177
rect 6825 42211 6883 42217
rect 6825 42177 6837 42211
rect 6871 42177 6883 42211
rect 6825 42171 6883 42177
rect 2682 42140 2688 42152
rect 2240 42112 2688 42140
rect 1636 42100 1642 42112
rect 2682 42100 2688 42112
rect 2740 42100 2746 42152
rect 4706 42100 4712 42152
rect 4764 42140 4770 42152
rect 6380 42140 6408 42171
rect 7006 42168 7012 42220
rect 7064 42168 7070 42220
rect 8128 42217 8156 42248
rect 7285 42211 7343 42217
rect 7285 42177 7297 42211
rect 7331 42177 7343 42211
rect 7285 42171 7343 42177
rect 7745 42211 7803 42217
rect 7745 42177 7757 42211
rect 7791 42177 7803 42211
rect 7745 42171 7803 42177
rect 8113 42211 8171 42217
rect 8113 42177 8125 42211
rect 8159 42177 8171 42211
rect 8113 42171 8171 42177
rect 4764 42112 6408 42140
rect 4764 42100 4770 42112
rect 5442 42032 5448 42084
rect 5500 42072 5506 42084
rect 7300 42072 7328 42171
rect 5500 42044 7328 42072
rect 5500 42032 5506 42044
rect 5074 41964 5080 42016
rect 5132 42004 5138 42016
rect 7760 42004 7788 42171
rect 5132 41976 7788 42004
rect 5132 41964 5138 41976
rect 1104 41914 8740 41936
rect 1104 41862 1950 41914
rect 2002 41862 2014 41914
rect 2066 41862 2078 41914
rect 2130 41862 2142 41914
rect 2194 41862 2206 41914
rect 2258 41862 7950 41914
rect 8002 41862 8014 41914
rect 8066 41862 8078 41914
rect 8130 41862 8142 41914
rect 8194 41862 8206 41914
rect 8258 41862 8740 41914
rect 1104 41840 8740 41862
rect 290 41760 296 41812
rect 348 41800 354 41812
rect 1765 41803 1823 41809
rect 1765 41800 1777 41803
rect 348 41772 1777 41800
rect 348 41760 354 41772
rect 1765 41769 1777 41772
rect 1811 41769 1823 41803
rect 1765 41763 1823 41769
rect 8297 41803 8355 41809
rect 8297 41769 8309 41803
rect 8343 41800 8355 41803
rect 8570 41800 8576 41812
rect 8343 41772 8576 41800
rect 8343 41769 8355 41772
rect 8297 41763 8355 41769
rect 8570 41760 8576 41772
rect 8628 41760 8634 41812
rect 750 41692 756 41744
rect 808 41732 814 41744
rect 1489 41735 1547 41741
rect 1489 41732 1501 41735
rect 808 41704 1501 41732
rect 808 41692 814 41704
rect 1489 41701 1501 41704
rect 1535 41701 1547 41735
rect 1489 41695 1547 41701
rect 7929 41735 7987 41741
rect 7929 41701 7941 41735
rect 7975 41732 7987 41735
rect 9030 41732 9036 41744
rect 7975 41704 9036 41732
rect 7975 41701 7987 41704
rect 7929 41695 7987 41701
rect 9030 41692 9036 41704
rect 9088 41692 9094 41744
rect 6086 41624 6092 41676
rect 6144 41664 6150 41676
rect 6144 41636 8156 41664
rect 6144 41624 6150 41636
rect 1670 41556 1676 41608
rect 1728 41556 1734 41608
rect 1854 41556 1860 41608
rect 1912 41596 1918 41608
rect 1949 41599 2007 41605
rect 1949 41596 1961 41599
rect 1912 41568 1961 41596
rect 1912 41556 1918 41568
rect 1949 41565 1961 41568
rect 1995 41565 2007 41599
rect 1949 41559 2007 41565
rect 7466 41556 7472 41608
rect 7524 41556 7530 41608
rect 8128 41605 8156 41636
rect 7745 41599 7803 41605
rect 7745 41565 7757 41599
rect 7791 41565 7803 41599
rect 7745 41559 7803 41565
rect 8113 41599 8171 41605
rect 8113 41565 8125 41599
rect 8159 41565 8171 41599
rect 8113 41559 8171 41565
rect 7098 41488 7104 41540
rect 7156 41528 7162 41540
rect 7760 41528 7788 41559
rect 7156 41500 7788 41528
rect 7156 41488 7162 41500
rect 7653 41463 7711 41469
rect 7653 41429 7665 41463
rect 7699 41460 7711 41463
rect 7834 41460 7840 41472
rect 7699 41432 7840 41460
rect 7699 41429 7711 41432
rect 7653 41423 7711 41429
rect 7834 41420 7840 41432
rect 7892 41420 7898 41472
rect 1104 41370 8740 41392
rect 1104 41318 3010 41370
rect 3062 41318 3074 41370
rect 3126 41318 3138 41370
rect 3190 41318 3202 41370
rect 3254 41318 3266 41370
rect 3318 41318 8740 41370
rect 1104 41296 8740 41318
rect 8297 41259 8355 41265
rect 8297 41225 8309 41259
rect 8343 41256 8355 41259
rect 9490 41256 9496 41268
rect 8343 41228 9496 41256
rect 8343 41225 8355 41228
rect 8297 41219 8355 41225
rect 9490 41216 9496 41228
rect 9548 41216 9554 41268
rect 7374 41080 7380 41132
rect 7432 41120 7438 41132
rect 7929 41123 7987 41129
rect 7929 41120 7941 41123
rect 7432 41092 7941 41120
rect 7432 41080 7438 41092
rect 7929 41089 7941 41092
rect 7975 41089 7987 41123
rect 7929 41083 7987 41089
rect 8113 41123 8171 41129
rect 8113 41089 8125 41123
rect 8159 41089 8171 41123
rect 8113 41083 8171 41089
rect 6730 41012 6736 41064
rect 6788 41052 6794 41064
rect 8128 41052 8156 41083
rect 6788 41024 8156 41052
rect 6788 41012 6794 41024
rect 7742 40876 7748 40928
rect 7800 40876 7806 40928
rect 1104 40826 8740 40848
rect 1104 40774 1950 40826
rect 2002 40774 2014 40826
rect 2066 40774 2078 40826
rect 2130 40774 2142 40826
rect 2194 40774 2206 40826
rect 2258 40774 7950 40826
rect 8002 40774 8014 40826
rect 8066 40774 8078 40826
rect 8130 40774 8142 40826
rect 8194 40774 8206 40826
rect 8258 40774 8740 40826
rect 1104 40752 8740 40774
rect 198 40468 204 40520
rect 256 40508 262 40520
rect 2041 40511 2099 40517
rect 2041 40508 2053 40511
rect 256 40480 2053 40508
rect 256 40468 262 40480
rect 2041 40477 2053 40480
rect 2087 40477 2099 40511
rect 2041 40471 2099 40477
rect 7650 40468 7656 40520
rect 7708 40468 7714 40520
rect 2225 40375 2283 40381
rect 2225 40341 2237 40375
rect 2271 40372 2283 40375
rect 5718 40372 5724 40384
rect 2271 40344 5724 40372
rect 2271 40341 2283 40344
rect 2225 40335 2283 40341
rect 5718 40332 5724 40344
rect 5776 40332 5782 40384
rect 7834 40332 7840 40384
rect 7892 40332 7898 40384
rect 1104 40282 8740 40304
rect 1104 40230 3010 40282
rect 3062 40230 3074 40282
rect 3126 40230 3138 40282
rect 3190 40230 3202 40282
rect 3254 40230 3266 40282
rect 3318 40230 8740 40282
rect 1104 40208 8740 40230
rect 7926 40060 7932 40112
rect 7984 40100 7990 40112
rect 7984 40072 8156 40100
rect 7984 40060 7990 40072
rect 7742 39992 7748 40044
rect 7800 39992 7806 40044
rect 8128 40041 8156 40072
rect 8113 40035 8171 40041
rect 8113 40001 8125 40035
rect 8159 40001 8171 40035
rect 8113 39995 8171 40001
rect 7926 39856 7932 39908
rect 7984 39856 7990 39908
rect 8294 39788 8300 39840
rect 8352 39788 8358 39840
rect 1104 39738 8740 39760
rect 1104 39686 1950 39738
rect 2002 39686 2014 39738
rect 2066 39686 2078 39738
rect 2130 39686 2142 39738
rect 2194 39686 2206 39738
rect 2258 39686 7950 39738
rect 8002 39686 8014 39738
rect 8066 39686 8078 39738
rect 8130 39686 8142 39738
rect 8194 39686 8206 39738
rect 8258 39686 8740 39738
rect 1104 39664 8740 39686
rect 106 39380 112 39432
rect 164 39420 170 39432
rect 2777 39423 2835 39429
rect 2777 39420 2789 39423
rect 164 39392 2789 39420
rect 164 39380 170 39392
rect 2777 39389 2789 39392
rect 2823 39389 2835 39423
rect 2777 39383 2835 39389
rect 5534 39380 5540 39432
rect 5592 39420 5598 39432
rect 7469 39423 7527 39429
rect 7469 39420 7481 39423
rect 5592 39392 7481 39420
rect 5592 39380 5598 39392
rect 7469 39389 7481 39392
rect 7515 39389 7527 39423
rect 7469 39383 7527 39389
rect 7745 39423 7803 39429
rect 7745 39389 7757 39423
rect 7791 39420 7803 39423
rect 7834 39420 7840 39432
rect 7791 39392 7840 39420
rect 7791 39389 7803 39392
rect 7745 39383 7803 39389
rect 7834 39380 7840 39392
rect 7892 39380 7898 39432
rect 8113 39423 8171 39429
rect 8113 39389 8125 39423
rect 8159 39389 8171 39423
rect 8113 39383 8171 39389
rect 8128 39352 8156 39383
rect 7668 39324 8156 39352
rect 2961 39287 3019 39293
rect 2961 39253 2973 39287
rect 3007 39284 3019 39287
rect 5994 39284 6000 39296
rect 3007 39256 6000 39284
rect 3007 39253 3019 39256
rect 2961 39247 3019 39253
rect 5994 39244 6000 39256
rect 6052 39244 6058 39296
rect 7668 39293 7696 39324
rect 7653 39287 7711 39293
rect 7653 39253 7665 39287
rect 7699 39253 7711 39287
rect 7653 39247 7711 39253
rect 7926 39244 7932 39296
rect 7984 39244 7990 39296
rect 8294 39244 8300 39296
rect 8352 39244 8358 39296
rect 1104 39194 8740 39216
rect 1104 39142 3010 39194
rect 3062 39142 3074 39194
rect 3126 39142 3138 39194
rect 3190 39142 3202 39194
rect 3254 39142 3266 39194
rect 3318 39142 8740 39194
rect 1104 39120 8740 39142
rect 7742 38904 7748 38956
rect 7800 38904 7806 38956
rect 7834 38904 7840 38956
rect 7892 38944 7898 38956
rect 8113 38947 8171 38953
rect 8113 38944 8125 38947
rect 7892 38916 8125 38944
rect 7892 38904 7898 38916
rect 8113 38913 8125 38916
rect 8159 38913 8171 38947
rect 8113 38907 8171 38913
rect 7926 38768 7932 38820
rect 7984 38768 7990 38820
rect 8294 38700 8300 38752
rect 8352 38700 8358 38752
rect 1104 38650 8740 38672
rect 1104 38598 1950 38650
rect 2002 38598 2014 38650
rect 2066 38598 2078 38650
rect 2130 38598 2142 38650
rect 2194 38598 2206 38650
rect 2258 38598 7950 38650
rect 8002 38598 8014 38650
rect 8066 38598 8078 38650
rect 8130 38598 8142 38650
rect 8194 38598 8206 38650
rect 8258 38598 8740 38650
rect 1104 38576 8740 38598
rect 7653 38539 7711 38545
rect 7653 38505 7665 38539
rect 7699 38536 7711 38539
rect 7742 38536 7748 38548
rect 7699 38508 7748 38536
rect 7699 38505 7711 38508
rect 7653 38499 7711 38505
rect 7742 38496 7748 38508
rect 7800 38496 7806 38548
rect 5718 38360 5724 38412
rect 5776 38400 5782 38412
rect 5776 38372 8156 38400
rect 5776 38360 5782 38372
rect 1302 38292 1308 38344
rect 1360 38332 1366 38344
rect 2685 38335 2743 38341
rect 2685 38332 2697 38335
rect 1360 38304 2697 38332
rect 1360 38292 1366 38304
rect 2685 38301 2697 38304
rect 2731 38301 2743 38335
rect 2685 38295 2743 38301
rect 5534 38292 5540 38344
rect 5592 38332 5598 38344
rect 7469 38335 7527 38341
rect 7469 38332 7481 38335
rect 5592 38304 7481 38332
rect 5592 38292 5598 38304
rect 7469 38301 7481 38304
rect 7515 38301 7527 38335
rect 7469 38295 7527 38301
rect 7742 38292 7748 38344
rect 7800 38292 7806 38344
rect 8128 38341 8156 38372
rect 8113 38335 8171 38341
rect 8113 38301 8125 38335
rect 8159 38301 8171 38335
rect 8113 38295 8171 38301
rect 2869 38199 2927 38205
rect 2869 38165 2881 38199
rect 2915 38196 2927 38199
rect 6822 38196 6828 38208
rect 2915 38168 6828 38196
rect 2915 38165 2927 38168
rect 2869 38159 2927 38165
rect 6822 38156 6828 38168
rect 6880 38156 6886 38208
rect 7926 38156 7932 38208
rect 7984 38156 7990 38208
rect 8294 38156 8300 38208
rect 8352 38156 8358 38208
rect 1104 38106 8740 38128
rect 1104 38054 3010 38106
rect 3062 38054 3074 38106
rect 3126 38054 3138 38106
rect 3190 38054 3202 38106
rect 3254 38054 3266 38106
rect 3318 38054 8740 38106
rect 1104 38032 8740 38054
rect 7653 37995 7711 38001
rect 7653 37961 7665 37995
rect 7699 37992 7711 37995
rect 7834 37992 7840 38004
rect 7699 37964 7840 37992
rect 7699 37961 7711 37964
rect 7653 37955 7711 37961
rect 7834 37952 7840 37964
rect 7892 37952 7898 38004
rect 5994 37884 6000 37936
rect 6052 37924 6058 37936
rect 6052 37896 8156 37924
rect 6052 37884 6058 37896
rect 7466 37816 7472 37868
rect 7524 37816 7530 37868
rect 7650 37816 7656 37868
rect 7708 37856 7714 37868
rect 8128 37865 8156 37896
rect 7745 37859 7803 37865
rect 7745 37856 7757 37859
rect 7708 37828 7757 37856
rect 7708 37816 7714 37828
rect 7745 37825 7757 37828
rect 7791 37825 7803 37859
rect 7745 37819 7803 37825
rect 8113 37859 8171 37865
rect 8113 37825 8125 37859
rect 8159 37825 8171 37859
rect 8113 37819 8171 37825
rect 7926 37680 7932 37732
rect 7984 37680 7990 37732
rect 8294 37612 8300 37664
rect 8352 37612 8358 37664
rect 1104 37562 8740 37584
rect 1104 37510 1950 37562
rect 2002 37510 2014 37562
rect 2066 37510 2078 37562
rect 2130 37510 2142 37562
rect 2194 37510 2206 37562
rect 2258 37510 7950 37562
rect 8002 37510 8014 37562
rect 8066 37510 8078 37562
rect 8130 37510 8142 37562
rect 8194 37510 8206 37562
rect 8258 37510 8740 37562
rect 1104 37488 8740 37510
rect 7653 37451 7711 37457
rect 7653 37417 7665 37451
rect 7699 37448 7711 37451
rect 7742 37448 7748 37460
rect 7699 37420 7748 37448
rect 7699 37417 7711 37420
rect 7653 37411 7711 37417
rect 7742 37408 7748 37420
rect 7800 37408 7806 37460
rect 6914 37204 6920 37256
rect 6972 37244 6978 37256
rect 7469 37247 7527 37253
rect 7469 37244 7481 37247
rect 6972 37216 7481 37244
rect 6972 37204 6978 37216
rect 7469 37213 7481 37216
rect 7515 37213 7527 37247
rect 7469 37207 7527 37213
rect 7745 37247 7803 37253
rect 7745 37213 7757 37247
rect 7791 37213 7803 37247
rect 8113 37247 8171 37253
rect 8113 37244 8125 37247
rect 7745 37207 7803 37213
rect 7852 37216 8125 37244
rect 6822 37136 6828 37188
rect 6880 37176 6886 37188
rect 7760 37176 7788 37207
rect 6880 37148 7788 37176
rect 6880 37136 6886 37148
rect 5718 37068 5724 37120
rect 5776 37108 5782 37120
rect 7852 37108 7880 37216
rect 8113 37213 8125 37216
rect 8159 37213 8171 37247
rect 8113 37207 8171 37213
rect 5776 37080 7880 37108
rect 5776 37068 5782 37080
rect 7926 37068 7932 37120
rect 7984 37068 7990 37120
rect 8294 37068 8300 37120
rect 8352 37068 8358 37120
rect 1104 37018 8740 37040
rect 1104 36966 3010 37018
rect 3062 36966 3074 37018
rect 3126 36966 3138 37018
rect 3190 36966 3202 37018
rect 3254 36966 3266 37018
rect 3318 36966 8740 37018
rect 1104 36944 8740 36966
rect 2593 36907 2651 36913
rect 2593 36873 2605 36907
rect 2639 36904 2651 36907
rect 2639 36876 2774 36904
rect 2639 36873 2651 36876
rect 2593 36867 2651 36873
rect 2406 36728 2412 36780
rect 2464 36728 2470 36780
rect 2746 36768 2774 36876
rect 7745 36771 7803 36777
rect 7745 36768 7757 36771
rect 2746 36740 7757 36768
rect 7745 36737 7757 36740
rect 7791 36737 7803 36771
rect 7745 36731 7803 36737
rect 8113 36771 8171 36777
rect 8113 36737 8125 36771
rect 8159 36737 8171 36771
rect 8113 36731 8171 36737
rect 3970 36660 3976 36712
rect 4028 36700 4034 36712
rect 8128 36700 8156 36731
rect 4028 36672 8156 36700
rect 4028 36660 4034 36672
rect 7926 36592 7932 36644
rect 7984 36592 7990 36644
rect 8294 36524 8300 36576
rect 8352 36524 8358 36576
rect 1104 36474 8740 36496
rect 1104 36422 1950 36474
rect 2002 36422 2014 36474
rect 2066 36422 2078 36474
rect 2130 36422 2142 36474
rect 2194 36422 2206 36474
rect 2258 36422 7950 36474
rect 8002 36422 8014 36474
rect 8066 36422 8078 36474
rect 8130 36422 8142 36474
rect 8194 36422 8206 36474
rect 8258 36422 8740 36474
rect 1104 36400 8740 36422
rect 2225 36295 2283 36301
rect 2225 36261 2237 36295
rect 2271 36292 2283 36295
rect 2271 36264 2774 36292
rect 2271 36261 2283 36264
rect 2225 36255 2283 36261
rect 842 36116 848 36168
rect 900 36156 906 36168
rect 2041 36159 2099 36165
rect 2041 36156 2053 36159
rect 900 36128 2053 36156
rect 900 36116 906 36128
rect 2041 36125 2053 36128
rect 2087 36125 2099 36159
rect 2746 36156 2774 36264
rect 7745 36159 7803 36165
rect 7745 36156 7757 36159
rect 2746 36128 7757 36156
rect 2041 36119 2099 36125
rect 7745 36125 7757 36128
rect 7791 36125 7803 36159
rect 7745 36119 7803 36125
rect 8113 36159 8171 36165
rect 8113 36125 8125 36159
rect 8159 36125 8171 36159
rect 8113 36119 8171 36125
rect 5350 36048 5356 36100
rect 5408 36088 5414 36100
rect 8128 36088 8156 36119
rect 5408 36060 8156 36088
rect 5408 36048 5414 36060
rect 7926 35980 7932 36032
rect 7984 35980 7990 36032
rect 8294 35980 8300 36032
rect 8352 35980 8358 36032
rect 1104 35930 8740 35952
rect 1104 35878 3010 35930
rect 3062 35878 3074 35930
rect 3126 35878 3138 35930
rect 3190 35878 3202 35930
rect 3254 35878 3266 35930
rect 3318 35878 8740 35930
rect 1104 35856 8740 35878
rect 4338 35640 4344 35692
rect 4396 35680 4402 35692
rect 7745 35683 7803 35689
rect 7745 35680 7757 35683
rect 4396 35652 7757 35680
rect 4396 35640 4402 35652
rect 7745 35649 7757 35652
rect 7791 35649 7803 35683
rect 7745 35643 7803 35649
rect 8113 35683 8171 35689
rect 8113 35649 8125 35683
rect 8159 35649 8171 35683
rect 8113 35643 8171 35649
rect 6178 35572 6184 35624
rect 6236 35612 6242 35624
rect 8128 35612 8156 35643
rect 6236 35584 8156 35612
rect 6236 35572 6242 35584
rect 7926 35504 7932 35556
rect 7984 35504 7990 35556
rect 8294 35436 8300 35488
rect 8352 35436 8358 35488
rect 1104 35386 8740 35408
rect 1104 35334 1950 35386
rect 2002 35334 2014 35386
rect 2066 35334 2078 35386
rect 2130 35334 2142 35386
rect 2194 35334 2206 35386
rect 2258 35334 7950 35386
rect 8002 35334 8014 35386
rect 8066 35334 8078 35386
rect 8130 35334 8142 35386
rect 8194 35334 8206 35386
rect 8258 35334 8740 35386
rect 1104 35312 8740 35334
rect 1765 35275 1823 35281
rect 1765 35241 1777 35275
rect 1811 35272 1823 35275
rect 5350 35272 5356 35284
rect 1811 35244 5356 35272
rect 1811 35241 1823 35244
rect 1765 35235 1823 35241
rect 5350 35232 5356 35244
rect 5408 35232 5414 35284
rect 7650 35232 7656 35284
rect 7708 35232 7714 35284
rect 3878 35096 3884 35148
rect 3936 35136 3942 35148
rect 3936 35108 8156 35136
rect 3936 35096 3942 35108
rect 290 35028 296 35080
rect 348 35068 354 35080
rect 1581 35071 1639 35077
rect 1581 35068 1593 35071
rect 348 35040 1593 35068
rect 348 35028 354 35040
rect 1581 35037 1593 35040
rect 1627 35037 1639 35071
rect 1581 35031 1639 35037
rect 7466 35028 7472 35080
rect 7524 35028 7530 35080
rect 8128 35077 8156 35108
rect 7745 35071 7803 35077
rect 7745 35037 7757 35071
rect 7791 35037 7803 35071
rect 7745 35031 7803 35037
rect 8113 35071 8171 35077
rect 8113 35037 8125 35071
rect 8159 35037 8171 35071
rect 8113 35031 8171 35037
rect 3694 34960 3700 35012
rect 3752 35000 3758 35012
rect 7760 35000 7788 35031
rect 3752 34972 7788 35000
rect 3752 34960 3758 34972
rect 7926 34892 7932 34944
rect 7984 34892 7990 34944
rect 8294 34892 8300 34944
rect 8352 34892 8358 34944
rect 1104 34842 8740 34864
rect 1104 34790 3010 34842
rect 3062 34790 3074 34842
rect 3126 34790 3138 34842
rect 3190 34790 3202 34842
rect 3254 34790 3266 34842
rect 3318 34790 8740 34842
rect 1104 34768 8740 34790
rect 7929 34731 7987 34737
rect 7929 34697 7941 34731
rect 7975 34728 7987 34731
rect 8846 34728 8852 34740
rect 7975 34700 8852 34728
rect 7975 34697 7987 34700
rect 7929 34691 7987 34697
rect 8846 34688 8852 34700
rect 8904 34688 8910 34740
rect 1762 34552 1768 34604
rect 1820 34592 1826 34604
rect 7745 34595 7803 34601
rect 7745 34592 7757 34595
rect 1820 34564 7757 34592
rect 1820 34552 1826 34564
rect 7745 34561 7757 34564
rect 7791 34561 7803 34595
rect 7745 34555 7803 34561
rect 8113 34595 8171 34601
rect 8113 34561 8125 34595
rect 8159 34561 8171 34595
rect 8113 34555 8171 34561
rect 2314 34484 2320 34536
rect 2372 34524 2378 34536
rect 8128 34524 8156 34555
rect 2372 34496 8156 34524
rect 2372 34484 2378 34496
rect 8294 34348 8300 34400
rect 8352 34348 8358 34400
rect 1104 34298 8740 34320
rect 1104 34246 1950 34298
rect 2002 34246 2014 34298
rect 2066 34246 2078 34298
rect 2130 34246 2142 34298
rect 2194 34246 2206 34298
rect 2258 34246 7950 34298
rect 8002 34246 8014 34298
rect 8066 34246 8078 34298
rect 8130 34246 8142 34298
rect 8194 34246 8206 34298
rect 8258 34246 8740 34298
rect 1104 34224 8740 34246
rect 658 33940 664 33992
rect 716 33980 722 33992
rect 2041 33983 2099 33989
rect 2041 33980 2053 33983
rect 716 33952 2053 33980
rect 716 33940 722 33952
rect 2041 33949 2053 33952
rect 2087 33949 2099 33983
rect 2041 33943 2099 33949
rect 6362 33940 6368 33992
rect 6420 33980 6426 33992
rect 7745 33983 7803 33989
rect 7745 33980 7757 33983
rect 6420 33952 7757 33980
rect 6420 33940 6426 33952
rect 7745 33949 7757 33952
rect 7791 33949 7803 33983
rect 7745 33943 7803 33949
rect 8110 33940 8116 33992
rect 8168 33940 8174 33992
rect 2225 33847 2283 33853
rect 2225 33813 2237 33847
rect 2271 33844 2283 33847
rect 7742 33844 7748 33856
rect 2271 33816 7748 33844
rect 2271 33813 2283 33816
rect 2225 33807 2283 33813
rect 7742 33804 7748 33816
rect 7800 33804 7806 33856
rect 7926 33804 7932 33856
rect 7984 33804 7990 33856
rect 8294 33804 8300 33856
rect 8352 33804 8358 33856
rect 1104 33754 8740 33776
rect 1104 33702 3010 33754
rect 3062 33702 3074 33754
rect 3126 33702 3138 33754
rect 3190 33702 3202 33754
rect 3254 33702 3266 33754
rect 3318 33702 8740 33754
rect 1104 33680 8740 33702
rect 1857 33643 1915 33649
rect 1857 33609 1869 33643
rect 1903 33640 1915 33643
rect 4338 33640 4344 33652
rect 1903 33612 4344 33640
rect 1903 33609 1915 33612
rect 1857 33603 1915 33609
rect 4338 33600 4344 33612
rect 4396 33600 4402 33652
rect 1486 33464 1492 33516
rect 1544 33504 1550 33516
rect 1673 33507 1731 33513
rect 1673 33504 1685 33507
rect 1544 33476 1685 33504
rect 1544 33464 1550 33476
rect 1673 33473 1685 33476
rect 1719 33473 1731 33507
rect 1673 33467 1731 33473
rect 7742 33464 7748 33516
rect 7800 33464 7806 33516
rect 7834 33464 7840 33516
rect 7892 33504 7898 33516
rect 8113 33507 8171 33513
rect 8113 33504 8125 33507
rect 7892 33476 8125 33504
rect 7892 33464 7898 33476
rect 8113 33473 8125 33476
rect 8159 33473 8171 33507
rect 8113 33467 8171 33473
rect 7926 33328 7932 33380
rect 7984 33328 7990 33380
rect 8294 33260 8300 33312
rect 8352 33260 8358 33312
rect 1104 33210 8740 33232
rect 1104 33158 1950 33210
rect 2002 33158 2014 33210
rect 2066 33158 2078 33210
rect 2130 33158 2142 33210
rect 2194 33158 2206 33210
rect 2258 33158 7950 33210
rect 8002 33158 8014 33210
rect 8066 33158 8078 33210
rect 8130 33158 8142 33210
rect 8194 33158 8206 33210
rect 8258 33158 8740 33210
rect 1104 33136 8740 33158
rect 2593 33099 2651 33105
rect 2593 33065 2605 33099
rect 2639 33096 2651 33099
rect 7834 33096 7840 33108
rect 2639 33068 7840 33096
rect 2639 33065 2651 33068
rect 2593 33059 2651 33065
rect 7834 33056 7840 33068
rect 7892 33056 7898 33108
rect 566 32852 572 32904
rect 624 32892 630 32904
rect 2409 32895 2467 32901
rect 2409 32892 2421 32895
rect 624 32864 2421 32892
rect 624 32852 630 32864
rect 2409 32861 2421 32864
rect 2455 32861 2467 32895
rect 2409 32855 2467 32861
rect 6270 32852 6276 32904
rect 6328 32892 6334 32904
rect 7469 32895 7527 32901
rect 7469 32892 7481 32895
rect 6328 32864 7481 32892
rect 6328 32852 6334 32864
rect 7469 32861 7481 32864
rect 7515 32861 7527 32895
rect 7469 32855 7527 32861
rect 7742 32852 7748 32904
rect 7800 32852 7806 32904
rect 8113 32895 8171 32901
rect 8113 32861 8125 32895
rect 8159 32861 8171 32895
rect 8113 32855 8171 32861
rect 3510 32784 3516 32836
rect 3568 32824 3574 32836
rect 8128 32824 8156 32855
rect 3568 32796 8156 32824
rect 3568 32784 3574 32796
rect 7653 32759 7711 32765
rect 7653 32725 7665 32759
rect 7699 32756 7711 32759
rect 7834 32756 7840 32768
rect 7699 32728 7840 32756
rect 7699 32725 7711 32728
rect 7653 32719 7711 32725
rect 7834 32716 7840 32728
rect 7892 32716 7898 32768
rect 7926 32716 7932 32768
rect 7984 32716 7990 32768
rect 8294 32716 8300 32768
rect 8352 32716 8358 32768
rect 1104 32666 8740 32688
rect 1104 32614 3010 32666
rect 3062 32614 3074 32666
rect 3126 32614 3138 32666
rect 3190 32614 3202 32666
rect 3254 32614 3266 32666
rect 3318 32614 8740 32666
rect 1104 32592 8740 32614
rect 2777 32555 2835 32561
rect 2777 32521 2789 32555
rect 2823 32552 2835 32555
rect 7742 32552 7748 32564
rect 2823 32524 7748 32552
rect 2823 32521 2835 32524
rect 2777 32515 2835 32521
rect 7742 32512 7748 32524
rect 7800 32512 7806 32564
rect 474 32376 480 32428
rect 532 32416 538 32428
rect 2593 32419 2651 32425
rect 2593 32416 2605 32419
rect 532 32388 2605 32416
rect 532 32376 538 32388
rect 2593 32385 2605 32388
rect 2639 32385 2651 32419
rect 2593 32379 2651 32385
rect 7742 32376 7748 32428
rect 7800 32376 7806 32428
rect 8113 32419 8171 32425
rect 8113 32385 8125 32419
rect 8159 32385 8171 32419
rect 8113 32379 8171 32385
rect 7190 32308 7196 32360
rect 7248 32348 7254 32360
rect 8128 32348 8156 32379
rect 7248 32320 8156 32348
rect 7248 32308 7254 32320
rect 7926 32240 7932 32292
rect 7984 32240 7990 32292
rect 8294 32172 8300 32224
rect 8352 32172 8358 32224
rect 1104 32122 8740 32144
rect 1104 32070 1950 32122
rect 2002 32070 2014 32122
rect 2066 32070 2078 32122
rect 2130 32070 2142 32122
rect 2194 32070 2206 32122
rect 2258 32070 7950 32122
rect 8002 32070 8014 32122
rect 8066 32070 8078 32122
rect 8130 32070 8142 32122
rect 8194 32070 8206 32122
rect 8258 32070 8740 32122
rect 1104 32048 8740 32070
rect 2961 32011 3019 32017
rect 2961 31977 2973 32011
rect 3007 32008 3019 32011
rect 3510 32008 3516 32020
rect 3007 31980 3516 32008
rect 3007 31977 3019 31980
rect 2961 31971 3019 31977
rect 3510 31968 3516 31980
rect 3568 31968 3574 32020
rect 7929 31943 7987 31949
rect 7929 31909 7941 31943
rect 7975 31940 7987 31943
rect 8846 31940 8852 31952
rect 7975 31912 8852 31940
rect 7975 31909 7987 31912
rect 7929 31903 7987 31909
rect 8846 31900 8852 31912
rect 8904 31900 8910 31952
rect 3510 31832 3516 31884
rect 3568 31872 3574 31884
rect 3694 31872 3700 31884
rect 3568 31844 3700 31872
rect 3568 31832 3574 31844
rect 3694 31832 3700 31844
rect 3752 31832 3758 31884
rect 2774 31764 2780 31816
rect 2832 31764 2838 31816
rect 4062 31764 4068 31816
rect 4120 31804 4126 31816
rect 7193 31807 7251 31813
rect 7193 31804 7205 31807
rect 4120 31776 7205 31804
rect 4120 31764 4126 31776
rect 7193 31773 7205 31776
rect 7239 31773 7251 31807
rect 7193 31767 7251 31773
rect 7466 31764 7472 31816
rect 7524 31804 7530 31816
rect 7745 31807 7803 31813
rect 7745 31804 7757 31807
rect 7524 31776 7757 31804
rect 7524 31764 7530 31776
rect 7745 31773 7757 31776
rect 7791 31773 7803 31807
rect 7745 31767 7803 31773
rect 7834 31764 7840 31816
rect 7892 31804 7898 31816
rect 8113 31807 8171 31813
rect 8113 31804 8125 31807
rect 7892 31776 8125 31804
rect 7892 31764 7898 31776
rect 8113 31773 8125 31776
rect 8159 31773 8171 31807
rect 8113 31767 8171 31773
rect 7374 31628 7380 31680
rect 7432 31628 7438 31680
rect 8294 31628 8300 31680
rect 8352 31628 8358 31680
rect 1104 31578 8740 31600
rect 1104 31526 3010 31578
rect 3062 31526 3074 31578
rect 3126 31526 3138 31578
rect 3190 31526 3202 31578
rect 3254 31526 3266 31578
rect 3318 31526 8740 31578
rect 1104 31504 8740 31526
rect 2225 31467 2283 31473
rect 2225 31433 2237 31467
rect 2271 31464 2283 31467
rect 7742 31464 7748 31476
rect 2271 31436 7748 31464
rect 2271 31433 2283 31436
rect 2225 31427 2283 31433
rect 7742 31424 7748 31436
rect 7800 31424 7806 31476
rect 198 31288 204 31340
rect 256 31328 262 31340
rect 2041 31331 2099 31337
rect 2041 31328 2053 31331
rect 256 31300 2053 31328
rect 256 31288 262 31300
rect 2041 31297 2053 31300
rect 2087 31297 2099 31331
rect 2041 31291 2099 31297
rect 7650 31288 7656 31340
rect 7708 31328 7714 31340
rect 7745 31331 7803 31337
rect 7745 31328 7757 31331
rect 7708 31300 7757 31328
rect 7708 31288 7714 31300
rect 7745 31297 7757 31300
rect 7791 31297 7803 31331
rect 7745 31291 7803 31297
rect 8113 31331 8171 31337
rect 8113 31297 8125 31331
rect 8159 31297 8171 31331
rect 8113 31291 8171 31297
rect 6638 31220 6644 31272
rect 6696 31260 6702 31272
rect 8128 31260 8156 31291
rect 6696 31232 8156 31260
rect 6696 31220 6702 31232
rect 7926 31152 7932 31204
rect 7984 31152 7990 31204
rect 2774 31084 2780 31136
rect 2832 31084 2838 31136
rect 8294 31084 8300 31136
rect 8352 31084 8358 31136
rect 1104 31034 8740 31056
rect 1104 30982 1950 31034
rect 2002 30982 2014 31034
rect 2066 30982 2078 31034
rect 2130 30982 2142 31034
rect 2194 30982 2206 31034
rect 2258 30982 7950 31034
rect 8002 30982 8014 31034
rect 8066 30982 8078 31034
rect 8130 30982 8142 31034
rect 8194 30982 8206 31034
rect 8258 30982 8740 31034
rect 1104 30960 8740 30982
rect 7006 30812 7012 30864
rect 7064 30852 7070 30864
rect 7064 30824 8156 30852
rect 7064 30812 7070 30824
rect 5166 30676 5172 30728
rect 5224 30716 5230 30728
rect 8128 30725 8156 30824
rect 7009 30719 7067 30725
rect 7009 30716 7021 30719
rect 5224 30688 7021 30716
rect 5224 30676 5230 30688
rect 7009 30685 7021 30688
rect 7055 30685 7067 30719
rect 7009 30679 7067 30685
rect 7745 30719 7803 30725
rect 7745 30685 7757 30719
rect 7791 30685 7803 30719
rect 7745 30679 7803 30685
rect 8113 30719 8171 30725
rect 8113 30685 8125 30719
rect 8159 30685 8171 30719
rect 8113 30679 8171 30685
rect 5350 30608 5356 30660
rect 5408 30648 5414 30660
rect 7760 30648 7788 30679
rect 5408 30620 7788 30648
rect 5408 30608 5414 30620
rect 7193 30583 7251 30589
rect 7193 30549 7205 30583
rect 7239 30580 7251 30583
rect 7834 30580 7840 30592
rect 7239 30552 7840 30580
rect 7239 30549 7251 30552
rect 7193 30543 7251 30549
rect 7834 30540 7840 30552
rect 7892 30540 7898 30592
rect 7926 30540 7932 30592
rect 7984 30540 7990 30592
rect 8294 30540 8300 30592
rect 8352 30540 8358 30592
rect 1104 30490 8740 30512
rect 1104 30438 3010 30490
rect 3062 30438 3074 30490
rect 3126 30438 3138 30490
rect 3190 30438 3202 30490
rect 3254 30438 3266 30490
rect 3318 30438 8740 30490
rect 1104 30416 8740 30438
rect 106 30200 112 30252
rect 164 30240 170 30252
rect 1581 30243 1639 30249
rect 1581 30240 1593 30243
rect 164 30212 1593 30240
rect 164 30200 170 30212
rect 1581 30209 1593 30212
rect 1627 30209 1639 30243
rect 1581 30203 1639 30209
rect 2593 30243 2651 30249
rect 2593 30209 2605 30243
rect 2639 30209 2651 30243
rect 2593 30203 2651 30209
rect 7101 30243 7159 30249
rect 7101 30209 7113 30243
rect 7147 30209 7159 30243
rect 7101 30203 7159 30209
rect 382 30132 388 30184
rect 440 30172 446 30184
rect 2608 30172 2636 30203
rect 440 30144 2636 30172
rect 7116 30172 7144 30203
rect 7374 30200 7380 30252
rect 7432 30240 7438 30252
rect 7745 30243 7803 30249
rect 7745 30240 7757 30243
rect 7432 30212 7757 30240
rect 7432 30200 7438 30212
rect 7745 30209 7757 30212
rect 7791 30209 7803 30243
rect 7745 30203 7803 30209
rect 7834 30200 7840 30252
rect 7892 30240 7898 30252
rect 8113 30243 8171 30249
rect 8113 30240 8125 30243
rect 7892 30212 8125 30240
rect 7892 30200 7898 30212
rect 8113 30209 8125 30212
rect 8159 30209 8171 30243
rect 8113 30203 8171 30209
rect 9122 30172 9128 30184
rect 7116 30144 9128 30172
rect 440 30132 446 30144
rect 9122 30132 9128 30144
rect 9180 30132 9186 30184
rect 1765 30107 1823 30113
rect 1765 30073 1777 30107
rect 1811 30104 1823 30107
rect 7466 30104 7472 30116
rect 1811 30076 7472 30104
rect 1811 30073 1823 30076
rect 1765 30067 1823 30073
rect 7466 30064 7472 30076
rect 7524 30064 7530 30116
rect 7926 30064 7932 30116
rect 7984 30064 7990 30116
rect 2777 30039 2835 30045
rect 2777 30005 2789 30039
rect 2823 30036 2835 30039
rect 7190 30036 7196 30048
rect 2823 30008 7196 30036
rect 2823 30005 2835 30008
rect 2777 29999 2835 30005
rect 7190 29996 7196 30008
rect 7248 29996 7254 30048
rect 7285 30039 7343 30045
rect 7285 30005 7297 30039
rect 7331 30036 7343 30039
rect 7742 30036 7748 30048
rect 7331 30008 7748 30036
rect 7331 30005 7343 30008
rect 7285 29999 7343 30005
rect 7742 29996 7748 30008
rect 7800 29996 7806 30048
rect 8294 29996 8300 30048
rect 8352 29996 8358 30048
rect 1104 29946 8740 29968
rect 1104 29894 1950 29946
rect 2002 29894 2014 29946
rect 2066 29894 2078 29946
rect 2130 29894 2142 29946
rect 2194 29894 2206 29946
rect 2258 29894 7950 29946
rect 8002 29894 8014 29946
rect 8066 29894 8078 29946
rect 8130 29894 8142 29946
rect 8194 29894 8206 29946
rect 8258 29894 8740 29946
rect 1104 29872 8740 29894
rect 9214 29696 9220 29708
rect 7300 29668 9220 29696
rect 7300 29637 7328 29668
rect 9214 29656 9220 29668
rect 9272 29656 9278 29708
rect 7285 29631 7343 29637
rect 7285 29597 7297 29631
rect 7331 29597 7343 29631
rect 7285 29591 7343 29597
rect 7742 29588 7748 29640
rect 7800 29588 7806 29640
rect 8113 29631 8171 29637
rect 8113 29597 8125 29631
rect 8159 29597 8171 29631
rect 8113 29591 8171 29597
rect 8128 29560 8156 29591
rect 7484 29532 8156 29560
rect 7484 29501 7512 29532
rect 7469 29495 7527 29501
rect 7469 29461 7481 29495
rect 7515 29461 7527 29495
rect 7469 29455 7527 29461
rect 7926 29452 7932 29504
rect 7984 29452 7990 29504
rect 8294 29452 8300 29504
rect 8352 29452 8358 29504
rect 1104 29402 8740 29424
rect 1104 29350 3010 29402
rect 3062 29350 3074 29402
rect 3126 29350 3138 29402
rect 3190 29350 3202 29402
rect 3254 29350 3266 29402
rect 3318 29350 8740 29402
rect 1104 29328 8740 29350
rect 2685 29291 2743 29297
rect 2685 29257 2697 29291
rect 2731 29288 2743 29291
rect 5718 29288 5724 29300
rect 2731 29260 5724 29288
rect 2731 29257 2743 29260
rect 2685 29251 2743 29257
rect 5718 29248 5724 29260
rect 5776 29248 5782 29300
rect 7285 29291 7343 29297
rect 7285 29257 7297 29291
rect 7331 29257 7343 29291
rect 7285 29251 7343 29257
rect 1302 29112 1308 29164
rect 1360 29152 1366 29164
rect 2501 29155 2559 29161
rect 2501 29152 2513 29155
rect 1360 29124 2513 29152
rect 1360 29112 1366 29124
rect 2501 29121 2513 29124
rect 2547 29121 2559 29155
rect 2501 29115 2559 29121
rect 7101 29155 7159 29161
rect 7101 29121 7113 29155
rect 7147 29121 7159 29155
rect 7300 29152 7328 29251
rect 7745 29155 7803 29161
rect 7745 29152 7757 29155
rect 7300 29124 7757 29152
rect 7101 29115 7159 29121
rect 7745 29121 7757 29124
rect 7791 29121 7803 29155
rect 7745 29115 7803 29121
rect 7116 29084 7144 29115
rect 7834 29112 7840 29164
rect 7892 29152 7898 29164
rect 8113 29155 8171 29161
rect 8113 29152 8125 29155
rect 7892 29124 8125 29152
rect 7892 29112 7898 29124
rect 8113 29121 8125 29124
rect 8159 29121 8171 29155
rect 8113 29115 8171 29121
rect 9490 29084 9496 29096
rect 7116 29056 9496 29084
rect 9490 29044 9496 29056
rect 9548 29044 9554 29096
rect 4798 28976 4804 29028
rect 4856 29016 4862 29028
rect 5902 29016 5908 29028
rect 4856 28988 5908 29016
rect 4856 28976 4862 28988
rect 5902 28976 5908 28988
rect 5960 28976 5966 29028
rect 7929 29019 7987 29025
rect 7929 28985 7941 29019
rect 7975 29016 7987 29019
rect 8938 29016 8944 29028
rect 7975 28988 8944 29016
rect 7975 28985 7987 28988
rect 7929 28979 7987 28985
rect 8938 28976 8944 28988
rect 8996 28976 9002 29028
rect 8294 28908 8300 28960
rect 8352 28908 8358 28960
rect 1104 28858 8740 28880
rect 1104 28806 1950 28858
rect 2002 28806 2014 28858
rect 2066 28806 2078 28858
rect 2130 28806 2142 28858
rect 2194 28806 2206 28858
rect 2258 28806 7950 28858
rect 8002 28806 8014 28858
rect 8066 28806 8078 28858
rect 8130 28806 8142 28858
rect 8194 28806 8206 28858
rect 8258 28806 8740 28858
rect 1104 28784 8740 28806
rect 7653 28747 7711 28753
rect 7653 28713 7665 28747
rect 7699 28744 7711 28747
rect 7834 28744 7840 28756
rect 7699 28716 7840 28744
rect 7699 28713 7711 28716
rect 7653 28707 7711 28713
rect 7834 28704 7840 28716
rect 7892 28704 7898 28756
rect 8662 28608 8668 28620
rect 7484 28580 8668 28608
rect 7484 28549 7512 28580
rect 8662 28568 8668 28580
rect 8720 28568 8726 28620
rect 7469 28543 7527 28549
rect 7469 28509 7481 28543
rect 7515 28509 7527 28543
rect 7469 28503 7527 28509
rect 7745 28543 7803 28549
rect 7745 28509 7757 28543
rect 7791 28509 7803 28543
rect 7745 28503 7803 28509
rect 7282 28432 7288 28484
rect 7340 28472 7346 28484
rect 7760 28472 7788 28503
rect 8110 28500 8116 28552
rect 8168 28500 8174 28552
rect 7340 28444 7788 28472
rect 7340 28432 7346 28444
rect 7926 28364 7932 28416
rect 7984 28364 7990 28416
rect 8294 28364 8300 28416
rect 8352 28364 8358 28416
rect 1104 28314 8740 28336
rect 1104 28262 3010 28314
rect 3062 28262 3074 28314
rect 3126 28262 3138 28314
rect 3190 28262 3202 28314
rect 3254 28262 3266 28314
rect 3318 28262 8740 28314
rect 1104 28240 8740 28262
rect 7653 28203 7711 28209
rect 7653 28169 7665 28203
rect 7699 28200 7711 28203
rect 8110 28200 8116 28212
rect 7699 28172 8116 28200
rect 7699 28169 7711 28172
rect 7653 28163 7711 28169
rect 8110 28160 8116 28172
rect 8168 28160 8174 28212
rect 7469 28067 7527 28073
rect 7469 28033 7481 28067
rect 7515 28033 7527 28067
rect 7469 28027 7527 28033
rect 7484 27996 7512 28027
rect 7742 28024 7748 28076
rect 7800 28024 7806 28076
rect 7834 28024 7840 28076
rect 7892 28064 7898 28076
rect 8113 28067 8171 28073
rect 8113 28064 8125 28067
rect 7892 28036 8125 28064
rect 7892 28024 7898 28036
rect 8113 28033 8125 28036
rect 8159 28033 8171 28067
rect 8113 28027 8171 28033
rect 8938 27996 8944 28008
rect 7484 27968 8944 27996
rect 8938 27956 8944 27968
rect 8996 27956 9002 28008
rect 7926 27888 7932 27940
rect 7984 27888 7990 27940
rect 8294 27820 8300 27872
rect 8352 27820 8358 27872
rect 1104 27770 8740 27792
rect 1104 27718 1950 27770
rect 2002 27718 2014 27770
rect 2066 27718 2078 27770
rect 2130 27718 2142 27770
rect 2194 27718 2206 27770
rect 2258 27718 7950 27770
rect 8002 27718 8014 27770
rect 8066 27718 8078 27770
rect 8130 27718 8142 27770
rect 8194 27718 8206 27770
rect 8258 27718 8740 27770
rect 1104 27696 8740 27718
rect 7653 27659 7711 27665
rect 7653 27625 7665 27659
rect 7699 27656 7711 27659
rect 7742 27656 7748 27668
rect 7699 27628 7748 27656
rect 7699 27625 7711 27628
rect 7653 27619 7711 27625
rect 7742 27616 7748 27628
rect 7800 27616 7806 27668
rect 2593 27591 2651 27597
rect 2593 27557 2605 27591
rect 2639 27588 2651 27591
rect 3970 27588 3976 27600
rect 2639 27560 3976 27588
rect 2639 27557 2651 27560
rect 2593 27551 2651 27557
rect 3970 27548 3976 27560
rect 4028 27548 4034 27600
rect 1210 27412 1216 27464
rect 1268 27452 1274 27464
rect 2409 27455 2467 27461
rect 2409 27452 2421 27455
rect 1268 27424 2421 27452
rect 1268 27412 1274 27424
rect 2409 27421 2421 27424
rect 2455 27421 2467 27455
rect 2409 27415 2467 27421
rect 6730 27412 6736 27464
rect 6788 27452 6794 27464
rect 7469 27455 7527 27461
rect 7469 27452 7481 27455
rect 6788 27424 7481 27452
rect 6788 27412 6794 27424
rect 7469 27421 7481 27424
rect 7515 27421 7527 27455
rect 7469 27415 7527 27421
rect 7558 27412 7564 27464
rect 7616 27452 7622 27464
rect 7745 27455 7803 27461
rect 7745 27452 7757 27455
rect 7616 27424 7757 27452
rect 7616 27412 7622 27424
rect 7745 27421 7757 27424
rect 7791 27421 7803 27455
rect 7745 27415 7803 27421
rect 8113 27455 8171 27461
rect 8113 27421 8125 27455
rect 8159 27421 8171 27455
rect 8113 27415 8171 27421
rect 7190 27344 7196 27396
rect 7248 27384 7254 27396
rect 8128 27384 8156 27415
rect 7248 27356 8156 27384
rect 7248 27344 7254 27356
rect 7926 27276 7932 27328
rect 7984 27276 7990 27328
rect 8294 27276 8300 27328
rect 8352 27276 8358 27328
rect 1104 27226 8740 27248
rect 1104 27174 3010 27226
rect 3062 27174 3074 27226
rect 3126 27174 3138 27226
rect 3190 27174 3202 27226
rect 3254 27174 3266 27226
rect 3318 27174 8740 27226
rect 1104 27152 8740 27174
rect 7469 27115 7527 27121
rect 7469 27081 7481 27115
rect 7515 27112 7527 27115
rect 7834 27112 7840 27124
rect 7515 27084 7840 27112
rect 7515 27081 7527 27084
rect 7469 27075 7527 27081
rect 7834 27072 7840 27084
rect 7892 27072 7898 27124
rect 7285 26979 7343 26985
rect 7285 26945 7297 26979
rect 7331 26976 7343 26979
rect 7374 26976 7380 26988
rect 7331 26948 7380 26976
rect 7331 26945 7343 26948
rect 7285 26939 7343 26945
rect 7374 26936 7380 26948
rect 7432 26936 7438 26988
rect 7742 26936 7748 26988
rect 7800 26936 7806 26988
rect 8113 26979 8171 26985
rect 8113 26945 8125 26979
rect 8159 26945 8171 26979
rect 8113 26939 8171 26945
rect 7466 26868 7472 26920
rect 7524 26908 7530 26920
rect 8128 26908 8156 26939
rect 7524 26880 8156 26908
rect 7524 26868 7530 26880
rect 7926 26800 7932 26852
rect 7984 26800 7990 26852
rect 8294 26732 8300 26784
rect 8352 26732 8358 26784
rect 1104 26682 8740 26704
rect 1104 26630 1950 26682
rect 2002 26630 2014 26682
rect 2066 26630 2078 26682
rect 2130 26630 2142 26682
rect 2194 26630 2206 26682
rect 2258 26630 7950 26682
rect 8002 26630 8014 26682
rect 8066 26630 8078 26682
rect 8130 26630 8142 26682
rect 8194 26630 8206 26682
rect 8258 26630 8740 26682
rect 1104 26608 8740 26630
rect 7193 26571 7251 26577
rect 7193 26537 7205 26571
rect 7239 26568 7251 26571
rect 7558 26568 7564 26580
rect 7239 26540 7564 26568
rect 7239 26537 7251 26540
rect 7193 26531 7251 26537
rect 7558 26528 7564 26540
rect 7616 26528 7622 26580
rect 7374 26460 7380 26512
rect 7432 26460 7438 26512
rect 7837 26503 7895 26509
rect 7837 26469 7849 26503
rect 7883 26500 7895 26503
rect 8754 26500 8760 26512
rect 7883 26472 8760 26500
rect 7883 26469 7895 26472
rect 7837 26463 7895 26469
rect 8754 26460 8760 26472
rect 8812 26460 8818 26512
rect 8570 26432 8576 26444
rect 7024 26404 8576 26432
rect 7024 26373 7052 26404
rect 8570 26392 8576 26404
rect 8628 26392 8634 26444
rect 7009 26367 7067 26373
rect 7009 26333 7021 26367
rect 7055 26333 7067 26367
rect 7009 26327 7067 26333
rect 8018 26324 8024 26376
rect 8076 26324 8082 26376
rect 8113 26367 8171 26373
rect 8113 26333 8125 26367
rect 8159 26333 8171 26367
rect 8113 26327 8171 26333
rect 2866 26256 2872 26308
rect 2924 26296 2930 26308
rect 7285 26299 7343 26305
rect 7285 26296 7297 26299
rect 2924 26268 7297 26296
rect 2924 26256 2930 26268
rect 7285 26265 7297 26268
rect 7331 26265 7343 26299
rect 7285 26259 7343 26265
rect 7374 26256 7380 26308
rect 7432 26296 7438 26308
rect 8128 26296 8156 26327
rect 7432 26268 8156 26296
rect 7432 26256 7438 26268
rect 8294 26188 8300 26240
rect 8352 26188 8358 26240
rect 1104 26138 8740 26160
rect 1104 26086 3010 26138
rect 3062 26086 3074 26138
rect 3126 26086 3138 26138
rect 3190 26086 3202 26138
rect 3254 26086 3266 26138
rect 3318 26086 8740 26138
rect 1104 26064 8740 26086
rect 2133 26027 2191 26033
rect 2133 25993 2145 26027
rect 2179 26024 2191 26027
rect 2682 26024 2688 26036
rect 2179 25996 2688 26024
rect 2179 25993 2191 25996
rect 2133 25987 2191 25993
rect 2682 25984 2688 25996
rect 2740 25984 2746 26036
rect 3145 26027 3203 26033
rect 3145 25993 3157 26027
rect 3191 26024 3203 26027
rect 5442 26024 5448 26036
rect 3191 25996 5448 26024
rect 3191 25993 3203 25996
rect 3145 25987 3203 25993
rect 5442 25984 5448 25996
rect 5500 25984 5506 26036
rect 7190 25984 7196 26036
rect 7248 25984 7254 26036
rect 8478 25956 8484 25968
rect 7024 25928 8484 25956
rect 1949 25891 2007 25897
rect 1949 25857 1961 25891
rect 1995 25888 2007 25891
rect 2498 25888 2504 25900
rect 1995 25860 2504 25888
rect 1995 25857 2007 25860
rect 1949 25851 2007 25857
rect 2498 25848 2504 25860
rect 2556 25848 2562 25900
rect 2961 25891 3019 25897
rect 2961 25857 2973 25891
rect 3007 25888 3019 25891
rect 3050 25888 3056 25900
rect 3007 25860 3056 25888
rect 3007 25857 3019 25860
rect 2961 25851 3019 25857
rect 3050 25848 3056 25860
rect 3108 25848 3114 25900
rect 7024 25897 7052 25928
rect 8478 25916 8484 25928
rect 8536 25916 8542 25968
rect 7009 25891 7067 25897
rect 7009 25857 7021 25891
rect 7055 25857 7067 25891
rect 7009 25851 7067 25857
rect 7558 25848 7564 25900
rect 7616 25888 7622 25900
rect 7745 25891 7803 25897
rect 7745 25888 7757 25891
rect 7616 25860 7757 25888
rect 7616 25848 7622 25860
rect 7745 25857 7757 25860
rect 7791 25857 7803 25891
rect 7745 25851 7803 25857
rect 8113 25891 8171 25897
rect 8113 25857 8125 25891
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 6546 25780 6552 25832
rect 6604 25820 6610 25832
rect 8128 25820 8156 25851
rect 6604 25792 8156 25820
rect 6604 25780 6610 25792
rect 7926 25712 7932 25764
rect 7984 25712 7990 25764
rect 8294 25644 8300 25696
rect 8352 25644 8358 25696
rect 1104 25594 8740 25616
rect 1104 25542 1950 25594
rect 2002 25542 2014 25594
rect 2066 25542 2078 25594
rect 2130 25542 2142 25594
rect 2194 25542 2206 25594
rect 2258 25542 7950 25594
rect 8002 25542 8014 25594
rect 8066 25542 8078 25594
rect 8130 25542 8142 25594
rect 8194 25542 8206 25594
rect 8258 25542 8740 25594
rect 1104 25520 8740 25542
rect 1854 25440 1860 25492
rect 1912 25440 1918 25492
rect 7377 25483 7435 25489
rect 7377 25449 7389 25483
rect 7423 25480 7435 25483
rect 7742 25480 7748 25492
rect 7423 25452 7748 25480
rect 7423 25449 7435 25452
rect 7377 25443 7435 25449
rect 7742 25440 7748 25452
rect 7800 25440 7806 25492
rect 9306 25344 9312 25356
rect 7208 25316 9312 25344
rect 1670 25236 1676 25288
rect 1728 25236 1734 25288
rect 7208 25285 7236 25316
rect 9306 25304 9312 25316
rect 9364 25304 9370 25356
rect 7193 25279 7251 25285
rect 7193 25245 7205 25279
rect 7239 25245 7251 25279
rect 7193 25239 7251 25245
rect 7742 25236 7748 25288
rect 7800 25236 7806 25288
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25245 8171 25279
rect 8113 25239 8171 25245
rect 3050 25168 3056 25220
rect 3108 25168 3114 25220
rect 6454 25168 6460 25220
rect 6512 25208 6518 25220
rect 8128 25208 8156 25239
rect 6512 25180 8156 25208
rect 6512 25168 6518 25180
rect 7926 25100 7932 25152
rect 7984 25100 7990 25152
rect 8294 25100 8300 25152
rect 8352 25100 8358 25152
rect 1104 25050 8740 25072
rect 1104 24998 3010 25050
rect 3062 24998 3074 25050
rect 3126 24998 3138 25050
rect 3190 24998 3202 25050
rect 3254 24998 3266 25050
rect 3318 24998 8740 25050
rect 1104 24976 8740 24998
rect 2406 24828 2412 24880
rect 2464 24868 2470 24880
rect 6362 24868 6368 24880
rect 2464 24840 6368 24868
rect 2464 24828 2470 24840
rect 6362 24828 6368 24840
rect 6420 24828 6426 24880
rect 7006 24760 7012 24812
rect 7064 24760 7070 24812
rect 7285 24803 7343 24809
rect 7285 24769 7297 24803
rect 7331 24800 7343 24803
rect 7745 24803 7803 24809
rect 7331 24772 7604 24800
rect 7331 24769 7343 24772
rect 7285 24763 7343 24769
rect 7098 24624 7104 24676
rect 7156 24664 7162 24676
rect 7193 24667 7251 24673
rect 7193 24664 7205 24667
rect 7156 24636 7205 24664
rect 7156 24624 7162 24636
rect 7193 24633 7205 24636
rect 7239 24633 7251 24667
rect 7193 24627 7251 24633
rect 7466 24624 7472 24676
rect 7524 24624 7530 24676
rect 7576 24664 7604 24772
rect 7745 24769 7757 24803
rect 7791 24800 7803 24803
rect 7834 24800 7840 24812
rect 7791 24772 7840 24800
rect 7791 24769 7803 24772
rect 7745 24763 7803 24769
rect 7834 24760 7840 24772
rect 7892 24760 7898 24812
rect 8113 24803 8171 24809
rect 8113 24769 8125 24803
rect 8159 24769 8171 24803
rect 8113 24763 8171 24769
rect 7650 24692 7656 24744
rect 7708 24732 7714 24744
rect 8128 24732 8156 24763
rect 7708 24704 8156 24732
rect 7708 24692 7714 24704
rect 9582 24664 9588 24676
rect 7576 24636 9588 24664
rect 9582 24624 9588 24636
rect 9640 24624 9646 24676
rect 7834 24556 7840 24608
rect 7892 24596 7898 24608
rect 7929 24599 7987 24605
rect 7929 24596 7941 24599
rect 7892 24568 7941 24596
rect 7892 24556 7898 24568
rect 7929 24565 7941 24568
rect 7975 24565 7987 24599
rect 7929 24559 7987 24565
rect 8297 24599 8355 24605
rect 8297 24565 8309 24599
rect 8343 24596 8355 24599
rect 9030 24596 9036 24608
rect 8343 24568 9036 24596
rect 8343 24565 8355 24568
rect 8297 24559 8355 24565
rect 9030 24556 9036 24568
rect 9088 24556 9094 24608
rect 1104 24506 8740 24528
rect 1104 24454 1950 24506
rect 2002 24454 2014 24506
rect 2066 24454 2078 24506
rect 2130 24454 2142 24506
rect 2194 24454 2206 24506
rect 2258 24454 7950 24506
rect 8002 24454 8014 24506
rect 8066 24454 8078 24506
rect 8130 24454 8142 24506
rect 8194 24454 8206 24506
rect 8258 24454 8740 24506
rect 1104 24432 8740 24454
rect 3418 24352 3424 24404
rect 3476 24352 3482 24404
rect 5074 24352 5080 24404
rect 5132 24352 5138 24404
rect 7190 24352 7196 24404
rect 7248 24392 7254 24404
rect 7466 24392 7472 24404
rect 7248 24364 7472 24392
rect 7248 24352 7254 24364
rect 7466 24352 7472 24364
rect 7524 24352 7530 24404
rect 7650 24352 7656 24404
rect 7708 24352 7714 24404
rect 3694 24324 3700 24336
rect 3436 24296 3700 24324
rect 3436 24268 3464 24296
rect 3694 24284 3700 24296
rect 3752 24284 3758 24336
rect 3418 24216 3424 24268
rect 3476 24216 3482 24268
rect 9398 24256 9404 24268
rect 7484 24228 9404 24256
rect 3605 24191 3663 24197
rect 3605 24157 3617 24191
rect 3651 24188 3663 24191
rect 3694 24188 3700 24200
rect 3651 24160 3700 24188
rect 3651 24157 3663 24160
rect 3605 24151 3663 24157
rect 3694 24148 3700 24160
rect 3752 24148 3758 24200
rect 4893 24191 4951 24197
rect 4893 24157 4905 24191
rect 4939 24188 4951 24191
rect 4982 24188 4988 24200
rect 4939 24160 4988 24188
rect 4939 24157 4951 24160
rect 4893 24151 4951 24157
rect 4982 24148 4988 24160
rect 5040 24148 5046 24200
rect 7484 24197 7512 24228
rect 9398 24216 9404 24228
rect 9456 24216 9462 24268
rect 7469 24191 7527 24197
rect 7469 24157 7481 24191
rect 7515 24157 7527 24191
rect 7469 24151 7527 24157
rect 7745 24191 7803 24197
rect 7745 24157 7757 24191
rect 7791 24157 7803 24191
rect 8113 24191 8171 24197
rect 8113 24188 8125 24191
rect 7745 24151 7803 24157
rect 7852 24160 8125 24188
rect 7006 24080 7012 24132
rect 7064 24080 7070 24132
rect 7098 24080 7104 24132
rect 7156 24120 7162 24132
rect 7760 24120 7788 24151
rect 7156 24092 7788 24120
rect 7156 24080 7162 24092
rect 6362 24012 6368 24064
rect 6420 24052 6426 24064
rect 7852 24052 7880 24160
rect 8113 24157 8125 24160
rect 8159 24157 8171 24191
rect 8113 24151 8171 24157
rect 6420 24024 7880 24052
rect 6420 24012 6426 24024
rect 7926 24012 7932 24064
rect 7984 24012 7990 24064
rect 8294 24012 8300 24064
rect 8352 24012 8358 24064
rect 1104 23962 8740 23984
rect 1104 23910 3010 23962
rect 3062 23910 3074 23962
rect 3126 23910 3138 23962
rect 3190 23910 3202 23962
rect 3254 23910 3266 23962
rect 3318 23910 8740 23962
rect 1104 23888 8740 23910
rect 1578 23808 1584 23860
rect 1636 23848 1642 23860
rect 1765 23851 1823 23857
rect 1765 23848 1777 23851
rect 1636 23820 1777 23848
rect 1636 23808 1642 23820
rect 1765 23817 1777 23820
rect 1811 23817 1823 23851
rect 1765 23811 1823 23817
rect 7006 23808 7012 23860
rect 7064 23848 7070 23860
rect 7190 23848 7196 23860
rect 7064 23820 7196 23848
rect 7064 23808 7070 23820
rect 7190 23808 7196 23820
rect 7248 23808 7254 23860
rect 1394 23672 1400 23724
rect 1452 23712 1458 23724
rect 1949 23715 2007 23721
rect 1949 23712 1961 23715
rect 1452 23684 1961 23712
rect 1452 23672 1458 23684
rect 1949 23681 1961 23684
rect 1995 23681 2007 23715
rect 1949 23675 2007 23681
rect 5258 23672 5264 23724
rect 5316 23712 5322 23724
rect 7745 23715 7803 23721
rect 7745 23712 7757 23715
rect 5316 23684 7757 23712
rect 5316 23672 5322 23684
rect 7745 23681 7757 23684
rect 7791 23681 7803 23715
rect 7745 23675 7803 23681
rect 7834 23672 7840 23724
rect 7892 23712 7898 23724
rect 8113 23715 8171 23721
rect 8113 23712 8125 23715
rect 7892 23684 8125 23712
rect 7892 23672 7898 23684
rect 8113 23681 8125 23684
rect 8159 23681 8171 23715
rect 8113 23675 8171 23681
rect 1026 23536 1032 23588
rect 1084 23576 1090 23588
rect 6270 23576 6276 23588
rect 1084 23548 6276 23576
rect 1084 23536 1090 23548
rect 6270 23536 6276 23548
rect 6328 23536 6334 23588
rect 7929 23579 7987 23585
rect 7929 23545 7941 23579
rect 7975 23576 7987 23579
rect 8846 23576 8852 23588
rect 7975 23548 8852 23576
rect 7975 23545 7987 23548
rect 7929 23539 7987 23545
rect 8846 23536 8852 23548
rect 8904 23536 8910 23588
rect 4982 23468 4988 23520
rect 5040 23468 5046 23520
rect 8297 23511 8355 23517
rect 8297 23477 8309 23511
rect 8343 23508 8355 23511
rect 9030 23508 9036 23520
rect 8343 23480 9036 23508
rect 8343 23477 8355 23480
rect 8297 23471 8355 23477
rect 9030 23468 9036 23480
rect 9088 23468 9094 23520
rect 1104 23418 8740 23440
rect 1104 23366 1950 23418
rect 2002 23366 2014 23418
rect 2066 23366 2078 23418
rect 2130 23366 2142 23418
rect 2194 23366 2206 23418
rect 2258 23366 7950 23418
rect 8002 23366 8014 23418
rect 8066 23366 8078 23418
rect 8130 23366 8142 23418
rect 8194 23366 8206 23418
rect 8258 23366 8740 23418
rect 1104 23344 8740 23366
rect 7653 23307 7711 23313
rect 7653 23273 7665 23307
rect 7699 23304 7711 23307
rect 7834 23304 7840 23316
rect 7699 23276 7840 23304
rect 7699 23273 7711 23276
rect 7653 23267 7711 23273
rect 7834 23264 7840 23276
rect 7892 23264 7898 23316
rect 7469 23103 7527 23109
rect 7469 23069 7481 23103
rect 7515 23100 7527 23103
rect 7650 23100 7656 23112
rect 7515 23072 7656 23100
rect 7515 23069 7527 23072
rect 7469 23063 7527 23069
rect 7650 23060 7656 23072
rect 7708 23060 7714 23112
rect 7745 23103 7803 23109
rect 7745 23069 7757 23103
rect 7791 23069 7803 23103
rect 7745 23063 7803 23069
rect 7190 22992 7196 23044
rect 7248 23032 7254 23044
rect 7760 23032 7788 23063
rect 8110 23060 8116 23112
rect 8168 23060 8174 23112
rect 7248 23004 7788 23032
rect 7248 22992 7254 23004
rect 7926 22924 7932 22976
rect 7984 22924 7990 22976
rect 8294 22924 8300 22976
rect 8352 22924 8358 22976
rect 1104 22874 8740 22896
rect 1104 22822 3010 22874
rect 3062 22822 3074 22874
rect 3126 22822 3138 22874
rect 3190 22822 3202 22874
rect 3254 22822 3266 22874
rect 3318 22822 8740 22874
rect 1104 22800 8740 22822
rect 3786 22720 3792 22772
rect 3844 22720 3850 22772
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 7193 22763 7251 22769
rect 7193 22760 7205 22763
rect 6972 22732 7205 22760
rect 6972 22720 6978 22732
rect 7193 22729 7205 22732
rect 7239 22729 7251 22763
rect 7193 22723 7251 22729
rect 7561 22763 7619 22769
rect 7561 22729 7573 22763
rect 7607 22760 7619 22763
rect 7650 22760 7656 22772
rect 7607 22732 7656 22760
rect 7607 22729 7619 22732
rect 7561 22723 7619 22729
rect 7650 22720 7656 22732
rect 7708 22720 7714 22772
rect 2682 22652 2688 22704
rect 2740 22692 2746 22704
rect 2740 22664 7788 22692
rect 2740 22652 2746 22664
rect 934 22584 940 22636
rect 992 22624 998 22636
rect 1857 22627 1915 22633
rect 1857 22624 1869 22627
rect 992 22596 1869 22624
rect 992 22584 998 22596
rect 1857 22593 1869 22596
rect 1903 22593 1915 22627
rect 1857 22587 1915 22593
rect 3605 22627 3663 22633
rect 3605 22593 3617 22627
rect 3651 22624 3663 22627
rect 3970 22624 3976 22636
rect 3651 22596 3976 22624
rect 3651 22593 3663 22596
rect 3605 22587 3663 22593
rect 3970 22584 3976 22596
rect 4028 22584 4034 22636
rect 7009 22627 7067 22633
rect 7009 22593 7021 22627
rect 7055 22624 7067 22627
rect 7650 22624 7656 22636
rect 7055 22596 7656 22624
rect 7055 22593 7067 22596
rect 7009 22587 7067 22593
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 7760 22633 7788 22664
rect 7745 22627 7803 22633
rect 7745 22593 7757 22627
rect 7791 22593 7803 22627
rect 7745 22587 7803 22593
rect 8113 22627 8171 22633
rect 8113 22593 8125 22627
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 5810 22516 5816 22568
rect 5868 22556 5874 22568
rect 8128 22556 8156 22587
rect 5868 22528 8156 22556
rect 5868 22516 5874 22528
rect 2041 22491 2099 22497
rect 2041 22457 2053 22491
rect 2087 22488 2099 22491
rect 6178 22488 6184 22500
rect 2087 22460 6184 22488
rect 2087 22457 2099 22460
rect 2041 22451 2099 22457
rect 6178 22448 6184 22460
rect 6236 22448 6242 22500
rect 7006 22448 7012 22500
rect 7064 22488 7070 22500
rect 7282 22488 7288 22500
rect 7064 22460 7288 22488
rect 7064 22448 7070 22460
rect 7282 22448 7288 22460
rect 7340 22448 7346 22500
rect 7834 22380 7840 22432
rect 7892 22420 7898 22432
rect 7929 22423 7987 22429
rect 7929 22420 7941 22423
rect 7892 22392 7941 22420
rect 7892 22380 7898 22392
rect 7929 22389 7941 22392
rect 7975 22389 7987 22423
rect 7929 22383 7987 22389
rect 8297 22423 8355 22429
rect 8297 22389 8309 22423
rect 8343 22420 8355 22423
rect 9030 22420 9036 22432
rect 8343 22392 9036 22420
rect 8343 22389 8355 22392
rect 8297 22383 8355 22389
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 1104 22330 8740 22352
rect 1104 22278 1950 22330
rect 2002 22278 2014 22330
rect 2066 22278 2078 22330
rect 2130 22278 2142 22330
rect 2194 22278 2206 22330
rect 2258 22278 7950 22330
rect 8002 22278 8014 22330
rect 8066 22278 8078 22330
rect 8130 22278 8142 22330
rect 8194 22278 8206 22330
rect 8258 22278 8740 22330
rect 1104 22256 8740 22278
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 6454 22216 6460 22228
rect 6236 22188 6460 22216
rect 6236 22176 6242 22188
rect 6454 22176 6460 22188
rect 6512 22176 6518 22228
rect 7374 22176 7380 22228
rect 7432 22216 7438 22228
rect 8386 22216 8392 22228
rect 7432 22188 8392 22216
rect 7432 22176 7438 22188
rect 8386 22176 8392 22188
rect 8444 22176 8450 22228
rect 7101 22151 7159 22157
rect 7101 22117 7113 22151
rect 7147 22148 7159 22151
rect 7650 22148 7656 22160
rect 7147 22120 7656 22148
rect 7147 22117 7159 22120
rect 7101 22111 7159 22117
rect 7650 22108 7656 22120
rect 7708 22148 7714 22160
rect 8202 22148 8208 22160
rect 7708 22120 8208 22148
rect 7708 22108 7714 22120
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 6564 22052 8156 22080
rect 6564 22024 6592 22052
rect 4522 21972 4528 22024
rect 4580 21972 4586 22024
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 6730 21972 6736 22024
rect 6788 21972 6794 22024
rect 7285 22015 7343 22021
rect 7285 21981 7297 22015
rect 7331 22012 7343 22015
rect 7374 22012 7380 22024
rect 7331 21984 7380 22012
rect 7331 21981 7343 21984
rect 7285 21975 7343 21981
rect 7374 21972 7380 21984
rect 7432 21972 7438 22024
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 22012 7803 22015
rect 8018 22012 8024 22024
rect 7791 21984 8024 22012
rect 7791 21981 7803 21984
rect 7745 21975 7803 21981
rect 8018 21972 8024 21984
rect 8076 21972 8082 22024
rect 8128 22021 8156 22052
rect 8113 22015 8171 22021
rect 8113 21981 8125 22015
rect 8159 21981 8171 22015
rect 8113 21975 8171 21981
rect 5902 21904 5908 21956
rect 5960 21944 5966 21956
rect 5960 21916 7512 21944
rect 5960 21904 5966 21916
rect 4706 21836 4712 21888
rect 4764 21836 4770 21888
rect 6822 21836 6828 21888
rect 6880 21876 6886 21888
rect 7484 21885 7512 21916
rect 6917 21879 6975 21885
rect 6917 21876 6929 21879
rect 6880 21848 6929 21876
rect 6880 21836 6886 21848
rect 6917 21845 6929 21848
rect 6963 21845 6975 21879
rect 6917 21839 6975 21845
rect 7469 21879 7527 21885
rect 7469 21845 7481 21879
rect 7515 21845 7527 21879
rect 7469 21839 7527 21845
rect 7926 21836 7932 21888
rect 7984 21836 7990 21888
rect 8294 21836 8300 21888
rect 8352 21836 8358 21888
rect 1104 21786 8740 21808
rect 1104 21734 3010 21786
rect 3062 21734 3074 21786
rect 3126 21734 3138 21786
rect 3190 21734 3202 21786
rect 3254 21734 3266 21786
rect 3318 21734 8740 21786
rect 1104 21712 8740 21734
rect 1765 21675 1823 21681
rect 1765 21641 1777 21675
rect 1811 21672 1823 21675
rect 3510 21672 3516 21684
rect 1811 21644 3516 21672
rect 1811 21641 1823 21644
rect 1765 21635 1823 21641
rect 3510 21632 3516 21644
rect 3568 21632 3574 21684
rect 7374 21632 7380 21684
rect 7432 21632 7438 21684
rect 750 21496 756 21548
rect 808 21536 814 21548
rect 1581 21539 1639 21545
rect 1581 21536 1593 21539
rect 808 21508 1593 21536
rect 808 21496 814 21508
rect 1581 21505 1593 21508
rect 1627 21505 1639 21539
rect 7745 21539 7803 21545
rect 7745 21536 7757 21539
rect 1581 21499 1639 21505
rect 6886 21508 7757 21536
rect 3786 21428 3792 21480
rect 3844 21468 3850 21480
rect 6886 21468 6914 21508
rect 7745 21505 7757 21508
rect 7791 21505 7803 21539
rect 7745 21499 7803 21505
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 3844 21440 6914 21468
rect 3844 21428 3850 21440
rect 7374 21428 7380 21480
rect 7432 21468 7438 21480
rect 8128 21468 8156 21499
rect 7432 21440 8156 21468
rect 7432 21428 7438 21440
rect 3697 21335 3755 21341
rect 3697 21301 3709 21335
rect 3743 21332 3755 21335
rect 3970 21332 3976 21344
rect 3743 21304 3976 21332
rect 3743 21301 3755 21304
rect 3697 21295 3755 21301
rect 3970 21292 3976 21304
rect 4028 21292 4034 21344
rect 5442 21292 5448 21344
rect 5500 21332 5506 21344
rect 7285 21335 7343 21341
rect 7285 21332 7297 21335
rect 5500 21304 7297 21332
rect 5500 21292 5506 21304
rect 7285 21301 7297 21304
rect 7331 21301 7343 21335
rect 7285 21295 7343 21301
rect 7834 21292 7840 21344
rect 7892 21332 7898 21344
rect 7929 21335 7987 21341
rect 7929 21332 7941 21335
rect 7892 21304 7941 21332
rect 7892 21292 7898 21304
rect 7929 21301 7941 21304
rect 7975 21301 7987 21335
rect 7929 21295 7987 21301
rect 8297 21335 8355 21341
rect 8297 21301 8309 21335
rect 8343 21332 8355 21335
rect 9030 21332 9036 21344
rect 8343 21304 9036 21332
rect 8343 21301 8355 21304
rect 8297 21295 8355 21301
rect 9030 21292 9036 21304
rect 9088 21292 9094 21344
rect 1104 21242 8740 21264
rect 1104 21190 1950 21242
rect 2002 21190 2014 21242
rect 2066 21190 2078 21242
rect 2130 21190 2142 21242
rect 2194 21190 2206 21242
rect 2258 21190 7950 21242
rect 8002 21190 8014 21242
rect 8066 21190 8078 21242
rect 8130 21190 8142 21242
rect 8194 21190 8206 21242
rect 8258 21190 8740 21242
rect 1104 21168 8740 21190
rect 6914 21088 6920 21140
rect 6972 21088 6978 21140
rect 7929 21063 7987 21069
rect 7929 21029 7941 21063
rect 7975 21060 7987 21063
rect 8846 21060 8852 21072
rect 7975 21032 8852 21060
rect 7975 21029 7987 21032
rect 7929 21023 7987 21029
rect 8846 21020 8852 21032
rect 8904 21020 8910 21072
rect 290 20884 296 20936
rect 348 20924 354 20936
rect 1670 20924 1676 20936
rect 348 20896 1676 20924
rect 348 20884 354 20896
rect 1670 20884 1676 20896
rect 1728 20884 1734 20936
rect 6730 20884 6736 20936
rect 6788 20884 6794 20936
rect 7742 20884 7748 20936
rect 7800 20884 7806 20936
rect 8110 20884 8116 20936
rect 8168 20884 8174 20936
rect 6546 20748 6552 20800
rect 6604 20788 6610 20800
rect 6822 20788 6828 20800
rect 6604 20760 6828 20788
rect 6604 20748 6610 20760
rect 6822 20748 6828 20760
rect 6880 20748 6886 20800
rect 8294 20748 8300 20800
rect 8352 20748 8358 20800
rect 1104 20698 8740 20720
rect 1104 20646 3010 20698
rect 3062 20646 3074 20698
rect 3126 20646 3138 20698
rect 3190 20646 3202 20698
rect 3254 20646 3266 20698
rect 3318 20646 8740 20698
rect 1104 20624 8740 20646
rect 5258 20544 5264 20596
rect 5316 20544 5322 20596
rect 5534 20544 5540 20596
rect 5592 20544 5598 20596
rect 5074 20408 5080 20460
rect 5132 20408 5138 20460
rect 5350 20408 5356 20460
rect 5408 20408 5414 20460
rect 7742 20408 7748 20460
rect 7800 20408 7806 20460
rect 8110 20408 8116 20460
rect 8168 20408 8174 20460
rect 7834 20204 7840 20256
rect 7892 20244 7898 20256
rect 7929 20247 7987 20253
rect 7929 20244 7941 20247
rect 7892 20216 7941 20244
rect 7892 20204 7898 20216
rect 7929 20213 7941 20216
rect 7975 20213 7987 20247
rect 7929 20207 7987 20213
rect 8297 20247 8355 20253
rect 8297 20213 8309 20247
rect 8343 20244 8355 20247
rect 9030 20244 9036 20256
rect 8343 20216 9036 20244
rect 8343 20213 8355 20216
rect 8297 20207 8355 20213
rect 9030 20204 9036 20216
rect 9088 20204 9094 20256
rect 1104 20154 8740 20176
rect 1104 20102 1950 20154
rect 2002 20102 2014 20154
rect 2066 20102 2078 20154
rect 2130 20102 2142 20154
rect 2194 20102 2206 20154
rect 2258 20102 7950 20154
rect 8002 20102 8014 20154
rect 8066 20102 8078 20154
rect 8130 20102 8142 20154
rect 8194 20102 8206 20154
rect 8258 20102 8740 20154
rect 1104 20080 8740 20102
rect 2590 20000 2596 20052
rect 2648 20000 2654 20052
rect 4890 20000 4896 20052
rect 4948 20000 4954 20052
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 7190 20040 7196 20052
rect 6972 20012 7196 20040
rect 6972 20000 6978 20012
rect 7190 20000 7196 20012
rect 7248 20000 7254 20052
rect 7558 20000 7564 20052
rect 7616 20040 7622 20052
rect 7926 20040 7932 20052
rect 7616 20012 7932 20040
rect 7616 20000 7622 20012
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 7190 19864 7196 19916
rect 7248 19904 7254 19916
rect 7248 19876 8156 19904
rect 7248 19864 7254 19876
rect 1670 19796 1676 19848
rect 1728 19836 1734 19848
rect 2409 19839 2467 19845
rect 2409 19836 2421 19839
rect 1728 19808 2421 19836
rect 1728 19796 1734 19808
rect 2409 19805 2421 19808
rect 2455 19805 2467 19839
rect 2409 19799 2467 19805
rect 4430 19796 4436 19848
rect 4488 19836 4494 19848
rect 4709 19839 4767 19845
rect 4709 19836 4721 19839
rect 4488 19808 4721 19836
rect 4488 19796 4494 19808
rect 4709 19805 4721 19808
rect 4755 19805 4767 19839
rect 4709 19799 4767 19805
rect 5902 19796 5908 19848
rect 5960 19836 5966 19848
rect 8128 19845 8156 19876
rect 7745 19839 7803 19845
rect 7745 19836 7757 19839
rect 5960 19808 7757 19836
rect 5960 19796 5966 19808
rect 7745 19805 7757 19808
rect 7791 19805 7803 19839
rect 7745 19799 7803 19805
rect 8113 19839 8171 19845
rect 8113 19805 8125 19839
rect 8159 19805 8171 19839
rect 8113 19799 8171 19805
rect 3878 19660 3884 19712
rect 3936 19700 3942 19712
rect 7558 19700 7564 19712
rect 3936 19672 7564 19700
rect 3936 19660 3942 19672
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 7926 19660 7932 19712
rect 7984 19660 7990 19712
rect 8294 19660 8300 19712
rect 8352 19660 8358 19712
rect 1104 19610 8740 19632
rect 1104 19558 3010 19610
rect 3062 19558 3074 19610
rect 3126 19558 3138 19610
rect 3190 19558 3202 19610
rect 3254 19558 3266 19610
rect 3318 19558 8740 19610
rect 1104 19536 8740 19558
rect 1857 19499 1915 19505
rect 1857 19465 1869 19499
rect 1903 19496 1915 19499
rect 3418 19496 3424 19508
rect 1903 19468 3424 19496
rect 1903 19465 1915 19468
rect 1857 19459 1915 19465
rect 3418 19456 3424 19468
rect 3476 19456 3482 19508
rect 3510 19456 3516 19508
rect 3568 19456 3574 19508
rect 3602 19456 3608 19508
rect 3660 19456 3666 19508
rect 6638 19456 6644 19508
rect 6696 19456 6702 19508
rect 7466 19456 7472 19508
rect 7524 19496 7530 19508
rect 7653 19499 7711 19505
rect 7653 19496 7665 19499
rect 7524 19468 7665 19496
rect 7524 19456 7530 19468
rect 7653 19465 7665 19468
rect 7699 19465 7711 19499
rect 7653 19459 7711 19465
rect 7837 19499 7895 19505
rect 7837 19465 7849 19499
rect 7883 19496 7895 19499
rect 8297 19499 8355 19505
rect 7883 19468 8248 19496
rect 7883 19465 7895 19468
rect 7837 19459 7895 19465
rect 5258 19388 5264 19440
rect 5316 19428 5322 19440
rect 8220 19428 8248 19468
rect 8297 19465 8309 19499
rect 8343 19496 8355 19499
rect 9030 19496 9036 19508
rect 8343 19468 9036 19496
rect 8343 19465 8355 19468
rect 8297 19459 8355 19465
rect 9030 19456 9036 19468
rect 9088 19456 9094 19508
rect 8754 19428 8760 19440
rect 5316 19400 8156 19428
rect 8220 19400 8760 19428
rect 5316 19388 5322 19400
rect 1118 19320 1124 19372
rect 1176 19360 1182 19372
rect 1673 19363 1731 19369
rect 1673 19360 1685 19363
rect 1176 19332 1685 19360
rect 1176 19320 1182 19332
rect 1673 19329 1685 19332
rect 1719 19329 1731 19363
rect 1673 19323 1731 19329
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3418 19360 3424 19372
rect 3375 19332 3424 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 3510 19320 3516 19372
rect 3568 19360 3574 19372
rect 3789 19363 3847 19369
rect 3789 19360 3801 19363
rect 3568 19332 3801 19360
rect 3568 19320 3574 19332
rect 3789 19329 3801 19332
rect 3835 19329 3847 19363
rect 3789 19323 3847 19329
rect 6454 19320 6460 19372
rect 6512 19320 6518 19372
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 7484 19292 7512 19323
rect 7558 19320 7564 19372
rect 7616 19360 7622 19372
rect 8128 19369 8156 19400
rect 8754 19388 8760 19400
rect 8812 19388 8818 19440
rect 8021 19363 8079 19369
rect 8021 19360 8033 19363
rect 7616 19332 8033 19360
rect 7616 19320 7622 19332
rect 8021 19329 8033 19332
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 8113 19363 8171 19369
rect 8113 19329 8125 19363
rect 8159 19329 8171 19363
rect 8113 19323 8171 19329
rect 8386 19292 8392 19304
rect 7484 19264 8392 19292
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 7466 19184 7472 19236
rect 7524 19224 7530 19236
rect 8202 19224 8208 19236
rect 7524 19196 8208 19224
rect 7524 19184 7530 19196
rect 8202 19184 8208 19196
rect 8260 19184 8266 19236
rect 1104 19066 8740 19088
rect 1104 19014 1950 19066
rect 2002 19014 2014 19066
rect 2066 19014 2078 19066
rect 2130 19014 2142 19066
rect 2194 19014 2206 19066
rect 2258 19014 7950 19066
rect 8002 19014 8014 19066
rect 8066 19014 8078 19066
rect 8130 19014 8142 19066
rect 8194 19014 8206 19066
rect 8258 19014 8740 19066
rect 1104 18992 8740 19014
rect 7282 18912 7288 18964
rect 7340 18912 7346 18964
rect 7374 18912 7380 18964
rect 7432 18952 7438 18964
rect 7653 18955 7711 18961
rect 7653 18952 7665 18955
rect 7432 18924 7665 18952
rect 7432 18912 7438 18924
rect 7653 18921 7665 18924
rect 7699 18921 7711 18955
rect 7653 18915 7711 18921
rect 6270 18844 6276 18896
rect 6328 18884 6334 18896
rect 6328 18856 8156 18884
rect 6328 18844 6334 18856
rect 7484 18788 8064 18816
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 7282 18748 7288 18760
rect 7147 18720 7288 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 7282 18708 7288 18720
rect 7340 18708 7346 18760
rect 7484 18757 7512 18788
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18717 7527 18751
rect 7469 18711 7527 18717
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 7760 18680 7788 18711
rect 6886 18652 7788 18680
rect 8036 18680 8064 18788
rect 8128 18757 8156 18856
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18717 8171 18751
rect 8113 18711 8171 18717
rect 9674 18680 9680 18692
rect 8036 18652 9680 18680
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 6886 18612 6914 18652
rect 9674 18640 9680 18652
rect 9732 18640 9738 18692
rect 6144 18584 6914 18612
rect 6144 18572 6150 18584
rect 7926 18572 7932 18624
rect 7984 18572 7990 18624
rect 8294 18572 8300 18624
rect 8352 18572 8358 18624
rect 1104 18522 8740 18544
rect 1104 18470 3010 18522
rect 3062 18470 3074 18522
rect 3126 18470 3138 18522
rect 3190 18470 3202 18522
rect 3254 18470 3266 18522
rect 3318 18470 8740 18522
rect 1104 18448 8740 18470
rect 4798 18368 4804 18420
rect 4856 18368 4862 18420
rect 7098 18368 7104 18420
rect 7156 18408 7162 18420
rect 7377 18411 7435 18417
rect 7377 18408 7389 18411
rect 7156 18380 7389 18408
rect 7156 18368 7162 18380
rect 7377 18377 7389 18380
rect 7423 18377 7435 18411
rect 7377 18371 7435 18377
rect 7282 18300 7288 18352
rect 7340 18340 7346 18352
rect 9030 18340 9036 18352
rect 7340 18312 9036 18340
rect 7340 18300 7346 18312
rect 9030 18300 9036 18312
rect 9088 18300 9094 18352
rect 4614 18232 4620 18284
rect 4672 18232 4678 18284
rect 7193 18275 7251 18281
rect 7193 18241 7205 18275
rect 7239 18272 7251 18275
rect 8754 18272 8760 18284
rect 7239 18244 8760 18272
rect 7239 18241 7251 18244
rect 7193 18235 7251 18241
rect 8754 18232 8760 18244
rect 8812 18232 8818 18284
rect 1104 17978 8740 18000
rect 1104 17926 1950 17978
rect 2002 17926 2014 17978
rect 2066 17926 2078 17978
rect 2130 17926 2142 17978
rect 2194 17926 2206 17978
rect 2258 17926 7950 17978
rect 8002 17926 8014 17978
rect 8066 17926 8078 17978
rect 8130 17926 8142 17978
rect 8194 17926 8206 17978
rect 8258 17926 8740 17978
rect 1104 17904 8740 17926
rect 1762 17824 1768 17876
rect 1820 17824 1826 17876
rect 6362 17824 6368 17876
rect 6420 17864 6426 17876
rect 6825 17867 6883 17873
rect 6825 17864 6837 17867
rect 6420 17836 6837 17864
rect 6420 17824 6426 17836
rect 6825 17833 6837 17836
rect 6871 17833 6883 17867
rect 6825 17827 6883 17833
rect 6178 17688 6184 17740
rect 6236 17728 6242 17740
rect 6362 17728 6368 17740
rect 6236 17700 6368 17728
rect 6236 17688 6242 17700
rect 6362 17688 6368 17700
rect 6420 17688 6426 17740
rect 842 17620 848 17672
rect 900 17660 906 17672
rect 1581 17663 1639 17669
rect 1581 17660 1593 17663
rect 900 17632 1593 17660
rect 900 17620 906 17632
rect 1581 17629 1593 17632
rect 1627 17629 1639 17663
rect 1581 17623 1639 17629
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17660 6699 17663
rect 7650 17660 7656 17672
rect 6687 17632 7656 17660
rect 6687 17629 6699 17632
rect 6641 17623 6699 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 1104 17434 8740 17456
rect 1104 17382 3010 17434
rect 3062 17382 3074 17434
rect 3126 17382 3138 17434
rect 3190 17382 3202 17434
rect 3254 17382 3266 17434
rect 3318 17382 8740 17434
rect 1104 17360 8740 17382
rect 7006 17280 7012 17332
rect 7064 17320 7070 17332
rect 7101 17323 7159 17329
rect 7101 17320 7113 17323
rect 7064 17292 7113 17320
rect 7064 17280 7070 17292
rect 7101 17289 7113 17292
rect 7147 17289 7159 17323
rect 7101 17283 7159 17289
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17153 6975 17187
rect 6917 17147 6975 17153
rect 6932 17060 6960 17147
rect 6914 17008 6920 17060
rect 6972 17008 6978 17060
rect 1104 16890 8740 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 7950 16890
rect 8002 16838 8014 16890
rect 8066 16838 8078 16890
rect 8130 16838 8142 16890
rect 8194 16838 8206 16890
rect 8258 16838 8740 16890
rect 1104 16816 8740 16838
rect 1104 16346 8740 16368
rect 1104 16294 3010 16346
rect 3062 16294 3074 16346
rect 3126 16294 3138 16346
rect 3190 16294 3202 16346
rect 3254 16294 3266 16346
rect 3318 16294 8740 16346
rect 1104 16272 8740 16294
rect 1854 16192 1860 16244
rect 1912 16192 1918 16244
rect 4890 16192 4896 16244
rect 4948 16192 4954 16244
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6420 16204 6561 16232
rect 6420 16192 6426 16204
rect 6549 16201 6561 16204
rect 6595 16201 6607 16235
rect 6549 16195 6607 16201
rect 7558 16192 7564 16244
rect 7616 16192 7622 16244
rect 1210 16056 1216 16108
rect 1268 16096 1274 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 1268 16068 2053 16096
rect 1268 16056 1274 16068
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 4709 16099 4767 16105
rect 4709 16065 4721 16099
rect 4755 16096 4767 16099
rect 4890 16096 4896 16108
rect 4755 16068 4896 16096
rect 4755 16065 4767 16068
rect 4709 16059 4767 16065
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 6365 16099 6423 16105
rect 6365 16065 6377 16099
rect 6411 16096 6423 16099
rect 7377 16099 7435 16105
rect 6411 16068 6914 16096
rect 6411 16065 6423 16068
rect 6365 16059 6423 16065
rect 6886 16028 6914 16068
rect 7377 16065 7389 16099
rect 7423 16096 7435 16099
rect 8754 16096 8760 16108
rect 7423 16068 8760 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 8754 16056 8760 16068
rect 8812 16056 8818 16108
rect 8570 16028 8576 16040
rect 6886 16000 8576 16028
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 1104 15802 8740 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 7950 15802
rect 8002 15750 8014 15802
rect 8066 15750 8078 15802
rect 8130 15750 8142 15802
rect 8194 15750 8206 15802
rect 8258 15750 8740 15802
rect 1104 15728 8740 15750
rect 2225 15691 2283 15697
rect 2225 15657 2237 15691
rect 2271 15688 2283 15691
rect 2314 15688 2320 15700
rect 2271 15660 2320 15688
rect 2271 15657 2283 15660
rect 2225 15651 2283 15657
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 750 15444 756 15496
rect 808 15484 814 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 808 15456 2053 15484
rect 808 15444 814 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 1104 15258 8740 15280
rect 1104 15206 3010 15258
rect 3062 15206 3074 15258
rect 3126 15206 3138 15258
rect 3190 15206 3202 15258
rect 3254 15206 3266 15258
rect 3318 15206 8740 15258
rect 1104 15184 8740 15206
rect 6546 15104 6552 15156
rect 6604 15104 6610 15156
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 8478 15008 8484 15020
rect 6411 14980 8484 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 6914 14764 6920 14816
rect 6972 14804 6978 14816
rect 7926 14804 7932 14816
rect 6972 14776 7932 14804
rect 6972 14764 6978 14776
rect 7926 14764 7932 14776
rect 7984 14764 7990 14816
rect 1104 14714 8740 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 7950 14714
rect 8002 14662 8014 14714
rect 8066 14662 8078 14714
rect 8130 14662 8142 14714
rect 8194 14662 8206 14714
rect 8258 14662 8740 14714
rect 1104 14640 8740 14662
rect 2133 14603 2191 14609
rect 2133 14569 2145 14603
rect 2179 14600 2191 14603
rect 2406 14600 2412 14612
rect 2179 14572 2412 14600
rect 2179 14569 2191 14572
rect 2133 14563 2191 14569
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 6914 14560 6920 14612
rect 6972 14560 6978 14612
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 7524 14572 8125 14600
rect 7524 14560 7530 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 1026 14356 1032 14408
rect 1084 14396 1090 14408
rect 1949 14399 2007 14405
rect 1949 14396 1961 14399
rect 1084 14368 1961 14396
rect 1084 14356 1090 14368
rect 1949 14365 1961 14368
rect 1995 14365 2007 14399
rect 1949 14359 2007 14365
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14396 6791 14399
rect 7929 14399 7987 14405
rect 6779 14368 6914 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 6886 14328 6914 14368
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 9490 14396 9496 14408
rect 7975 14368 9496 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 9490 14356 9496 14368
rect 9548 14356 9554 14408
rect 8294 14328 8300 14340
rect 6886 14300 8300 14328
rect 8294 14288 8300 14300
rect 8352 14288 8358 14340
rect 1104 14170 8740 14192
rect 1104 14118 3010 14170
rect 3062 14118 3074 14170
rect 3126 14118 3138 14170
rect 3190 14118 3202 14170
rect 3254 14118 3266 14170
rect 3318 14118 8740 14170
rect 1104 14096 8740 14118
rect 1104 13626 8740 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 7950 13626
rect 8002 13574 8014 13626
rect 8066 13574 8078 13626
rect 8130 13574 8142 13626
rect 8194 13574 8206 13626
rect 8258 13574 8740 13626
rect 1104 13552 8740 13574
rect 1854 13472 1860 13524
rect 1912 13472 1918 13524
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 7892 13484 8033 13512
rect 7892 13472 7898 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 8021 13475 8079 13481
rect 750 13268 756 13320
rect 808 13308 814 13320
rect 1673 13311 1731 13317
rect 1673 13308 1685 13311
rect 808 13280 1685 13308
rect 808 13268 814 13280
rect 1673 13277 1685 13280
rect 1719 13277 1731 13311
rect 1673 13271 1731 13277
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13308 7895 13311
rect 8754 13308 8760 13320
rect 7883 13280 8760 13308
rect 7883 13277 7895 13280
rect 7837 13271 7895 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 1104 13082 8740 13104
rect 1104 13030 3010 13082
rect 3062 13030 3074 13082
rect 3126 13030 3138 13082
rect 3190 13030 3202 13082
rect 3254 13030 3266 13082
rect 3318 13030 8740 13082
rect 1104 13008 8740 13030
rect 1104 12538 8740 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 7950 12538
rect 8002 12486 8014 12538
rect 8066 12486 8078 12538
rect 8130 12486 8142 12538
rect 8194 12486 8206 12538
rect 8258 12486 8740 12538
rect 1104 12464 8740 12486
rect 2682 12384 2688 12436
rect 2740 12424 2746 12436
rect 5905 12427 5963 12433
rect 5905 12424 5917 12427
rect 2740 12396 5917 12424
rect 2740 12384 2746 12396
rect 5905 12393 5917 12396
rect 5951 12393 5963 12427
rect 5905 12387 5963 12393
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 7653 12427 7711 12433
rect 7653 12424 7665 12427
rect 6880 12396 7665 12424
rect 6880 12384 6886 12396
rect 7653 12393 7665 12396
rect 7699 12393 7711 12427
rect 7653 12387 7711 12393
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12220 5779 12223
rect 7469 12223 7527 12229
rect 5767 12192 6914 12220
rect 5767 12189 5779 12192
rect 5721 12183 5779 12189
rect 6886 12152 6914 12192
rect 7469 12189 7481 12223
rect 7515 12220 7527 12223
rect 8754 12220 8760 12232
rect 7515 12192 8760 12220
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 8478 12152 8484 12164
rect 6886 12124 8484 12152
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 1104 11994 8740 12016
rect 1104 11942 3010 11994
rect 3062 11942 3074 11994
rect 3126 11942 3138 11994
rect 3190 11942 3202 11994
rect 3254 11942 3266 11994
rect 3318 11942 8740 11994
rect 1104 11920 8740 11942
rect 7837 11883 7895 11889
rect 7837 11849 7849 11883
rect 7883 11880 7895 11883
rect 8386 11880 8392 11892
rect 7883 11852 8392 11880
rect 7883 11849 7895 11852
rect 7837 11843 7895 11849
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11744 8079 11747
rect 8938 11744 8944 11756
rect 8067 11716 8944 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 1104 11450 8740 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 7950 11450
rect 8002 11398 8014 11450
rect 8066 11398 8078 11450
rect 8130 11398 8142 11450
rect 8194 11398 8206 11450
rect 8258 11398 8740 11450
rect 1104 11376 8740 11398
rect 1854 11296 1860 11348
rect 1912 11296 1918 11348
rect 5810 11296 5816 11348
rect 5868 11296 5874 11348
rect 1118 11092 1124 11144
rect 1176 11132 1182 11144
rect 2041 11135 2099 11141
rect 2041 11132 2053 11135
rect 1176 11104 2053 11132
rect 1176 11092 1182 11104
rect 2041 11101 2053 11104
rect 2087 11101 2099 11135
rect 2041 11095 2099 11101
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11132 5687 11135
rect 8294 11132 8300 11144
rect 5675 11104 8300 11132
rect 5675 11101 5687 11104
rect 5629 11095 5687 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 1104 10906 8740 10928
rect 1104 10854 3010 10906
rect 3062 10854 3074 10906
rect 3126 10854 3138 10906
rect 3190 10854 3202 10906
rect 3254 10854 3266 10906
rect 3318 10854 8740 10906
rect 1104 10832 8740 10854
rect 6917 10795 6975 10801
rect 6917 10761 6929 10795
rect 6963 10792 6975 10795
rect 7006 10792 7012 10804
rect 6963 10764 7012 10792
rect 6963 10761 6975 10764
rect 6917 10755 6975 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 8386 10656 8392 10668
rect 6779 10628 8392 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 1104 10362 8740 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 7950 10362
rect 8002 10310 8014 10362
rect 8066 10310 8078 10362
rect 8130 10310 8142 10362
rect 8194 10310 8206 10362
rect 8258 10310 8740 10362
rect 1104 10288 8740 10310
rect 1104 9818 8740 9840
rect 1104 9766 3010 9818
rect 3062 9766 3074 9818
rect 3126 9766 3138 9818
rect 3190 9766 3202 9818
rect 3254 9766 3266 9818
rect 3318 9766 8740 9818
rect 1104 9744 8740 9766
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7098 9392 7104 9444
rect 7156 9392 7162 9444
rect 1104 9274 8740 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 7950 9274
rect 8002 9222 8014 9274
rect 8066 9222 8078 9274
rect 8130 9222 8142 9274
rect 8194 9222 8206 9274
rect 8258 9222 8740 9274
rect 1104 9200 8740 9222
rect 5166 9120 5172 9172
rect 5224 9160 5230 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 5224 9132 7297 9160
rect 5224 9120 5230 9132
rect 7285 9129 7297 9132
rect 7331 9129 7343 9163
rect 7285 9123 7343 9129
rect 7098 8916 7104 8968
rect 7156 8916 7162 8968
rect 1104 8730 8740 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 8740 8730
rect 1104 8656 8740 8678
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 5960 8588 6561 8616
rect 5960 8576 5966 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 6549 8579 6607 8585
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 8386 8480 8392 8492
rect 6411 8452 8392 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 1104 8186 8740 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 8740 8186
rect 1104 8112 8740 8134
rect 7190 8032 7196 8084
rect 7248 8032 7254 8084
rect 7006 7828 7012 7880
rect 7064 7828 7070 7880
rect 1104 7642 8740 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 8740 7642
rect 1104 7568 8740 7590
rect 1104 7098 8740 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 8740 7098
rect 1104 7024 8740 7046
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7892 6752 7941 6780
rect 7892 6740 7898 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 7742 6604 7748 6656
rect 7800 6604 7806 6656
rect 1104 6554 8740 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 8740 6554
rect 1104 6480 8740 6502
rect 7374 6400 7380 6452
rect 7432 6400 7438 6452
rect 7190 6264 7196 6316
rect 7248 6264 7254 6316
rect 1104 6010 8740 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 8740 6010
rect 1104 5936 8740 5958
rect 5994 5856 6000 5908
rect 6052 5856 6058 5908
rect 5810 5652 5816 5704
rect 5868 5652 5874 5704
rect 1104 5466 8740 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 8740 5466
rect 1104 5392 8740 5414
rect 1104 4922 8740 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 8740 4922
rect 1104 4848 8740 4870
rect 6178 4768 6184 4820
rect 6236 4768 6242 4820
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4604 6055 4607
rect 6730 4604 6736 4616
rect 6043 4576 6736 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 1104 4378 8740 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 8740 4378
rect 1104 4304 8740 4326
rect 7282 4088 7288 4140
rect 7340 4088 7346 4140
rect 3786 3952 3792 4004
rect 3844 3992 3850 4004
rect 7469 3995 7527 4001
rect 7469 3992 7481 3995
rect 3844 3964 7481 3992
rect 3844 3952 3850 3964
rect 7469 3961 7481 3964
rect 7515 3961 7527 3995
rect 7469 3955 7527 3961
rect 1104 3834 8740 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 8740 3834
rect 1104 3760 8740 3782
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 3936 3692 7941 3720
rect 3936 3680 3942 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 7892 3488 8125 3516
rect 7892 3476 7898 3488
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 3418 3408 3424 3460
rect 3476 3448 3482 3460
rect 6730 3448 6736 3460
rect 3476 3420 6736 3448
rect 3476 3408 3482 3420
rect 6730 3408 6736 3420
rect 6788 3408 6794 3460
rect 1104 3290 8740 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 8740 3290
rect 1104 3216 8740 3238
rect 6086 3136 6092 3188
rect 6144 3136 6150 3188
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6328 3148 6561 3176
rect 6328 3136 6334 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 5902 3000 5908 3052
rect 5960 3000 5966 3052
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7800 3012 7849 3040
rect 7800 3000 7806 3012
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 5258 2864 5264 2916
rect 5316 2904 5322 2916
rect 8021 2907 8079 2913
rect 8021 2904 8033 2907
rect 5316 2876 8033 2904
rect 5316 2864 5322 2876
rect 8021 2873 8033 2876
rect 8067 2873 8079 2907
rect 8021 2867 8079 2873
rect 1104 2746 8740 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 8740 2746
rect 1104 2672 8740 2694
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 2682 2632 2688 2644
rect 2188 2604 2688 2632
rect 2188 2592 2194 2604
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 8570 2632 8576 2644
rect 5500 2604 8576 2632
rect 5500 2592 5506 2604
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 1104 2202 8740 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 8740 2202
rect 1104 2128 8740 2150
rect 1670 2048 1676 2100
rect 1728 2088 1734 2100
rect 2590 2088 2596 2100
rect 1728 2060 2596 2088
rect 1728 2048 1734 2060
rect 2590 2048 2596 2060
rect 2648 2048 2654 2100
rect 4522 416 4528 468
rect 4580 456 4586 468
rect 6270 456 6276 468
rect 4580 428 6276 456
rect 4580 416 4586 428
rect 6270 416 6276 428
rect 6328 416 6334 468
<< via1 >>
rect 3010 42406 3062 42458
rect 3074 42406 3126 42458
rect 3138 42406 3190 42458
rect 3202 42406 3254 42458
rect 3266 42406 3318 42458
rect 1216 42304 1268 42356
rect 1676 42304 1728 42356
rect 2136 42304 2188 42356
rect 2596 42304 2648 42356
rect 2872 42304 2924 42356
rect 3516 42304 3568 42356
rect 3976 42304 4028 42356
rect 4436 42304 4488 42356
rect 4896 42304 4948 42356
rect 5356 42304 5408 42356
rect 5816 42304 5868 42356
rect 6276 42304 6328 42356
rect 6736 42304 6788 42356
rect 7196 42304 7248 42356
rect 7656 42304 7708 42356
rect 8116 42304 8168 42356
rect 4528 42236 4580 42288
rect 1676 42211 1728 42220
rect 1676 42177 1685 42211
rect 1685 42177 1719 42211
rect 1719 42177 1728 42211
rect 1676 42168 1728 42177
rect 1584 42100 1636 42152
rect 2596 42211 2648 42220
rect 2596 42177 2605 42211
rect 2605 42177 2639 42211
rect 2639 42177 2648 42211
rect 2596 42168 2648 42177
rect 3424 42168 3476 42220
rect 3608 42211 3660 42220
rect 3608 42177 3617 42211
rect 3617 42177 3651 42211
rect 3651 42177 3660 42211
rect 3608 42168 3660 42177
rect 3792 42168 3844 42220
rect 4896 42168 4948 42220
rect 4988 42211 5040 42220
rect 4988 42177 4997 42211
rect 4997 42177 5031 42211
rect 5031 42177 5040 42211
rect 4988 42168 5040 42177
rect 5632 42168 5684 42220
rect 5908 42211 5960 42220
rect 5908 42177 5917 42211
rect 5917 42177 5951 42211
rect 5951 42177 5960 42211
rect 5908 42168 5960 42177
rect 2688 42100 2740 42152
rect 4712 42100 4764 42152
rect 7012 42168 7064 42220
rect 5448 42032 5500 42084
rect 5080 41964 5132 42016
rect 1950 41862 2002 41914
rect 2014 41862 2066 41914
rect 2078 41862 2130 41914
rect 2142 41862 2194 41914
rect 2206 41862 2258 41914
rect 7950 41862 8002 41914
rect 8014 41862 8066 41914
rect 8078 41862 8130 41914
rect 8142 41862 8194 41914
rect 8206 41862 8258 41914
rect 296 41760 348 41812
rect 8576 41760 8628 41812
rect 756 41692 808 41744
rect 9036 41692 9088 41744
rect 6092 41624 6144 41676
rect 1676 41599 1728 41608
rect 1676 41565 1685 41599
rect 1685 41565 1719 41599
rect 1719 41565 1728 41599
rect 1676 41556 1728 41565
rect 1860 41556 1912 41608
rect 7472 41599 7524 41608
rect 7472 41565 7481 41599
rect 7481 41565 7515 41599
rect 7515 41565 7524 41599
rect 7472 41556 7524 41565
rect 7104 41488 7156 41540
rect 7840 41420 7892 41472
rect 3010 41318 3062 41370
rect 3074 41318 3126 41370
rect 3138 41318 3190 41370
rect 3202 41318 3254 41370
rect 3266 41318 3318 41370
rect 9496 41216 9548 41268
rect 7380 41080 7432 41132
rect 6736 41012 6788 41064
rect 7748 40919 7800 40928
rect 7748 40885 7757 40919
rect 7757 40885 7791 40919
rect 7791 40885 7800 40919
rect 7748 40876 7800 40885
rect 1950 40774 2002 40826
rect 2014 40774 2066 40826
rect 2078 40774 2130 40826
rect 2142 40774 2194 40826
rect 2206 40774 2258 40826
rect 7950 40774 8002 40826
rect 8014 40774 8066 40826
rect 8078 40774 8130 40826
rect 8142 40774 8194 40826
rect 8206 40774 8258 40826
rect 204 40468 256 40520
rect 7656 40511 7708 40520
rect 7656 40477 7665 40511
rect 7665 40477 7699 40511
rect 7699 40477 7708 40511
rect 7656 40468 7708 40477
rect 5724 40332 5776 40384
rect 7840 40375 7892 40384
rect 7840 40341 7849 40375
rect 7849 40341 7883 40375
rect 7883 40341 7892 40375
rect 7840 40332 7892 40341
rect 3010 40230 3062 40282
rect 3074 40230 3126 40282
rect 3138 40230 3190 40282
rect 3202 40230 3254 40282
rect 3266 40230 3318 40282
rect 7932 40060 7984 40112
rect 7748 40035 7800 40044
rect 7748 40001 7757 40035
rect 7757 40001 7791 40035
rect 7791 40001 7800 40035
rect 7748 39992 7800 40001
rect 7932 39899 7984 39908
rect 7932 39865 7941 39899
rect 7941 39865 7975 39899
rect 7975 39865 7984 39899
rect 7932 39856 7984 39865
rect 8300 39831 8352 39840
rect 8300 39797 8309 39831
rect 8309 39797 8343 39831
rect 8343 39797 8352 39831
rect 8300 39788 8352 39797
rect 1950 39686 2002 39738
rect 2014 39686 2066 39738
rect 2078 39686 2130 39738
rect 2142 39686 2194 39738
rect 2206 39686 2258 39738
rect 7950 39686 8002 39738
rect 8014 39686 8066 39738
rect 8078 39686 8130 39738
rect 8142 39686 8194 39738
rect 8206 39686 8258 39738
rect 112 39380 164 39432
rect 5540 39380 5592 39432
rect 7840 39380 7892 39432
rect 6000 39244 6052 39296
rect 7932 39287 7984 39296
rect 7932 39253 7941 39287
rect 7941 39253 7975 39287
rect 7975 39253 7984 39287
rect 7932 39244 7984 39253
rect 8300 39287 8352 39296
rect 8300 39253 8309 39287
rect 8309 39253 8343 39287
rect 8343 39253 8352 39287
rect 8300 39244 8352 39253
rect 3010 39142 3062 39194
rect 3074 39142 3126 39194
rect 3138 39142 3190 39194
rect 3202 39142 3254 39194
rect 3266 39142 3318 39194
rect 7748 38947 7800 38956
rect 7748 38913 7757 38947
rect 7757 38913 7791 38947
rect 7791 38913 7800 38947
rect 7748 38904 7800 38913
rect 7840 38904 7892 38956
rect 7932 38811 7984 38820
rect 7932 38777 7941 38811
rect 7941 38777 7975 38811
rect 7975 38777 7984 38811
rect 7932 38768 7984 38777
rect 8300 38743 8352 38752
rect 8300 38709 8309 38743
rect 8309 38709 8343 38743
rect 8343 38709 8352 38743
rect 8300 38700 8352 38709
rect 1950 38598 2002 38650
rect 2014 38598 2066 38650
rect 2078 38598 2130 38650
rect 2142 38598 2194 38650
rect 2206 38598 2258 38650
rect 7950 38598 8002 38650
rect 8014 38598 8066 38650
rect 8078 38598 8130 38650
rect 8142 38598 8194 38650
rect 8206 38598 8258 38650
rect 7748 38496 7800 38548
rect 5724 38360 5776 38412
rect 1308 38292 1360 38344
rect 5540 38292 5592 38344
rect 7748 38335 7800 38344
rect 7748 38301 7757 38335
rect 7757 38301 7791 38335
rect 7791 38301 7800 38335
rect 7748 38292 7800 38301
rect 6828 38156 6880 38208
rect 7932 38199 7984 38208
rect 7932 38165 7941 38199
rect 7941 38165 7975 38199
rect 7975 38165 7984 38199
rect 7932 38156 7984 38165
rect 8300 38199 8352 38208
rect 8300 38165 8309 38199
rect 8309 38165 8343 38199
rect 8343 38165 8352 38199
rect 8300 38156 8352 38165
rect 3010 38054 3062 38106
rect 3074 38054 3126 38106
rect 3138 38054 3190 38106
rect 3202 38054 3254 38106
rect 3266 38054 3318 38106
rect 7840 37952 7892 38004
rect 6000 37884 6052 37936
rect 7472 37859 7524 37868
rect 7472 37825 7481 37859
rect 7481 37825 7515 37859
rect 7515 37825 7524 37859
rect 7472 37816 7524 37825
rect 7656 37816 7708 37868
rect 7932 37723 7984 37732
rect 7932 37689 7941 37723
rect 7941 37689 7975 37723
rect 7975 37689 7984 37723
rect 7932 37680 7984 37689
rect 8300 37655 8352 37664
rect 8300 37621 8309 37655
rect 8309 37621 8343 37655
rect 8343 37621 8352 37655
rect 8300 37612 8352 37621
rect 1950 37510 2002 37562
rect 2014 37510 2066 37562
rect 2078 37510 2130 37562
rect 2142 37510 2194 37562
rect 2206 37510 2258 37562
rect 7950 37510 8002 37562
rect 8014 37510 8066 37562
rect 8078 37510 8130 37562
rect 8142 37510 8194 37562
rect 8206 37510 8258 37562
rect 7748 37408 7800 37460
rect 6920 37204 6972 37256
rect 6828 37136 6880 37188
rect 5724 37068 5776 37120
rect 7932 37111 7984 37120
rect 7932 37077 7941 37111
rect 7941 37077 7975 37111
rect 7975 37077 7984 37111
rect 7932 37068 7984 37077
rect 8300 37111 8352 37120
rect 8300 37077 8309 37111
rect 8309 37077 8343 37111
rect 8343 37077 8352 37111
rect 8300 37068 8352 37077
rect 3010 36966 3062 37018
rect 3074 36966 3126 37018
rect 3138 36966 3190 37018
rect 3202 36966 3254 37018
rect 3266 36966 3318 37018
rect 2412 36771 2464 36780
rect 2412 36737 2421 36771
rect 2421 36737 2455 36771
rect 2455 36737 2464 36771
rect 2412 36728 2464 36737
rect 3976 36660 4028 36712
rect 7932 36635 7984 36644
rect 7932 36601 7941 36635
rect 7941 36601 7975 36635
rect 7975 36601 7984 36635
rect 7932 36592 7984 36601
rect 8300 36567 8352 36576
rect 8300 36533 8309 36567
rect 8309 36533 8343 36567
rect 8343 36533 8352 36567
rect 8300 36524 8352 36533
rect 1950 36422 2002 36474
rect 2014 36422 2066 36474
rect 2078 36422 2130 36474
rect 2142 36422 2194 36474
rect 2206 36422 2258 36474
rect 7950 36422 8002 36474
rect 8014 36422 8066 36474
rect 8078 36422 8130 36474
rect 8142 36422 8194 36474
rect 8206 36422 8258 36474
rect 848 36116 900 36168
rect 5356 36048 5408 36100
rect 7932 36023 7984 36032
rect 7932 35989 7941 36023
rect 7941 35989 7975 36023
rect 7975 35989 7984 36023
rect 7932 35980 7984 35989
rect 8300 36023 8352 36032
rect 8300 35989 8309 36023
rect 8309 35989 8343 36023
rect 8343 35989 8352 36023
rect 8300 35980 8352 35989
rect 3010 35878 3062 35930
rect 3074 35878 3126 35930
rect 3138 35878 3190 35930
rect 3202 35878 3254 35930
rect 3266 35878 3318 35930
rect 4344 35640 4396 35692
rect 6184 35572 6236 35624
rect 7932 35547 7984 35556
rect 7932 35513 7941 35547
rect 7941 35513 7975 35547
rect 7975 35513 7984 35547
rect 7932 35504 7984 35513
rect 8300 35479 8352 35488
rect 8300 35445 8309 35479
rect 8309 35445 8343 35479
rect 8343 35445 8352 35479
rect 8300 35436 8352 35445
rect 1950 35334 2002 35386
rect 2014 35334 2066 35386
rect 2078 35334 2130 35386
rect 2142 35334 2194 35386
rect 2206 35334 2258 35386
rect 7950 35334 8002 35386
rect 8014 35334 8066 35386
rect 8078 35334 8130 35386
rect 8142 35334 8194 35386
rect 8206 35334 8258 35386
rect 5356 35232 5408 35284
rect 7656 35275 7708 35284
rect 7656 35241 7665 35275
rect 7665 35241 7699 35275
rect 7699 35241 7708 35275
rect 7656 35232 7708 35241
rect 3884 35096 3936 35148
rect 296 35028 348 35080
rect 7472 35071 7524 35080
rect 7472 35037 7481 35071
rect 7481 35037 7515 35071
rect 7515 35037 7524 35071
rect 7472 35028 7524 35037
rect 3700 34960 3752 35012
rect 7932 34935 7984 34944
rect 7932 34901 7941 34935
rect 7941 34901 7975 34935
rect 7975 34901 7984 34935
rect 7932 34892 7984 34901
rect 8300 34935 8352 34944
rect 8300 34901 8309 34935
rect 8309 34901 8343 34935
rect 8343 34901 8352 34935
rect 8300 34892 8352 34901
rect 3010 34790 3062 34842
rect 3074 34790 3126 34842
rect 3138 34790 3190 34842
rect 3202 34790 3254 34842
rect 3266 34790 3318 34842
rect 8852 34688 8904 34740
rect 1768 34552 1820 34604
rect 2320 34484 2372 34536
rect 8300 34391 8352 34400
rect 8300 34357 8309 34391
rect 8309 34357 8343 34391
rect 8343 34357 8352 34391
rect 8300 34348 8352 34357
rect 1950 34246 2002 34298
rect 2014 34246 2066 34298
rect 2078 34246 2130 34298
rect 2142 34246 2194 34298
rect 2206 34246 2258 34298
rect 7950 34246 8002 34298
rect 8014 34246 8066 34298
rect 8078 34246 8130 34298
rect 8142 34246 8194 34298
rect 8206 34246 8258 34298
rect 664 33940 716 33992
rect 6368 33940 6420 33992
rect 8116 33983 8168 33992
rect 8116 33949 8125 33983
rect 8125 33949 8159 33983
rect 8159 33949 8168 33983
rect 8116 33940 8168 33949
rect 7748 33804 7800 33856
rect 7932 33847 7984 33856
rect 7932 33813 7941 33847
rect 7941 33813 7975 33847
rect 7975 33813 7984 33847
rect 7932 33804 7984 33813
rect 8300 33847 8352 33856
rect 8300 33813 8309 33847
rect 8309 33813 8343 33847
rect 8343 33813 8352 33847
rect 8300 33804 8352 33813
rect 3010 33702 3062 33754
rect 3074 33702 3126 33754
rect 3138 33702 3190 33754
rect 3202 33702 3254 33754
rect 3266 33702 3318 33754
rect 4344 33600 4396 33652
rect 1492 33464 1544 33516
rect 7748 33507 7800 33516
rect 7748 33473 7757 33507
rect 7757 33473 7791 33507
rect 7791 33473 7800 33507
rect 7748 33464 7800 33473
rect 7840 33464 7892 33516
rect 7932 33371 7984 33380
rect 7932 33337 7941 33371
rect 7941 33337 7975 33371
rect 7975 33337 7984 33371
rect 7932 33328 7984 33337
rect 8300 33303 8352 33312
rect 8300 33269 8309 33303
rect 8309 33269 8343 33303
rect 8343 33269 8352 33303
rect 8300 33260 8352 33269
rect 1950 33158 2002 33210
rect 2014 33158 2066 33210
rect 2078 33158 2130 33210
rect 2142 33158 2194 33210
rect 2206 33158 2258 33210
rect 7950 33158 8002 33210
rect 8014 33158 8066 33210
rect 8078 33158 8130 33210
rect 8142 33158 8194 33210
rect 8206 33158 8258 33210
rect 7840 33056 7892 33108
rect 572 32852 624 32904
rect 6276 32852 6328 32904
rect 7748 32895 7800 32904
rect 7748 32861 7757 32895
rect 7757 32861 7791 32895
rect 7791 32861 7800 32895
rect 7748 32852 7800 32861
rect 3516 32784 3568 32836
rect 7840 32716 7892 32768
rect 7932 32759 7984 32768
rect 7932 32725 7941 32759
rect 7941 32725 7975 32759
rect 7975 32725 7984 32759
rect 7932 32716 7984 32725
rect 8300 32759 8352 32768
rect 8300 32725 8309 32759
rect 8309 32725 8343 32759
rect 8343 32725 8352 32759
rect 8300 32716 8352 32725
rect 3010 32614 3062 32666
rect 3074 32614 3126 32666
rect 3138 32614 3190 32666
rect 3202 32614 3254 32666
rect 3266 32614 3318 32666
rect 7748 32512 7800 32564
rect 480 32376 532 32428
rect 7748 32419 7800 32428
rect 7748 32385 7757 32419
rect 7757 32385 7791 32419
rect 7791 32385 7800 32419
rect 7748 32376 7800 32385
rect 7196 32308 7248 32360
rect 7932 32283 7984 32292
rect 7932 32249 7941 32283
rect 7941 32249 7975 32283
rect 7975 32249 7984 32283
rect 7932 32240 7984 32249
rect 8300 32215 8352 32224
rect 8300 32181 8309 32215
rect 8309 32181 8343 32215
rect 8343 32181 8352 32215
rect 8300 32172 8352 32181
rect 1950 32070 2002 32122
rect 2014 32070 2066 32122
rect 2078 32070 2130 32122
rect 2142 32070 2194 32122
rect 2206 32070 2258 32122
rect 7950 32070 8002 32122
rect 8014 32070 8066 32122
rect 8078 32070 8130 32122
rect 8142 32070 8194 32122
rect 8206 32070 8258 32122
rect 3516 31968 3568 32020
rect 8852 31900 8904 31952
rect 3516 31832 3568 31884
rect 3700 31832 3752 31884
rect 2780 31807 2832 31816
rect 2780 31773 2789 31807
rect 2789 31773 2823 31807
rect 2823 31773 2832 31807
rect 2780 31764 2832 31773
rect 4068 31764 4120 31816
rect 7472 31764 7524 31816
rect 7840 31764 7892 31816
rect 7380 31671 7432 31680
rect 7380 31637 7389 31671
rect 7389 31637 7423 31671
rect 7423 31637 7432 31671
rect 7380 31628 7432 31637
rect 8300 31671 8352 31680
rect 8300 31637 8309 31671
rect 8309 31637 8343 31671
rect 8343 31637 8352 31671
rect 8300 31628 8352 31637
rect 3010 31526 3062 31578
rect 3074 31526 3126 31578
rect 3138 31526 3190 31578
rect 3202 31526 3254 31578
rect 3266 31526 3318 31578
rect 7748 31424 7800 31476
rect 204 31288 256 31340
rect 7656 31288 7708 31340
rect 6644 31220 6696 31272
rect 7932 31195 7984 31204
rect 7932 31161 7941 31195
rect 7941 31161 7975 31195
rect 7975 31161 7984 31195
rect 7932 31152 7984 31161
rect 2780 31127 2832 31136
rect 2780 31093 2789 31127
rect 2789 31093 2823 31127
rect 2823 31093 2832 31127
rect 2780 31084 2832 31093
rect 8300 31127 8352 31136
rect 8300 31093 8309 31127
rect 8309 31093 8343 31127
rect 8343 31093 8352 31127
rect 8300 31084 8352 31093
rect 1950 30982 2002 31034
rect 2014 30982 2066 31034
rect 2078 30982 2130 31034
rect 2142 30982 2194 31034
rect 2206 30982 2258 31034
rect 7950 30982 8002 31034
rect 8014 30982 8066 31034
rect 8078 30982 8130 31034
rect 8142 30982 8194 31034
rect 8206 30982 8258 31034
rect 7012 30812 7064 30864
rect 5172 30676 5224 30728
rect 5356 30608 5408 30660
rect 7840 30540 7892 30592
rect 7932 30583 7984 30592
rect 7932 30549 7941 30583
rect 7941 30549 7975 30583
rect 7975 30549 7984 30583
rect 7932 30540 7984 30549
rect 8300 30583 8352 30592
rect 8300 30549 8309 30583
rect 8309 30549 8343 30583
rect 8343 30549 8352 30583
rect 8300 30540 8352 30549
rect 3010 30438 3062 30490
rect 3074 30438 3126 30490
rect 3138 30438 3190 30490
rect 3202 30438 3254 30490
rect 3266 30438 3318 30490
rect 112 30200 164 30252
rect 388 30132 440 30184
rect 7380 30200 7432 30252
rect 7840 30200 7892 30252
rect 9128 30132 9180 30184
rect 7472 30064 7524 30116
rect 7932 30107 7984 30116
rect 7932 30073 7941 30107
rect 7941 30073 7975 30107
rect 7975 30073 7984 30107
rect 7932 30064 7984 30073
rect 7196 29996 7248 30048
rect 7748 29996 7800 30048
rect 8300 30039 8352 30048
rect 8300 30005 8309 30039
rect 8309 30005 8343 30039
rect 8343 30005 8352 30039
rect 8300 29996 8352 30005
rect 1950 29894 2002 29946
rect 2014 29894 2066 29946
rect 2078 29894 2130 29946
rect 2142 29894 2194 29946
rect 2206 29894 2258 29946
rect 7950 29894 8002 29946
rect 8014 29894 8066 29946
rect 8078 29894 8130 29946
rect 8142 29894 8194 29946
rect 8206 29894 8258 29946
rect 9220 29656 9272 29708
rect 7748 29631 7800 29640
rect 7748 29597 7757 29631
rect 7757 29597 7791 29631
rect 7791 29597 7800 29631
rect 7748 29588 7800 29597
rect 7932 29495 7984 29504
rect 7932 29461 7941 29495
rect 7941 29461 7975 29495
rect 7975 29461 7984 29495
rect 7932 29452 7984 29461
rect 8300 29495 8352 29504
rect 8300 29461 8309 29495
rect 8309 29461 8343 29495
rect 8343 29461 8352 29495
rect 8300 29452 8352 29461
rect 3010 29350 3062 29402
rect 3074 29350 3126 29402
rect 3138 29350 3190 29402
rect 3202 29350 3254 29402
rect 3266 29350 3318 29402
rect 5724 29248 5776 29300
rect 1308 29112 1360 29164
rect 7840 29112 7892 29164
rect 9496 29044 9548 29096
rect 4804 28976 4856 29028
rect 5908 28976 5960 29028
rect 8944 28976 8996 29028
rect 8300 28951 8352 28960
rect 8300 28917 8309 28951
rect 8309 28917 8343 28951
rect 8343 28917 8352 28951
rect 8300 28908 8352 28917
rect 1950 28806 2002 28858
rect 2014 28806 2066 28858
rect 2078 28806 2130 28858
rect 2142 28806 2194 28858
rect 2206 28806 2258 28858
rect 7950 28806 8002 28858
rect 8014 28806 8066 28858
rect 8078 28806 8130 28858
rect 8142 28806 8194 28858
rect 8206 28806 8258 28858
rect 7840 28704 7892 28756
rect 8668 28568 8720 28620
rect 7288 28432 7340 28484
rect 8116 28543 8168 28552
rect 8116 28509 8125 28543
rect 8125 28509 8159 28543
rect 8159 28509 8168 28543
rect 8116 28500 8168 28509
rect 7932 28407 7984 28416
rect 7932 28373 7941 28407
rect 7941 28373 7975 28407
rect 7975 28373 7984 28407
rect 7932 28364 7984 28373
rect 8300 28407 8352 28416
rect 8300 28373 8309 28407
rect 8309 28373 8343 28407
rect 8343 28373 8352 28407
rect 8300 28364 8352 28373
rect 3010 28262 3062 28314
rect 3074 28262 3126 28314
rect 3138 28262 3190 28314
rect 3202 28262 3254 28314
rect 3266 28262 3318 28314
rect 8116 28160 8168 28212
rect 7748 28067 7800 28076
rect 7748 28033 7757 28067
rect 7757 28033 7791 28067
rect 7791 28033 7800 28067
rect 7748 28024 7800 28033
rect 7840 28024 7892 28076
rect 8944 27956 8996 28008
rect 7932 27931 7984 27940
rect 7932 27897 7941 27931
rect 7941 27897 7975 27931
rect 7975 27897 7984 27931
rect 7932 27888 7984 27897
rect 8300 27863 8352 27872
rect 8300 27829 8309 27863
rect 8309 27829 8343 27863
rect 8343 27829 8352 27863
rect 8300 27820 8352 27829
rect 1950 27718 2002 27770
rect 2014 27718 2066 27770
rect 2078 27718 2130 27770
rect 2142 27718 2194 27770
rect 2206 27718 2258 27770
rect 7950 27718 8002 27770
rect 8014 27718 8066 27770
rect 8078 27718 8130 27770
rect 8142 27718 8194 27770
rect 8206 27718 8258 27770
rect 7748 27616 7800 27668
rect 3976 27548 4028 27600
rect 1216 27412 1268 27464
rect 6736 27412 6788 27464
rect 7564 27412 7616 27464
rect 7196 27344 7248 27396
rect 7932 27319 7984 27328
rect 7932 27285 7941 27319
rect 7941 27285 7975 27319
rect 7975 27285 7984 27319
rect 7932 27276 7984 27285
rect 8300 27319 8352 27328
rect 8300 27285 8309 27319
rect 8309 27285 8343 27319
rect 8343 27285 8352 27319
rect 8300 27276 8352 27285
rect 3010 27174 3062 27226
rect 3074 27174 3126 27226
rect 3138 27174 3190 27226
rect 3202 27174 3254 27226
rect 3266 27174 3318 27226
rect 7840 27072 7892 27124
rect 7380 26936 7432 26988
rect 7748 26979 7800 26988
rect 7748 26945 7757 26979
rect 7757 26945 7791 26979
rect 7791 26945 7800 26979
rect 7748 26936 7800 26945
rect 7472 26868 7524 26920
rect 7932 26843 7984 26852
rect 7932 26809 7941 26843
rect 7941 26809 7975 26843
rect 7975 26809 7984 26843
rect 7932 26800 7984 26809
rect 8300 26775 8352 26784
rect 8300 26741 8309 26775
rect 8309 26741 8343 26775
rect 8343 26741 8352 26775
rect 8300 26732 8352 26741
rect 1950 26630 2002 26682
rect 2014 26630 2066 26682
rect 2078 26630 2130 26682
rect 2142 26630 2194 26682
rect 2206 26630 2258 26682
rect 7950 26630 8002 26682
rect 8014 26630 8066 26682
rect 8078 26630 8130 26682
rect 8142 26630 8194 26682
rect 8206 26630 8258 26682
rect 7564 26528 7616 26580
rect 7380 26503 7432 26512
rect 7380 26469 7389 26503
rect 7389 26469 7423 26503
rect 7423 26469 7432 26503
rect 7380 26460 7432 26469
rect 8760 26460 8812 26512
rect 8576 26392 8628 26444
rect 8024 26367 8076 26376
rect 8024 26333 8033 26367
rect 8033 26333 8067 26367
rect 8067 26333 8076 26367
rect 8024 26324 8076 26333
rect 2872 26256 2924 26308
rect 7380 26256 7432 26308
rect 8300 26231 8352 26240
rect 8300 26197 8309 26231
rect 8309 26197 8343 26231
rect 8343 26197 8352 26231
rect 8300 26188 8352 26197
rect 3010 26086 3062 26138
rect 3074 26086 3126 26138
rect 3138 26086 3190 26138
rect 3202 26086 3254 26138
rect 3266 26086 3318 26138
rect 2688 25984 2740 26036
rect 5448 25984 5500 26036
rect 7196 26027 7248 26036
rect 7196 25993 7205 26027
rect 7205 25993 7239 26027
rect 7239 25993 7248 26027
rect 7196 25984 7248 25993
rect 2504 25848 2556 25900
rect 3056 25848 3108 25900
rect 8484 25916 8536 25968
rect 7564 25848 7616 25900
rect 6552 25780 6604 25832
rect 7932 25755 7984 25764
rect 7932 25721 7941 25755
rect 7941 25721 7975 25755
rect 7975 25721 7984 25755
rect 7932 25712 7984 25721
rect 8300 25687 8352 25696
rect 8300 25653 8309 25687
rect 8309 25653 8343 25687
rect 8343 25653 8352 25687
rect 8300 25644 8352 25653
rect 1950 25542 2002 25594
rect 2014 25542 2066 25594
rect 2078 25542 2130 25594
rect 2142 25542 2194 25594
rect 2206 25542 2258 25594
rect 7950 25542 8002 25594
rect 8014 25542 8066 25594
rect 8078 25542 8130 25594
rect 8142 25542 8194 25594
rect 8206 25542 8258 25594
rect 1860 25483 1912 25492
rect 1860 25449 1869 25483
rect 1869 25449 1903 25483
rect 1903 25449 1912 25483
rect 1860 25440 1912 25449
rect 7748 25440 7800 25492
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 9312 25304 9364 25356
rect 7748 25279 7800 25288
rect 7748 25245 7757 25279
rect 7757 25245 7791 25279
rect 7791 25245 7800 25279
rect 7748 25236 7800 25245
rect 3056 25211 3108 25220
rect 3056 25177 3065 25211
rect 3065 25177 3099 25211
rect 3099 25177 3108 25211
rect 3056 25168 3108 25177
rect 6460 25168 6512 25220
rect 7932 25143 7984 25152
rect 7932 25109 7941 25143
rect 7941 25109 7975 25143
rect 7975 25109 7984 25143
rect 7932 25100 7984 25109
rect 8300 25143 8352 25152
rect 8300 25109 8309 25143
rect 8309 25109 8343 25143
rect 8343 25109 8352 25143
rect 8300 25100 8352 25109
rect 3010 24998 3062 25050
rect 3074 24998 3126 25050
rect 3138 24998 3190 25050
rect 3202 24998 3254 25050
rect 3266 24998 3318 25050
rect 2412 24828 2464 24880
rect 6368 24828 6420 24880
rect 7012 24803 7064 24812
rect 7012 24769 7021 24803
rect 7021 24769 7055 24803
rect 7055 24769 7064 24803
rect 7012 24760 7064 24769
rect 7104 24624 7156 24676
rect 7472 24667 7524 24676
rect 7472 24633 7481 24667
rect 7481 24633 7515 24667
rect 7515 24633 7524 24667
rect 7472 24624 7524 24633
rect 7840 24760 7892 24812
rect 7656 24692 7708 24744
rect 9588 24624 9640 24676
rect 7840 24556 7892 24608
rect 9036 24556 9088 24608
rect 1950 24454 2002 24506
rect 2014 24454 2066 24506
rect 2078 24454 2130 24506
rect 2142 24454 2194 24506
rect 2206 24454 2258 24506
rect 7950 24454 8002 24506
rect 8014 24454 8066 24506
rect 8078 24454 8130 24506
rect 8142 24454 8194 24506
rect 8206 24454 8258 24506
rect 3424 24395 3476 24404
rect 3424 24361 3433 24395
rect 3433 24361 3467 24395
rect 3467 24361 3476 24395
rect 3424 24352 3476 24361
rect 5080 24395 5132 24404
rect 5080 24361 5089 24395
rect 5089 24361 5123 24395
rect 5123 24361 5132 24395
rect 5080 24352 5132 24361
rect 7196 24352 7248 24404
rect 7472 24352 7524 24404
rect 7656 24395 7708 24404
rect 7656 24361 7665 24395
rect 7665 24361 7699 24395
rect 7699 24361 7708 24395
rect 7656 24352 7708 24361
rect 3700 24284 3752 24336
rect 3424 24216 3476 24268
rect 3700 24148 3752 24200
rect 4988 24148 5040 24200
rect 9404 24216 9456 24268
rect 7012 24123 7064 24132
rect 7012 24089 7021 24123
rect 7021 24089 7055 24123
rect 7055 24089 7064 24123
rect 7012 24080 7064 24089
rect 7104 24080 7156 24132
rect 6368 24012 6420 24064
rect 7932 24055 7984 24064
rect 7932 24021 7941 24055
rect 7941 24021 7975 24055
rect 7975 24021 7984 24055
rect 7932 24012 7984 24021
rect 8300 24055 8352 24064
rect 8300 24021 8309 24055
rect 8309 24021 8343 24055
rect 8343 24021 8352 24055
rect 8300 24012 8352 24021
rect 3010 23910 3062 23962
rect 3074 23910 3126 23962
rect 3138 23910 3190 23962
rect 3202 23910 3254 23962
rect 3266 23910 3318 23962
rect 1584 23808 1636 23860
rect 7012 23808 7064 23860
rect 7196 23808 7248 23860
rect 1400 23672 1452 23724
rect 5264 23672 5316 23724
rect 7840 23672 7892 23724
rect 1032 23536 1084 23588
rect 6276 23536 6328 23588
rect 8852 23536 8904 23588
rect 4988 23511 5040 23520
rect 4988 23477 4997 23511
rect 4997 23477 5031 23511
rect 5031 23477 5040 23511
rect 4988 23468 5040 23477
rect 9036 23468 9088 23520
rect 1950 23366 2002 23418
rect 2014 23366 2066 23418
rect 2078 23366 2130 23418
rect 2142 23366 2194 23418
rect 2206 23366 2258 23418
rect 7950 23366 8002 23418
rect 8014 23366 8066 23418
rect 8078 23366 8130 23418
rect 8142 23366 8194 23418
rect 8206 23366 8258 23418
rect 7840 23264 7892 23316
rect 7656 23060 7708 23112
rect 7196 22992 7248 23044
rect 8116 23103 8168 23112
rect 8116 23069 8125 23103
rect 8125 23069 8159 23103
rect 8159 23069 8168 23103
rect 8116 23060 8168 23069
rect 7932 22967 7984 22976
rect 7932 22933 7941 22967
rect 7941 22933 7975 22967
rect 7975 22933 7984 22967
rect 7932 22924 7984 22933
rect 8300 22967 8352 22976
rect 8300 22933 8309 22967
rect 8309 22933 8343 22967
rect 8343 22933 8352 22967
rect 8300 22924 8352 22933
rect 3010 22822 3062 22874
rect 3074 22822 3126 22874
rect 3138 22822 3190 22874
rect 3202 22822 3254 22874
rect 3266 22822 3318 22874
rect 3792 22763 3844 22772
rect 3792 22729 3801 22763
rect 3801 22729 3835 22763
rect 3835 22729 3844 22763
rect 3792 22720 3844 22729
rect 6920 22720 6972 22772
rect 7656 22720 7708 22772
rect 2688 22652 2740 22704
rect 940 22584 992 22636
rect 3976 22584 4028 22636
rect 7656 22584 7708 22636
rect 5816 22516 5868 22568
rect 6184 22448 6236 22500
rect 7012 22448 7064 22500
rect 7288 22448 7340 22500
rect 7840 22380 7892 22432
rect 9036 22380 9088 22432
rect 1950 22278 2002 22330
rect 2014 22278 2066 22330
rect 2078 22278 2130 22330
rect 2142 22278 2194 22330
rect 2206 22278 2258 22330
rect 7950 22278 8002 22330
rect 8014 22278 8066 22330
rect 8078 22278 8130 22330
rect 8142 22278 8194 22330
rect 8206 22278 8258 22330
rect 6184 22176 6236 22228
rect 6460 22176 6512 22228
rect 7380 22176 7432 22228
rect 8392 22176 8444 22228
rect 7656 22108 7708 22160
rect 8208 22108 8260 22160
rect 4528 22015 4580 22024
rect 4528 21981 4537 22015
rect 4537 21981 4571 22015
rect 4571 21981 4580 22015
rect 4528 21972 4580 21981
rect 6552 21972 6604 22024
rect 6736 22015 6788 22024
rect 6736 21981 6745 22015
rect 6745 21981 6779 22015
rect 6779 21981 6788 22015
rect 6736 21972 6788 21981
rect 7380 21972 7432 22024
rect 8024 21972 8076 22024
rect 5908 21904 5960 21956
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 6828 21836 6880 21888
rect 7932 21879 7984 21888
rect 7932 21845 7941 21879
rect 7941 21845 7975 21879
rect 7975 21845 7984 21879
rect 7932 21836 7984 21845
rect 8300 21879 8352 21888
rect 8300 21845 8309 21879
rect 8309 21845 8343 21879
rect 8343 21845 8352 21879
rect 8300 21836 8352 21845
rect 3010 21734 3062 21786
rect 3074 21734 3126 21786
rect 3138 21734 3190 21786
rect 3202 21734 3254 21786
rect 3266 21734 3318 21786
rect 3516 21632 3568 21684
rect 7380 21675 7432 21684
rect 7380 21641 7389 21675
rect 7389 21641 7423 21675
rect 7423 21641 7432 21675
rect 7380 21632 7432 21641
rect 756 21496 808 21548
rect 3792 21428 3844 21480
rect 7380 21428 7432 21480
rect 3976 21292 4028 21344
rect 5448 21292 5500 21344
rect 7840 21292 7892 21344
rect 9036 21292 9088 21344
rect 1950 21190 2002 21242
rect 2014 21190 2066 21242
rect 2078 21190 2130 21242
rect 2142 21190 2194 21242
rect 2206 21190 2258 21242
rect 7950 21190 8002 21242
rect 8014 21190 8066 21242
rect 8078 21190 8130 21242
rect 8142 21190 8194 21242
rect 8206 21190 8258 21242
rect 6920 21131 6972 21140
rect 6920 21097 6929 21131
rect 6929 21097 6963 21131
rect 6963 21097 6972 21131
rect 6920 21088 6972 21097
rect 8852 21020 8904 21072
rect 296 20884 348 20936
rect 1676 20884 1728 20936
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 7748 20927 7800 20936
rect 7748 20893 7757 20927
rect 7757 20893 7791 20927
rect 7791 20893 7800 20927
rect 7748 20884 7800 20893
rect 8116 20927 8168 20936
rect 8116 20893 8125 20927
rect 8125 20893 8159 20927
rect 8159 20893 8168 20927
rect 8116 20884 8168 20893
rect 6552 20748 6604 20800
rect 6828 20748 6880 20800
rect 8300 20791 8352 20800
rect 8300 20757 8309 20791
rect 8309 20757 8343 20791
rect 8343 20757 8352 20791
rect 8300 20748 8352 20757
rect 3010 20646 3062 20698
rect 3074 20646 3126 20698
rect 3138 20646 3190 20698
rect 3202 20646 3254 20698
rect 3266 20646 3318 20698
rect 5264 20587 5316 20596
rect 5264 20553 5273 20587
rect 5273 20553 5307 20587
rect 5307 20553 5316 20587
rect 5264 20544 5316 20553
rect 5540 20587 5592 20596
rect 5540 20553 5549 20587
rect 5549 20553 5583 20587
rect 5583 20553 5592 20587
rect 5540 20544 5592 20553
rect 5080 20451 5132 20460
rect 5080 20417 5089 20451
rect 5089 20417 5123 20451
rect 5123 20417 5132 20451
rect 5080 20408 5132 20417
rect 5356 20451 5408 20460
rect 5356 20417 5365 20451
rect 5365 20417 5399 20451
rect 5399 20417 5408 20451
rect 5356 20408 5408 20417
rect 7748 20451 7800 20460
rect 7748 20417 7757 20451
rect 7757 20417 7791 20451
rect 7791 20417 7800 20451
rect 7748 20408 7800 20417
rect 8116 20451 8168 20460
rect 8116 20417 8125 20451
rect 8125 20417 8159 20451
rect 8159 20417 8168 20451
rect 8116 20408 8168 20417
rect 7840 20204 7892 20256
rect 9036 20204 9088 20256
rect 1950 20102 2002 20154
rect 2014 20102 2066 20154
rect 2078 20102 2130 20154
rect 2142 20102 2194 20154
rect 2206 20102 2258 20154
rect 7950 20102 8002 20154
rect 8014 20102 8066 20154
rect 8078 20102 8130 20154
rect 8142 20102 8194 20154
rect 8206 20102 8258 20154
rect 2596 20043 2648 20052
rect 2596 20009 2605 20043
rect 2605 20009 2639 20043
rect 2639 20009 2648 20043
rect 2596 20000 2648 20009
rect 4896 20043 4948 20052
rect 4896 20009 4905 20043
rect 4905 20009 4939 20043
rect 4939 20009 4948 20043
rect 4896 20000 4948 20009
rect 6920 20000 6972 20052
rect 7196 20000 7248 20052
rect 7564 20000 7616 20052
rect 7932 20000 7984 20052
rect 7196 19864 7248 19916
rect 1676 19796 1728 19848
rect 4436 19796 4488 19848
rect 5908 19796 5960 19848
rect 3884 19660 3936 19712
rect 7564 19660 7616 19712
rect 7932 19703 7984 19712
rect 7932 19669 7941 19703
rect 7941 19669 7975 19703
rect 7975 19669 7984 19703
rect 7932 19660 7984 19669
rect 8300 19703 8352 19712
rect 8300 19669 8309 19703
rect 8309 19669 8343 19703
rect 8343 19669 8352 19703
rect 8300 19660 8352 19669
rect 3010 19558 3062 19610
rect 3074 19558 3126 19610
rect 3138 19558 3190 19610
rect 3202 19558 3254 19610
rect 3266 19558 3318 19610
rect 3424 19456 3476 19508
rect 3516 19499 3568 19508
rect 3516 19465 3525 19499
rect 3525 19465 3559 19499
rect 3559 19465 3568 19499
rect 3516 19456 3568 19465
rect 3608 19499 3660 19508
rect 3608 19465 3617 19499
rect 3617 19465 3651 19499
rect 3651 19465 3660 19499
rect 3608 19456 3660 19465
rect 6644 19499 6696 19508
rect 6644 19465 6653 19499
rect 6653 19465 6687 19499
rect 6687 19465 6696 19499
rect 6644 19456 6696 19465
rect 7472 19456 7524 19508
rect 5264 19388 5316 19440
rect 9036 19456 9088 19508
rect 1124 19320 1176 19372
rect 3424 19320 3476 19372
rect 3516 19320 3568 19372
rect 6460 19363 6512 19372
rect 6460 19329 6469 19363
rect 6469 19329 6503 19363
rect 6503 19329 6512 19363
rect 6460 19320 6512 19329
rect 7564 19320 7616 19372
rect 8760 19388 8812 19440
rect 8392 19252 8444 19304
rect 7472 19184 7524 19236
rect 8208 19184 8260 19236
rect 1950 19014 2002 19066
rect 2014 19014 2066 19066
rect 2078 19014 2130 19066
rect 2142 19014 2194 19066
rect 2206 19014 2258 19066
rect 7950 19014 8002 19066
rect 8014 19014 8066 19066
rect 8078 19014 8130 19066
rect 8142 19014 8194 19066
rect 8206 19014 8258 19066
rect 7288 18955 7340 18964
rect 7288 18921 7297 18955
rect 7297 18921 7331 18955
rect 7331 18921 7340 18955
rect 7288 18912 7340 18921
rect 7380 18912 7432 18964
rect 6276 18844 6328 18896
rect 7288 18708 7340 18760
rect 6092 18572 6144 18624
rect 9680 18640 9732 18692
rect 7932 18615 7984 18624
rect 7932 18581 7941 18615
rect 7941 18581 7975 18615
rect 7975 18581 7984 18615
rect 7932 18572 7984 18581
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 3010 18470 3062 18522
rect 3074 18470 3126 18522
rect 3138 18470 3190 18522
rect 3202 18470 3254 18522
rect 3266 18470 3318 18522
rect 4804 18411 4856 18420
rect 4804 18377 4813 18411
rect 4813 18377 4847 18411
rect 4847 18377 4856 18411
rect 4804 18368 4856 18377
rect 7104 18368 7156 18420
rect 7288 18300 7340 18352
rect 9036 18300 9088 18352
rect 4620 18275 4672 18284
rect 4620 18241 4629 18275
rect 4629 18241 4663 18275
rect 4663 18241 4672 18275
rect 4620 18232 4672 18241
rect 8760 18232 8812 18284
rect 1950 17926 2002 17978
rect 2014 17926 2066 17978
rect 2078 17926 2130 17978
rect 2142 17926 2194 17978
rect 2206 17926 2258 17978
rect 7950 17926 8002 17978
rect 8014 17926 8066 17978
rect 8078 17926 8130 17978
rect 8142 17926 8194 17978
rect 8206 17926 8258 17978
rect 1768 17867 1820 17876
rect 1768 17833 1777 17867
rect 1777 17833 1811 17867
rect 1811 17833 1820 17867
rect 1768 17824 1820 17833
rect 6368 17824 6420 17876
rect 6184 17688 6236 17740
rect 6368 17688 6420 17740
rect 848 17620 900 17672
rect 7656 17620 7708 17672
rect 3010 17382 3062 17434
rect 3074 17382 3126 17434
rect 3138 17382 3190 17434
rect 3202 17382 3254 17434
rect 3266 17382 3318 17434
rect 7012 17280 7064 17332
rect 6920 17008 6972 17060
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 7950 16838 8002 16890
rect 8014 16838 8066 16890
rect 8078 16838 8130 16890
rect 8142 16838 8194 16890
rect 8206 16838 8258 16890
rect 3010 16294 3062 16346
rect 3074 16294 3126 16346
rect 3138 16294 3190 16346
rect 3202 16294 3254 16346
rect 3266 16294 3318 16346
rect 1860 16235 1912 16244
rect 1860 16201 1869 16235
rect 1869 16201 1903 16235
rect 1903 16201 1912 16235
rect 1860 16192 1912 16201
rect 4896 16235 4948 16244
rect 4896 16201 4905 16235
rect 4905 16201 4939 16235
rect 4939 16201 4948 16235
rect 4896 16192 4948 16201
rect 6368 16192 6420 16244
rect 7564 16235 7616 16244
rect 7564 16201 7573 16235
rect 7573 16201 7607 16235
rect 7607 16201 7616 16235
rect 7564 16192 7616 16201
rect 1216 16056 1268 16108
rect 4896 16056 4948 16108
rect 8760 16056 8812 16108
rect 8576 15988 8628 16040
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 7950 15750 8002 15802
rect 8014 15750 8066 15802
rect 8078 15750 8130 15802
rect 8142 15750 8194 15802
rect 8206 15750 8258 15802
rect 2320 15648 2372 15700
rect 756 15444 808 15496
rect 3010 15206 3062 15258
rect 3074 15206 3126 15258
rect 3138 15206 3190 15258
rect 3202 15206 3254 15258
rect 3266 15206 3318 15258
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 8484 14968 8536 15020
rect 6920 14764 6972 14816
rect 7932 14764 7984 14816
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 7950 14662 8002 14714
rect 8014 14662 8066 14714
rect 8078 14662 8130 14714
rect 8142 14662 8194 14714
rect 8206 14662 8258 14714
rect 2412 14560 2464 14612
rect 6920 14603 6972 14612
rect 6920 14569 6929 14603
rect 6929 14569 6963 14603
rect 6963 14569 6972 14603
rect 6920 14560 6972 14569
rect 7472 14560 7524 14612
rect 1032 14356 1084 14408
rect 9496 14356 9548 14408
rect 8300 14288 8352 14340
rect 3010 14118 3062 14170
rect 3074 14118 3126 14170
rect 3138 14118 3190 14170
rect 3202 14118 3254 14170
rect 3266 14118 3318 14170
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 7950 13574 8002 13626
rect 8014 13574 8066 13626
rect 8078 13574 8130 13626
rect 8142 13574 8194 13626
rect 8206 13574 8258 13626
rect 1860 13515 1912 13524
rect 1860 13481 1869 13515
rect 1869 13481 1903 13515
rect 1903 13481 1912 13515
rect 1860 13472 1912 13481
rect 7840 13472 7892 13524
rect 756 13268 808 13320
rect 8760 13268 8812 13320
rect 3010 13030 3062 13082
rect 3074 13030 3126 13082
rect 3138 13030 3190 13082
rect 3202 13030 3254 13082
rect 3266 13030 3318 13082
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 7950 12486 8002 12538
rect 8014 12486 8066 12538
rect 8078 12486 8130 12538
rect 8142 12486 8194 12538
rect 8206 12486 8258 12538
rect 2688 12384 2740 12436
rect 6828 12384 6880 12436
rect 8760 12180 8812 12232
rect 8484 12112 8536 12164
rect 3010 11942 3062 11994
rect 3074 11942 3126 11994
rect 3138 11942 3190 11994
rect 3202 11942 3254 11994
rect 3266 11942 3318 11994
rect 8392 11840 8444 11892
rect 8944 11704 8996 11756
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 7950 11398 8002 11450
rect 8014 11398 8066 11450
rect 8078 11398 8130 11450
rect 8142 11398 8194 11450
rect 8206 11398 8258 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 5816 11339 5868 11348
rect 5816 11305 5825 11339
rect 5825 11305 5859 11339
rect 5859 11305 5868 11339
rect 5816 11296 5868 11305
rect 1124 11092 1176 11144
rect 8300 11092 8352 11144
rect 3010 10854 3062 10906
rect 3074 10854 3126 10906
rect 3138 10854 3190 10906
rect 3202 10854 3254 10906
rect 3266 10854 3318 10906
rect 7012 10752 7064 10804
rect 8392 10616 8444 10668
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 7950 10310 8002 10362
rect 8014 10310 8066 10362
rect 8078 10310 8130 10362
rect 8142 10310 8194 10362
rect 8206 10310 8258 10362
rect 3010 9766 3062 9818
rect 3074 9766 3126 9818
rect 3138 9766 3190 9818
rect 3202 9766 3254 9818
rect 3266 9766 3318 9818
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7104 9435 7156 9444
rect 7104 9401 7113 9435
rect 7113 9401 7147 9435
rect 7147 9401 7156 9435
rect 7104 9392 7156 9401
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 7950 9222 8002 9274
rect 8014 9222 8066 9274
rect 8078 9222 8130 9274
rect 8142 9222 8194 9274
rect 8206 9222 8258 9274
rect 5172 9120 5224 9172
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 5908 8576 5960 8628
rect 8392 8440 8444 8492
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 7840 6740 7892 6792
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 7380 6443 7432 6452
rect 7380 6409 7389 6443
rect 7389 6409 7423 6443
rect 7423 6409 7432 6443
rect 7380 6400 7432 6409
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 6000 5899 6052 5908
rect 6000 5865 6009 5899
rect 6009 5865 6043 5899
rect 6043 5865 6052 5899
rect 6000 5856 6052 5865
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 6184 4811 6236 4820
rect 6184 4777 6193 4811
rect 6193 4777 6227 4811
rect 6227 4777 6236 4811
rect 6184 4768 6236 4777
rect 6736 4564 6788 4616
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 3792 3952 3844 4004
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 3884 3680 3936 3732
rect 7840 3476 7892 3528
rect 3424 3408 3476 3460
rect 6736 3408 6788 3460
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 6092 3179 6144 3188
rect 6092 3145 6101 3179
rect 6101 3145 6135 3179
rect 6135 3145 6144 3179
rect 6092 3136 6144 3145
rect 6276 3136 6328 3188
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 7748 3000 7800 3052
rect 5264 2864 5316 2916
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 2136 2592 2188 2644
rect 2688 2592 2740 2644
rect 5448 2592 5500 2644
rect 8576 2592 8628 2644
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 1676 2048 1728 2100
rect 2596 2048 2648 2100
rect 4528 416 4580 468
rect 6276 416 6328 468
<< metal2 >>
rect 294 44960 350 45016
rect 754 44960 810 45016
rect 1214 44960 1270 45016
rect 1674 44960 1730 45016
rect 2134 44960 2190 45016
rect 2594 44960 2650 45016
rect 2884 44974 3004 45002
rect 308 41818 336 44960
rect 296 41812 348 41818
rect 296 41754 348 41760
rect 768 41750 796 44960
rect 1228 42362 1256 44960
rect 1688 42362 1716 44960
rect 2148 42362 2176 44960
rect 2608 42362 2636 44960
rect 2884 42362 2912 44974
rect 2976 44962 3004 44974
rect 3054 44962 3110 45016
rect 2976 44960 3110 44962
rect 3514 44960 3570 45016
rect 3974 44960 4030 45016
rect 4434 44960 4490 45016
rect 4894 44960 4950 45016
rect 5354 44960 5410 45016
rect 5814 44960 5870 45016
rect 6274 44960 6330 45016
rect 6734 44960 6790 45016
rect 7194 44960 7250 45016
rect 7654 44960 7710 45016
rect 8114 44960 8170 45016
rect 8574 44960 8630 45016
rect 9034 44960 9090 45016
rect 9494 44960 9550 45016
rect 2976 44934 3096 44960
rect 3010 42460 3318 42469
rect 3010 42458 3016 42460
rect 3072 42458 3096 42460
rect 3152 42458 3176 42460
rect 3232 42458 3256 42460
rect 3312 42458 3318 42460
rect 3072 42406 3074 42458
rect 3254 42406 3256 42458
rect 3010 42404 3016 42406
rect 3072 42404 3096 42406
rect 3152 42404 3176 42406
rect 3232 42404 3256 42406
rect 3312 42404 3318 42406
rect 3010 42395 3318 42404
rect 3528 42362 3556 44960
rect 3988 42362 4016 44960
rect 4448 42362 4476 44960
rect 4908 42362 4936 44960
rect 5368 42362 5396 44960
rect 5828 42362 5856 44960
rect 6288 42362 6316 44960
rect 6748 42362 6776 44960
rect 7208 42362 7236 44960
rect 7378 43616 7434 43625
rect 7378 43551 7434 43560
rect 1216 42356 1268 42362
rect 1216 42298 1268 42304
rect 1676 42356 1728 42362
rect 1676 42298 1728 42304
rect 2136 42356 2188 42362
rect 2136 42298 2188 42304
rect 2596 42356 2648 42362
rect 2596 42298 2648 42304
rect 2872 42356 2924 42362
rect 2872 42298 2924 42304
rect 3516 42356 3568 42362
rect 3516 42298 3568 42304
rect 3976 42356 4028 42362
rect 3976 42298 4028 42304
rect 4436 42356 4488 42362
rect 4436 42298 4488 42304
rect 4896 42356 4948 42362
rect 4896 42298 4948 42304
rect 5356 42356 5408 42362
rect 5356 42298 5408 42304
rect 5816 42356 5868 42362
rect 5816 42298 5868 42304
rect 6276 42356 6328 42362
rect 6276 42298 6328 42304
rect 6736 42356 6788 42362
rect 6736 42298 6788 42304
rect 7196 42356 7248 42362
rect 7196 42298 7248 42304
rect 4528 42288 4580 42294
rect 4528 42230 4580 42236
rect 1676 42220 1728 42226
rect 1676 42162 1728 42168
rect 2596 42220 2648 42226
rect 2596 42162 2648 42168
rect 3424 42220 3476 42226
rect 3424 42162 3476 42168
rect 3608 42220 3660 42226
rect 3608 42162 3660 42168
rect 3792 42220 3844 42226
rect 3792 42162 3844 42168
rect 1584 42152 1636 42158
rect 1584 42094 1636 42100
rect 756 41744 808 41750
rect 756 41686 808 41692
rect 204 40520 256 40526
rect 204 40462 256 40468
rect 112 39432 164 39438
rect 112 39374 164 39380
rect 124 31385 152 39374
rect 216 34105 244 40462
rect 1308 38344 1360 38350
rect 1308 38286 1360 38292
rect 848 36168 900 36174
rect 848 36110 900 36116
rect 296 35080 348 35086
rect 296 35022 348 35028
rect 202 34096 258 34105
rect 202 34031 258 34040
rect 110 31376 166 31385
rect 110 31311 166 31320
rect 204 31340 256 31346
rect 204 31282 256 31288
rect 112 30252 164 30258
rect 112 30194 164 30200
rect 124 2825 152 30194
rect 216 5545 244 31282
rect 308 23225 336 35022
rect 664 33992 716 33998
rect 664 33934 716 33940
rect 572 32904 624 32910
rect 572 32846 624 32852
rect 480 32428 532 32434
rect 480 32370 532 32376
rect 388 30184 440 30190
rect 388 30126 440 30132
rect 294 23216 350 23225
rect 294 23151 350 23160
rect 296 20936 348 20942
rect 296 20878 348 20884
rect 202 5536 258 5545
rect 202 5471 258 5480
rect 110 2816 166 2825
rect 110 2751 166 2760
rect 308 56 336 20878
rect 400 4185 428 30126
rect 492 8265 520 32370
rect 584 9625 612 32846
rect 676 16130 704 33934
rect 860 24585 888 36110
rect 1320 30025 1348 38286
rect 1492 33516 1544 33522
rect 1492 33458 1544 33464
rect 1306 30016 1362 30025
rect 1306 29951 1362 29960
rect 1308 29164 1360 29170
rect 1308 29106 1360 29112
rect 1320 28665 1348 29106
rect 1306 28656 1362 28665
rect 1306 28591 1362 28600
rect 1216 27464 1268 27470
rect 1216 27406 1268 27412
rect 1228 25945 1256 27406
rect 1214 25936 1270 25945
rect 1214 25871 1270 25880
rect 846 24576 902 24585
rect 846 24511 902 24520
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1032 23588 1084 23594
rect 1032 23530 1084 23536
rect 940 22636 992 22642
rect 940 22578 992 22584
rect 756 21548 808 21554
rect 756 21490 808 21496
rect 768 19145 796 21490
rect 952 20505 980 22578
rect 938 20496 994 20505
rect 938 20431 994 20440
rect 754 19136 810 19145
rect 754 19071 810 19080
rect 1044 18850 1072 23530
rect 1124 19372 1176 19378
rect 1124 19314 1176 19320
rect 768 18822 1072 18850
rect 768 16266 796 18822
rect 1136 17785 1164 19314
rect 1122 17776 1178 17785
rect 1122 17711 1178 17720
rect 848 17672 900 17678
rect 848 17614 900 17620
rect 860 16425 888 17614
rect 846 16416 902 16425
rect 846 16351 902 16360
rect 768 16238 1164 16266
rect 676 16102 980 16130
rect 756 15496 808 15502
rect 756 15438 808 15444
rect 768 15065 796 15438
rect 754 15056 810 15065
rect 754 14991 810 15000
rect 756 13320 808 13326
rect 756 13262 808 13268
rect 768 12345 796 13262
rect 754 12336 810 12345
rect 754 12271 810 12280
rect 952 10985 980 16102
rect 1032 14408 1084 14414
rect 1032 14350 1084 14356
rect 1044 13705 1072 14350
rect 1030 13696 1086 13705
rect 1030 13631 1086 13640
rect 1136 12434 1164 16238
rect 1216 16108 1268 16114
rect 1216 16050 1268 16056
rect 1044 12406 1164 12434
rect 938 10976 994 10985
rect 938 10911 994 10920
rect 570 9616 626 9625
rect 570 9551 626 9560
rect 478 8256 534 8265
rect 478 8191 534 8200
rect 1044 7562 1072 12406
rect 1124 11144 1176 11150
rect 1124 11086 1176 11092
rect 676 7534 1072 7562
rect 386 4176 442 4185
rect 386 4111 442 4120
rect 676 1465 704 7534
rect 1136 2774 1164 11086
rect 768 2746 1164 2774
rect 662 1456 718 1465
rect 662 1391 718 1400
rect 768 56 796 2746
rect 1228 56 1256 16050
rect 294 0 350 56
rect 754 0 810 56
rect 1214 0 1270 56
rect 1412 42 1440 23666
rect 1504 21865 1532 33458
rect 1596 23866 1624 42094
rect 1688 41721 1716 42162
rect 1950 41916 2258 41925
rect 1950 41914 1956 41916
rect 2012 41914 2036 41916
rect 2092 41914 2116 41916
rect 2172 41914 2196 41916
rect 2252 41914 2258 41916
rect 2012 41862 2014 41914
rect 2194 41862 2196 41914
rect 1950 41860 1956 41862
rect 2012 41860 2036 41862
rect 2092 41860 2116 41862
rect 2172 41860 2196 41862
rect 2252 41860 2258 41862
rect 1950 41851 2258 41860
rect 1674 41712 1730 41721
rect 1674 41647 1730 41656
rect 1676 41608 1728 41614
rect 1676 41550 1728 41556
rect 1860 41608 1912 41614
rect 1860 41550 1912 41556
rect 1688 41449 1716 41550
rect 1674 41440 1730 41449
rect 1674 41375 1730 41384
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1490 21856 1546 21865
rect 1490 21791 1546 21800
rect 1688 20942 1716 25230
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1688 2106 1716 19790
rect 1780 17882 1808 34546
rect 1872 25498 1900 41550
rect 1950 40828 2258 40837
rect 1950 40826 1956 40828
rect 2012 40826 2036 40828
rect 2092 40826 2116 40828
rect 2172 40826 2196 40828
rect 2252 40826 2258 40828
rect 2012 40774 2014 40826
rect 2194 40774 2196 40826
rect 1950 40772 1956 40774
rect 2012 40772 2036 40774
rect 2092 40772 2116 40774
rect 2172 40772 2196 40774
rect 2252 40772 2258 40774
rect 1950 40763 2258 40772
rect 1950 39740 2258 39749
rect 1950 39738 1956 39740
rect 2012 39738 2036 39740
rect 2092 39738 2116 39740
rect 2172 39738 2196 39740
rect 2252 39738 2258 39740
rect 2012 39686 2014 39738
rect 2194 39686 2196 39738
rect 1950 39684 1956 39686
rect 2012 39684 2036 39686
rect 2092 39684 2116 39686
rect 2172 39684 2196 39686
rect 2252 39684 2258 39686
rect 1950 39675 2258 39684
rect 1950 38652 2258 38661
rect 1950 38650 1956 38652
rect 2012 38650 2036 38652
rect 2092 38650 2116 38652
rect 2172 38650 2196 38652
rect 2252 38650 2258 38652
rect 2012 38598 2014 38650
rect 2194 38598 2196 38650
rect 1950 38596 1956 38598
rect 2012 38596 2036 38598
rect 2092 38596 2116 38598
rect 2172 38596 2196 38598
rect 2252 38596 2258 38598
rect 1950 38587 2258 38596
rect 1950 37564 2258 37573
rect 1950 37562 1956 37564
rect 2012 37562 2036 37564
rect 2092 37562 2116 37564
rect 2172 37562 2196 37564
rect 2252 37562 2258 37564
rect 2012 37510 2014 37562
rect 2194 37510 2196 37562
rect 1950 37508 1956 37510
rect 2012 37508 2036 37510
rect 2092 37508 2116 37510
rect 2172 37508 2196 37510
rect 2252 37508 2258 37510
rect 1950 37499 2258 37508
rect 2412 36780 2464 36786
rect 2412 36722 2464 36728
rect 1950 36476 2258 36485
rect 1950 36474 1956 36476
rect 2012 36474 2036 36476
rect 2092 36474 2116 36476
rect 2172 36474 2196 36476
rect 2252 36474 2258 36476
rect 2012 36422 2014 36474
rect 2194 36422 2196 36474
rect 1950 36420 1956 36422
rect 2012 36420 2036 36422
rect 2092 36420 2116 36422
rect 2172 36420 2196 36422
rect 2252 36420 2258 36422
rect 1950 36411 2258 36420
rect 1950 35388 2258 35397
rect 1950 35386 1956 35388
rect 2012 35386 2036 35388
rect 2092 35386 2116 35388
rect 2172 35386 2196 35388
rect 2252 35386 2258 35388
rect 2012 35334 2014 35386
rect 2194 35334 2196 35386
rect 1950 35332 1956 35334
rect 2012 35332 2036 35334
rect 2092 35332 2116 35334
rect 2172 35332 2196 35334
rect 2252 35332 2258 35334
rect 1950 35323 2258 35332
rect 2320 34536 2372 34542
rect 2320 34478 2372 34484
rect 1950 34300 2258 34309
rect 1950 34298 1956 34300
rect 2012 34298 2036 34300
rect 2092 34298 2116 34300
rect 2172 34298 2196 34300
rect 2252 34298 2258 34300
rect 2012 34246 2014 34298
rect 2194 34246 2196 34298
rect 1950 34244 1956 34246
rect 2012 34244 2036 34246
rect 2092 34244 2116 34246
rect 2172 34244 2196 34246
rect 2252 34244 2258 34246
rect 1950 34235 2258 34244
rect 1950 33212 2258 33221
rect 1950 33210 1956 33212
rect 2012 33210 2036 33212
rect 2092 33210 2116 33212
rect 2172 33210 2196 33212
rect 2252 33210 2258 33212
rect 2012 33158 2014 33210
rect 2194 33158 2196 33210
rect 1950 33156 1956 33158
rect 2012 33156 2036 33158
rect 2092 33156 2116 33158
rect 2172 33156 2196 33158
rect 2252 33156 2258 33158
rect 1950 33147 2258 33156
rect 1950 32124 2258 32133
rect 1950 32122 1956 32124
rect 2012 32122 2036 32124
rect 2092 32122 2116 32124
rect 2172 32122 2196 32124
rect 2252 32122 2258 32124
rect 2012 32070 2014 32122
rect 2194 32070 2196 32122
rect 1950 32068 1956 32070
rect 2012 32068 2036 32070
rect 2092 32068 2116 32070
rect 2172 32068 2196 32070
rect 2252 32068 2258 32070
rect 1950 32059 2258 32068
rect 1950 31036 2258 31045
rect 1950 31034 1956 31036
rect 2012 31034 2036 31036
rect 2092 31034 2116 31036
rect 2172 31034 2196 31036
rect 2252 31034 2258 31036
rect 2012 30982 2014 31034
rect 2194 30982 2196 31034
rect 1950 30980 1956 30982
rect 2012 30980 2036 30982
rect 2092 30980 2116 30982
rect 2172 30980 2196 30982
rect 2252 30980 2258 30982
rect 1950 30971 2258 30980
rect 1950 29948 2258 29957
rect 1950 29946 1956 29948
rect 2012 29946 2036 29948
rect 2092 29946 2116 29948
rect 2172 29946 2196 29948
rect 2252 29946 2258 29948
rect 2012 29894 2014 29946
rect 2194 29894 2196 29946
rect 1950 29892 1956 29894
rect 2012 29892 2036 29894
rect 2092 29892 2116 29894
rect 2172 29892 2196 29894
rect 2252 29892 2258 29894
rect 1950 29883 2258 29892
rect 1950 28860 2258 28869
rect 1950 28858 1956 28860
rect 2012 28858 2036 28860
rect 2092 28858 2116 28860
rect 2172 28858 2196 28860
rect 2252 28858 2258 28860
rect 2012 28806 2014 28858
rect 2194 28806 2196 28858
rect 1950 28804 1956 28806
rect 2012 28804 2036 28806
rect 2092 28804 2116 28806
rect 2172 28804 2196 28806
rect 2252 28804 2258 28806
rect 1950 28795 2258 28804
rect 1950 27772 2258 27781
rect 1950 27770 1956 27772
rect 2012 27770 2036 27772
rect 2092 27770 2116 27772
rect 2172 27770 2196 27772
rect 2252 27770 2258 27772
rect 2012 27718 2014 27770
rect 2194 27718 2196 27770
rect 1950 27716 1956 27718
rect 2012 27716 2036 27718
rect 2092 27716 2116 27718
rect 2172 27716 2196 27718
rect 2252 27716 2258 27718
rect 1950 27707 2258 27716
rect 1950 26684 2258 26693
rect 1950 26682 1956 26684
rect 2012 26682 2036 26684
rect 2092 26682 2116 26684
rect 2172 26682 2196 26684
rect 2252 26682 2258 26684
rect 2012 26630 2014 26682
rect 2194 26630 2196 26682
rect 1950 26628 1956 26630
rect 2012 26628 2036 26630
rect 2092 26628 2116 26630
rect 2172 26628 2196 26630
rect 2252 26628 2258 26630
rect 1950 26619 2258 26628
rect 1950 25596 2258 25605
rect 1950 25594 1956 25596
rect 2012 25594 2036 25596
rect 2092 25594 2116 25596
rect 2172 25594 2196 25596
rect 2252 25594 2258 25596
rect 2012 25542 2014 25594
rect 2194 25542 2196 25594
rect 1950 25540 1956 25542
rect 2012 25540 2036 25542
rect 2092 25540 2116 25542
rect 2172 25540 2196 25542
rect 2252 25540 2258 25542
rect 1950 25531 2258 25540
rect 1860 25492 1912 25498
rect 1860 25434 1912 25440
rect 1950 24508 2258 24517
rect 1950 24506 1956 24508
rect 2012 24506 2036 24508
rect 2092 24506 2116 24508
rect 2172 24506 2196 24508
rect 2252 24506 2258 24508
rect 2012 24454 2014 24506
rect 2194 24454 2196 24506
rect 1950 24452 1956 24454
rect 2012 24452 2036 24454
rect 2092 24452 2116 24454
rect 2172 24452 2196 24454
rect 2252 24452 2258 24454
rect 1950 24443 2258 24452
rect 1950 23420 2258 23429
rect 1950 23418 1956 23420
rect 2012 23418 2036 23420
rect 2092 23418 2116 23420
rect 2172 23418 2196 23420
rect 2252 23418 2258 23420
rect 2012 23366 2014 23418
rect 2194 23366 2196 23418
rect 1950 23364 1956 23366
rect 2012 23364 2036 23366
rect 2092 23364 2116 23366
rect 2172 23364 2196 23366
rect 2252 23364 2258 23366
rect 1950 23355 2258 23364
rect 1950 22332 2258 22341
rect 1950 22330 1956 22332
rect 2012 22330 2036 22332
rect 2092 22330 2116 22332
rect 2172 22330 2196 22332
rect 2252 22330 2258 22332
rect 2012 22278 2014 22330
rect 2194 22278 2196 22330
rect 1950 22276 1956 22278
rect 2012 22276 2036 22278
rect 2092 22276 2116 22278
rect 2172 22276 2196 22278
rect 2252 22276 2258 22278
rect 1950 22267 2258 22276
rect 1950 21244 2258 21253
rect 1950 21242 1956 21244
rect 2012 21242 2036 21244
rect 2092 21242 2116 21244
rect 2172 21242 2196 21244
rect 2252 21242 2258 21244
rect 2012 21190 2014 21242
rect 2194 21190 2196 21242
rect 1950 21188 1956 21190
rect 2012 21188 2036 21190
rect 2092 21188 2116 21190
rect 2172 21188 2196 21190
rect 2252 21188 2258 21190
rect 1950 21179 2258 21188
rect 1950 20156 2258 20165
rect 1950 20154 1956 20156
rect 2012 20154 2036 20156
rect 2092 20154 2116 20156
rect 2172 20154 2196 20156
rect 2252 20154 2258 20156
rect 2012 20102 2014 20154
rect 2194 20102 2196 20154
rect 1950 20100 1956 20102
rect 2012 20100 2036 20102
rect 2092 20100 2116 20102
rect 2172 20100 2196 20102
rect 2252 20100 2258 20102
rect 1950 20091 2258 20100
rect 1950 19068 2258 19077
rect 1950 19066 1956 19068
rect 2012 19066 2036 19068
rect 2092 19066 2116 19068
rect 2172 19066 2196 19068
rect 2252 19066 2258 19068
rect 2012 19014 2014 19066
rect 2194 19014 2196 19066
rect 1950 19012 1956 19014
rect 2012 19012 2036 19014
rect 2092 19012 2116 19014
rect 2172 19012 2196 19014
rect 2252 19012 2258 19014
rect 1950 19003 2258 19012
rect 1950 17980 2258 17989
rect 1950 17978 1956 17980
rect 2012 17978 2036 17980
rect 2092 17978 2116 17980
rect 2172 17978 2196 17980
rect 2252 17978 2258 17980
rect 2012 17926 2014 17978
rect 2194 17926 2196 17978
rect 1950 17924 1956 17926
rect 2012 17924 2036 17926
rect 2092 17924 2116 17926
rect 2172 17924 2196 17926
rect 2252 17924 2258 17926
rect 1950 17915 2258 17924
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 1858 16280 1914 16289
rect 1858 16215 1860 16224
rect 1912 16215 1914 16224
rect 1860 16186 1912 16192
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 2332 15706 2360 34478
rect 2424 27305 2452 36722
rect 2410 27296 2466 27305
rect 2410 27231 2466 27240
rect 2504 25900 2556 25906
rect 2504 25842 2556 25848
rect 2412 24880 2464 24886
rect 2412 24822 2464 24828
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 2424 14618 2452 24822
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 1858 13832 1914 13841
rect 1858 13767 1914 13776
rect 1872 13530 1900 13767
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 1858 11656 1914 11665
rect 1858 11591 1914 11600
rect 1872 11354 1900 11591
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 2516 8294 2544 25842
rect 2608 20058 2636 42162
rect 2688 42152 2740 42158
rect 2688 42094 2740 42100
rect 2700 26042 2728 42094
rect 3010 41372 3318 41381
rect 3010 41370 3016 41372
rect 3072 41370 3096 41372
rect 3152 41370 3176 41372
rect 3232 41370 3256 41372
rect 3312 41370 3318 41372
rect 3072 41318 3074 41370
rect 3254 41318 3256 41370
rect 3010 41316 3016 41318
rect 3072 41316 3096 41318
rect 3152 41316 3176 41318
rect 3232 41316 3256 41318
rect 3312 41316 3318 41318
rect 3010 41307 3318 41316
rect 3010 40284 3318 40293
rect 3010 40282 3016 40284
rect 3072 40282 3096 40284
rect 3152 40282 3176 40284
rect 3232 40282 3256 40284
rect 3312 40282 3318 40284
rect 3072 40230 3074 40282
rect 3254 40230 3256 40282
rect 3010 40228 3016 40230
rect 3072 40228 3096 40230
rect 3152 40228 3176 40230
rect 3232 40228 3256 40230
rect 3312 40228 3318 40230
rect 3010 40219 3318 40228
rect 3010 39196 3318 39205
rect 3010 39194 3016 39196
rect 3072 39194 3096 39196
rect 3152 39194 3176 39196
rect 3232 39194 3256 39196
rect 3312 39194 3318 39196
rect 3072 39142 3074 39194
rect 3254 39142 3256 39194
rect 3010 39140 3016 39142
rect 3072 39140 3096 39142
rect 3152 39140 3176 39142
rect 3232 39140 3256 39142
rect 3312 39140 3318 39142
rect 3010 39131 3318 39140
rect 3010 38108 3318 38117
rect 3010 38106 3016 38108
rect 3072 38106 3096 38108
rect 3152 38106 3176 38108
rect 3232 38106 3256 38108
rect 3312 38106 3318 38108
rect 3072 38054 3074 38106
rect 3254 38054 3256 38106
rect 3010 38052 3016 38054
rect 3072 38052 3096 38054
rect 3152 38052 3176 38054
rect 3232 38052 3256 38054
rect 3312 38052 3318 38054
rect 3010 38043 3318 38052
rect 3010 37020 3318 37029
rect 3010 37018 3016 37020
rect 3072 37018 3096 37020
rect 3152 37018 3176 37020
rect 3232 37018 3256 37020
rect 3312 37018 3318 37020
rect 3072 36966 3074 37018
rect 3254 36966 3256 37018
rect 3010 36964 3016 36966
rect 3072 36964 3096 36966
rect 3152 36964 3176 36966
rect 3232 36964 3256 36966
rect 3312 36964 3318 36966
rect 3010 36955 3318 36964
rect 3010 35932 3318 35941
rect 3010 35930 3016 35932
rect 3072 35930 3096 35932
rect 3152 35930 3176 35932
rect 3232 35930 3256 35932
rect 3312 35930 3318 35932
rect 3072 35878 3074 35930
rect 3254 35878 3256 35930
rect 3010 35876 3016 35878
rect 3072 35876 3096 35878
rect 3152 35876 3176 35878
rect 3232 35876 3256 35878
rect 3312 35876 3318 35878
rect 3010 35867 3318 35876
rect 3010 34844 3318 34853
rect 3010 34842 3016 34844
rect 3072 34842 3096 34844
rect 3152 34842 3176 34844
rect 3232 34842 3256 34844
rect 3312 34842 3318 34844
rect 3072 34790 3074 34842
rect 3254 34790 3256 34842
rect 3010 34788 3016 34790
rect 3072 34788 3096 34790
rect 3152 34788 3176 34790
rect 3232 34788 3256 34790
rect 3312 34788 3318 34790
rect 3010 34779 3318 34788
rect 3010 33756 3318 33765
rect 3010 33754 3016 33756
rect 3072 33754 3096 33756
rect 3152 33754 3176 33756
rect 3232 33754 3256 33756
rect 3312 33754 3318 33756
rect 3072 33702 3074 33754
rect 3254 33702 3256 33754
rect 3010 33700 3016 33702
rect 3072 33700 3096 33702
rect 3152 33700 3176 33702
rect 3232 33700 3256 33702
rect 3312 33700 3318 33702
rect 3010 33691 3318 33700
rect 3010 32668 3318 32677
rect 3010 32666 3016 32668
rect 3072 32666 3096 32668
rect 3152 32666 3176 32668
rect 3232 32666 3256 32668
rect 3312 32666 3318 32668
rect 3072 32614 3074 32666
rect 3254 32614 3256 32666
rect 3010 32612 3016 32614
rect 3072 32612 3096 32614
rect 3152 32612 3176 32614
rect 3232 32612 3256 32614
rect 3312 32612 3318 32614
rect 3010 32603 3318 32612
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2792 31142 2820 31758
rect 3010 31580 3318 31589
rect 3010 31578 3016 31580
rect 3072 31578 3096 31580
rect 3152 31578 3176 31580
rect 3232 31578 3256 31580
rect 3312 31578 3318 31580
rect 3072 31526 3074 31578
rect 3254 31526 3256 31578
rect 3010 31524 3016 31526
rect 3072 31524 3096 31526
rect 3152 31524 3176 31526
rect 3232 31524 3256 31526
rect 3312 31524 3318 31526
rect 3010 31515 3318 31524
rect 2780 31136 2832 31142
rect 2780 31078 2832 31084
rect 2688 26036 2740 26042
rect 2688 25978 2740 25984
rect 2688 22704 2740 22710
rect 2688 22646 2740 22652
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2700 12442 2728 22646
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2516 8266 2728 8294
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2700 2650 2728 8266
rect 2792 6905 2820 31078
rect 3010 30492 3318 30501
rect 3010 30490 3016 30492
rect 3072 30490 3096 30492
rect 3152 30490 3176 30492
rect 3232 30490 3256 30492
rect 3312 30490 3318 30492
rect 3072 30438 3074 30490
rect 3254 30438 3256 30490
rect 3010 30436 3016 30438
rect 3072 30436 3096 30438
rect 3152 30436 3176 30438
rect 3232 30436 3256 30438
rect 3312 30436 3318 30438
rect 3010 30427 3318 30436
rect 3010 29404 3318 29413
rect 3010 29402 3016 29404
rect 3072 29402 3096 29404
rect 3152 29402 3176 29404
rect 3232 29402 3256 29404
rect 3312 29402 3318 29404
rect 3072 29350 3074 29402
rect 3254 29350 3256 29402
rect 3010 29348 3016 29350
rect 3072 29348 3096 29350
rect 3152 29348 3176 29350
rect 3232 29348 3256 29350
rect 3312 29348 3318 29350
rect 3010 29339 3318 29348
rect 3010 28316 3318 28325
rect 3010 28314 3016 28316
rect 3072 28314 3096 28316
rect 3152 28314 3176 28316
rect 3232 28314 3256 28316
rect 3312 28314 3318 28316
rect 3072 28262 3074 28314
rect 3254 28262 3256 28314
rect 3010 28260 3016 28262
rect 3072 28260 3096 28262
rect 3152 28260 3176 28262
rect 3232 28260 3256 28262
rect 3312 28260 3318 28262
rect 3010 28251 3318 28260
rect 3010 27228 3318 27237
rect 3010 27226 3016 27228
rect 3072 27226 3096 27228
rect 3152 27226 3176 27228
rect 3232 27226 3256 27228
rect 3312 27226 3318 27228
rect 3072 27174 3074 27226
rect 3254 27174 3256 27226
rect 3010 27172 3016 27174
rect 3072 27172 3096 27174
rect 3152 27172 3176 27174
rect 3232 27172 3256 27174
rect 3312 27172 3318 27174
rect 3010 27163 3318 27172
rect 2872 26308 2924 26314
rect 2872 26250 2924 26256
rect 2884 11121 2912 26250
rect 3010 26140 3318 26149
rect 3010 26138 3016 26140
rect 3072 26138 3096 26140
rect 3152 26138 3176 26140
rect 3232 26138 3256 26140
rect 3312 26138 3318 26140
rect 3072 26086 3074 26138
rect 3254 26086 3256 26138
rect 3010 26084 3016 26086
rect 3072 26084 3096 26086
rect 3152 26084 3176 26086
rect 3232 26084 3256 26086
rect 3312 26084 3318 26086
rect 3010 26075 3318 26084
rect 3056 25900 3108 25906
rect 3056 25842 3108 25848
rect 3068 25265 3096 25842
rect 3054 25256 3110 25265
rect 3054 25191 3056 25200
rect 3108 25191 3110 25200
rect 3056 25162 3108 25168
rect 3010 25052 3318 25061
rect 3010 25050 3016 25052
rect 3072 25050 3096 25052
rect 3152 25050 3176 25052
rect 3232 25050 3256 25052
rect 3312 25050 3318 25052
rect 3072 24998 3074 25050
rect 3254 24998 3256 25050
rect 3010 24996 3016 24998
rect 3072 24996 3096 24998
rect 3152 24996 3176 24998
rect 3232 24996 3256 24998
rect 3312 24996 3318 24998
rect 3010 24987 3318 24996
rect 3436 24410 3464 42162
rect 3516 32836 3568 32842
rect 3516 32778 3568 32784
rect 3528 32026 3556 32778
rect 3516 32020 3568 32026
rect 3516 31962 3568 31968
rect 3516 31884 3568 31890
rect 3516 31826 3568 31832
rect 3424 24404 3476 24410
rect 3424 24346 3476 24352
rect 3424 24268 3476 24274
rect 3424 24210 3476 24216
rect 3010 23964 3318 23973
rect 3010 23962 3016 23964
rect 3072 23962 3096 23964
rect 3152 23962 3176 23964
rect 3232 23962 3256 23964
rect 3312 23962 3318 23964
rect 3072 23910 3074 23962
rect 3254 23910 3256 23962
rect 3010 23908 3016 23910
rect 3072 23908 3096 23910
rect 3152 23908 3176 23910
rect 3232 23908 3256 23910
rect 3312 23908 3318 23910
rect 3010 23899 3318 23908
rect 3010 22876 3318 22885
rect 3010 22874 3016 22876
rect 3072 22874 3096 22876
rect 3152 22874 3176 22876
rect 3232 22874 3256 22876
rect 3312 22874 3318 22876
rect 3072 22822 3074 22874
rect 3254 22822 3256 22874
rect 3010 22820 3016 22822
rect 3072 22820 3096 22822
rect 3152 22820 3176 22822
rect 3232 22820 3256 22822
rect 3312 22820 3318 22822
rect 3010 22811 3318 22820
rect 3010 21788 3318 21797
rect 3010 21786 3016 21788
rect 3072 21786 3096 21788
rect 3152 21786 3176 21788
rect 3232 21786 3256 21788
rect 3312 21786 3318 21788
rect 3072 21734 3074 21786
rect 3254 21734 3256 21786
rect 3010 21732 3016 21734
rect 3072 21732 3096 21734
rect 3152 21732 3176 21734
rect 3232 21732 3256 21734
rect 3312 21732 3318 21734
rect 3010 21723 3318 21732
rect 3010 20700 3318 20709
rect 3010 20698 3016 20700
rect 3072 20698 3096 20700
rect 3152 20698 3176 20700
rect 3232 20698 3256 20700
rect 3312 20698 3318 20700
rect 3072 20646 3074 20698
rect 3254 20646 3256 20698
rect 3010 20644 3016 20646
rect 3072 20644 3096 20646
rect 3152 20644 3176 20646
rect 3232 20644 3256 20646
rect 3312 20644 3318 20646
rect 3010 20635 3318 20644
rect 3010 19612 3318 19621
rect 3010 19610 3016 19612
rect 3072 19610 3096 19612
rect 3152 19610 3176 19612
rect 3232 19610 3256 19612
rect 3312 19610 3318 19612
rect 3072 19558 3074 19610
rect 3254 19558 3256 19610
rect 3010 19556 3016 19558
rect 3072 19556 3096 19558
rect 3152 19556 3176 19558
rect 3232 19556 3256 19558
rect 3312 19556 3318 19558
rect 3010 19547 3318 19556
rect 3436 19514 3464 24210
rect 3528 21690 3556 31826
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3514 19544 3570 19553
rect 3424 19508 3476 19514
rect 3620 19514 3648 42162
rect 3700 35012 3752 35018
rect 3700 34954 3752 34960
rect 3712 31890 3740 34954
rect 3700 31884 3752 31890
rect 3700 31826 3752 31832
rect 3698 31784 3754 31793
rect 3698 31719 3754 31728
rect 3712 24342 3740 31719
rect 3700 24336 3752 24342
rect 3700 24278 3752 24284
rect 3700 24200 3752 24206
rect 3700 24142 3752 24148
rect 3712 23497 3740 24142
rect 3698 23488 3754 23497
rect 3698 23423 3754 23432
rect 3804 22778 3832 42162
rect 3976 36712 4028 36718
rect 3976 36654 4028 36660
rect 3884 35148 3936 35154
rect 3884 35090 3936 35096
rect 3896 31793 3924 35090
rect 3882 31784 3938 31793
rect 3882 31719 3938 31728
rect 3988 27606 4016 36654
rect 4344 35692 4396 35698
rect 4344 35634 4396 35640
rect 4356 33658 4384 35634
rect 4344 33652 4396 33658
rect 4344 33594 4396 33600
rect 4068 31816 4120 31822
rect 4068 31758 4120 31764
rect 3976 27600 4028 27606
rect 3976 27542 4028 27548
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 3792 21480 3844 21486
rect 3792 21422 3844 21428
rect 3514 19479 3516 19488
rect 3424 19450 3476 19456
rect 3568 19479 3570 19488
rect 3608 19508 3660 19514
rect 3516 19450 3568 19456
rect 3608 19450 3660 19456
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3010 18524 3318 18533
rect 3010 18522 3016 18524
rect 3072 18522 3096 18524
rect 3152 18522 3176 18524
rect 3232 18522 3256 18524
rect 3312 18522 3318 18524
rect 3072 18470 3074 18522
rect 3254 18470 3256 18522
rect 3010 18468 3016 18470
rect 3072 18468 3096 18470
rect 3152 18468 3176 18470
rect 3232 18468 3256 18470
rect 3312 18468 3318 18470
rect 3010 18459 3318 18468
rect 3010 17436 3318 17445
rect 3010 17434 3016 17436
rect 3072 17434 3096 17436
rect 3152 17434 3176 17436
rect 3232 17434 3256 17436
rect 3312 17434 3318 17436
rect 3072 17382 3074 17434
rect 3254 17382 3256 17434
rect 3010 17380 3016 17382
rect 3072 17380 3096 17382
rect 3152 17380 3176 17382
rect 3232 17380 3256 17382
rect 3312 17380 3318 17382
rect 3010 17371 3318 17380
rect 3010 16348 3318 16357
rect 3010 16346 3016 16348
rect 3072 16346 3096 16348
rect 3152 16346 3176 16348
rect 3232 16346 3256 16348
rect 3312 16346 3318 16348
rect 3072 16294 3074 16346
rect 3254 16294 3256 16346
rect 3010 16292 3016 16294
rect 3072 16292 3096 16294
rect 3152 16292 3176 16294
rect 3232 16292 3256 16294
rect 3312 16292 3318 16294
rect 3010 16283 3318 16292
rect 3010 15260 3318 15269
rect 3010 15258 3016 15260
rect 3072 15258 3096 15260
rect 3152 15258 3176 15260
rect 3232 15258 3256 15260
rect 3312 15258 3318 15260
rect 3072 15206 3074 15258
rect 3254 15206 3256 15258
rect 3010 15204 3016 15206
rect 3072 15204 3096 15206
rect 3152 15204 3176 15206
rect 3232 15204 3256 15206
rect 3312 15204 3318 15206
rect 3010 15195 3318 15204
rect 3010 14172 3318 14181
rect 3010 14170 3016 14172
rect 3072 14170 3096 14172
rect 3152 14170 3176 14172
rect 3232 14170 3256 14172
rect 3312 14170 3318 14172
rect 3072 14118 3074 14170
rect 3254 14118 3256 14170
rect 3010 14116 3016 14118
rect 3072 14116 3096 14118
rect 3152 14116 3176 14118
rect 3232 14116 3256 14118
rect 3312 14116 3318 14118
rect 3010 14107 3318 14116
rect 3010 13084 3318 13093
rect 3010 13082 3016 13084
rect 3072 13082 3096 13084
rect 3152 13082 3176 13084
rect 3232 13082 3256 13084
rect 3312 13082 3318 13084
rect 3072 13030 3074 13082
rect 3254 13030 3256 13082
rect 3010 13028 3016 13030
rect 3072 13028 3096 13030
rect 3152 13028 3176 13030
rect 3232 13028 3256 13030
rect 3312 13028 3318 13030
rect 3010 13019 3318 13028
rect 3010 11996 3318 12005
rect 3010 11994 3016 11996
rect 3072 11994 3096 11996
rect 3152 11994 3176 11996
rect 3232 11994 3256 11996
rect 3312 11994 3318 11996
rect 3072 11942 3074 11994
rect 3254 11942 3256 11994
rect 3010 11940 3016 11942
rect 3072 11940 3096 11942
rect 3152 11940 3176 11942
rect 3232 11940 3256 11942
rect 3312 11940 3318 11942
rect 3010 11931 3318 11940
rect 2870 11112 2926 11121
rect 2870 11047 2926 11056
rect 3010 10908 3318 10917
rect 3010 10906 3016 10908
rect 3072 10906 3096 10908
rect 3152 10906 3176 10908
rect 3232 10906 3256 10908
rect 3312 10906 3318 10908
rect 3072 10854 3074 10906
rect 3254 10854 3256 10906
rect 3010 10852 3016 10854
rect 3072 10852 3096 10854
rect 3152 10852 3176 10854
rect 3232 10852 3256 10854
rect 3312 10852 3318 10854
rect 3010 10843 3318 10852
rect 3010 9820 3318 9829
rect 3010 9818 3016 9820
rect 3072 9818 3096 9820
rect 3152 9818 3176 9820
rect 3232 9818 3256 9820
rect 3312 9818 3318 9820
rect 3072 9766 3074 9818
rect 3254 9766 3256 9818
rect 3010 9764 3016 9766
rect 3072 9764 3096 9766
rect 3152 9764 3176 9766
rect 3232 9764 3256 9766
rect 3312 9764 3318 9766
rect 3010 9755 3318 9764
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 3436 3466 3464 19314
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 1596 56 1716 82
rect 2148 56 2176 2586
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 2596 2100 2648 2106
rect 2596 2042 2648 2048
rect 2608 56 2636 2042
rect 3054 1320 3110 1329
rect 3054 1255 3110 1264
rect 3068 56 3096 1255
rect 3528 56 3556 19314
rect 3804 4010 3832 21422
rect 3988 21350 4016 22578
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3896 3738 3924 19654
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3988 56 4016 21286
rect 4080 16153 4108 31758
rect 4540 29073 4568 42230
rect 4896 42220 4948 42226
rect 4896 42162 4948 42168
rect 4988 42220 5040 42226
rect 4988 42162 5040 42168
rect 5632 42220 5684 42226
rect 5632 42162 5684 42168
rect 5908 42220 5960 42226
rect 5908 42162 5960 42168
rect 7012 42220 7064 42226
rect 7012 42162 7064 42168
rect 4712 42152 4764 42158
rect 4712 42094 4764 42100
rect 4526 29064 4582 29073
rect 4526 28999 4582 29008
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 4448 56 4476 19790
rect 4540 474 4568 21966
rect 4724 21894 4752 42094
rect 4804 29028 4856 29034
rect 4804 28970 4856 28976
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4816 18426 4844 28970
rect 4908 20058 4936 42162
rect 5000 41449 5028 42162
rect 5448 42084 5500 42090
rect 5448 42026 5500 42032
rect 5080 42016 5132 42022
rect 5080 41958 5132 41964
rect 4986 41440 5042 41449
rect 4986 41375 5042 41384
rect 5092 24410 5120 41958
rect 5356 36100 5408 36106
rect 5356 36042 5408 36048
rect 5368 35290 5396 36042
rect 5356 35284 5408 35290
rect 5356 35226 5408 35232
rect 5172 30728 5224 30734
rect 5172 30670 5224 30676
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 5000 23526 5028 24142
rect 4988 23520 5040 23526
rect 4986 23488 4988 23497
rect 5040 23488 5042 23497
rect 4986 23423 5042 23432
rect 5184 23338 5212 30670
rect 5356 30660 5408 30666
rect 5356 30602 5408 30608
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5000 23310 5212 23338
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4632 8265 4660 18226
rect 5000 16425 5028 23310
rect 5276 22930 5304 23666
rect 5184 22902 5304 22930
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 4986 16416 5042 16425
rect 4986 16351 5042 16360
rect 4894 16280 4950 16289
rect 4894 16215 4896 16224
rect 4948 16215 4950 16224
rect 4896 16186 4948 16192
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4618 8256 4674 8265
rect 4618 8191 4674 8200
rect 4528 468 4580 474
rect 4528 410 4580 416
rect 4908 56 4936 16050
rect 5092 15609 5120 20402
rect 5078 15600 5134 15609
rect 5078 15535 5134 15544
rect 5184 9178 5212 22902
rect 5368 22094 5396 30602
rect 5460 26042 5488 42026
rect 5538 39536 5594 39545
rect 5538 39471 5594 39480
rect 5552 39438 5580 39471
rect 5540 39432 5592 39438
rect 5540 39374 5592 39380
rect 5540 38344 5592 38350
rect 5538 38312 5540 38321
rect 5592 38312 5594 38321
rect 5538 38247 5594 38256
rect 5448 26036 5500 26042
rect 5448 25978 5500 25984
rect 5644 22094 5672 42162
rect 5724 40384 5776 40390
rect 5724 40326 5776 40332
rect 5736 38418 5764 40326
rect 5724 38412 5776 38418
rect 5724 38354 5776 38360
rect 5724 37120 5776 37126
rect 5724 37062 5776 37068
rect 5736 29306 5764 37062
rect 5724 29300 5776 29306
rect 5724 29242 5776 29248
rect 5920 29034 5948 42162
rect 6092 41676 6144 41682
rect 6092 41618 6144 41624
rect 6000 39296 6052 39302
rect 6000 39238 6052 39244
rect 6012 37942 6040 39238
rect 6000 37936 6052 37942
rect 6000 37878 6052 37884
rect 5908 29028 5960 29034
rect 5908 28970 5960 28976
rect 5816 22568 5868 22574
rect 5816 22510 5868 22516
rect 5276 22066 5396 22094
rect 5552 22066 5672 22094
rect 5276 20602 5304 22066
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5276 2922 5304 19382
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 5368 56 5396 20402
rect 5460 2650 5488 21286
rect 5552 20602 5580 22066
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 5828 11354 5856 22510
rect 6104 22094 6132 41618
rect 6736 41064 6788 41070
rect 6736 41006 6788 41012
rect 6184 35624 6236 35630
rect 6184 35566 6236 35572
rect 6196 22506 6224 35566
rect 6368 33992 6420 33998
rect 6368 33934 6420 33940
rect 6276 32904 6328 32910
rect 6276 32846 6328 32852
rect 6288 23594 6316 32846
rect 6380 24886 6408 33934
rect 6748 31754 6776 41006
rect 6828 38208 6880 38214
rect 6828 38150 6880 38156
rect 6840 37194 6868 38150
rect 6920 37256 6972 37262
rect 6920 37198 6972 37204
rect 6828 37188 6880 37194
rect 6828 37130 6880 37136
rect 6932 35601 6960 37198
rect 6918 35592 6974 35601
rect 6918 35527 6974 35536
rect 7024 31754 7052 42162
rect 7104 41540 7156 41546
rect 7104 41482 7156 41488
rect 6748 31726 6868 31754
rect 6644 31272 6696 31278
rect 6644 31214 6696 31220
rect 6552 25832 6604 25838
rect 6552 25774 6604 25780
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 6368 24880 6420 24886
rect 6368 24822 6420 24828
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6276 23588 6328 23594
rect 6276 23530 6328 23536
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 5920 22066 6132 22094
rect 5920 21962 5948 22066
rect 5908 21956 5960 21962
rect 5908 21898 5960 21904
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5920 8634 5948 19790
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 5998 11656 6054 11665
rect 5998 11591 6054 11600
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5722 8256 5778 8265
rect 5722 8191 5778 8200
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5736 2122 5764 8191
rect 5814 7304 5870 7313
rect 5814 7239 5870 7248
rect 5828 5710 5856 7239
rect 5906 6216 5962 6225
rect 5906 6151 5962 6160
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5920 3058 5948 6151
rect 6012 5914 6040 11591
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6104 3194 6132 18566
rect 6196 17746 6224 22170
rect 6276 18896 6328 18902
rect 6276 18838 6328 18844
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6182 13832 6238 13841
rect 6182 13767 6238 13776
rect 6196 4826 6224 13767
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6288 3194 6316 18838
rect 6380 17882 6408 24006
rect 6472 22234 6500 25162
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 6564 22094 6592 25774
rect 6472 22066 6592 22094
rect 6472 20618 6500 22066
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6564 20806 6592 21966
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6472 20590 6592 20618
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6380 16250 6408 17682
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6472 15473 6500 19314
rect 6458 15464 6514 15473
rect 6458 15399 6514 15408
rect 6564 15162 6592 20590
rect 6656 19514 6684 31214
rect 6736 27464 6788 27470
rect 6736 27406 6788 27412
rect 6748 23497 6776 27406
rect 6734 23488 6790 23497
rect 6734 23423 6790 23432
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6748 21049 6776 21966
rect 6840 21894 6868 31726
rect 6932 31726 7052 31754
rect 6932 22778 6960 31726
rect 7012 30864 7064 30870
rect 7012 30806 7064 30812
rect 7024 24993 7052 30806
rect 7010 24984 7066 24993
rect 7010 24919 7066 24928
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7024 24138 7052 24754
rect 7116 24682 7144 41482
rect 7392 41138 7420 43551
rect 7668 42362 7696 44960
rect 8128 42362 8156 44960
rect 7656 42356 7708 42362
rect 7656 42298 7708 42304
rect 8116 42356 8168 42362
rect 8116 42298 8168 42304
rect 7470 42256 7526 42265
rect 7470 42191 7526 42200
rect 7484 41614 7512 42191
rect 7950 41916 8258 41925
rect 7950 41914 7956 41916
rect 8012 41914 8036 41916
rect 8092 41914 8116 41916
rect 8172 41914 8196 41916
rect 8252 41914 8258 41916
rect 8012 41862 8014 41914
rect 8194 41862 8196 41914
rect 7950 41860 7956 41862
rect 8012 41860 8036 41862
rect 8092 41860 8116 41862
rect 8172 41860 8196 41862
rect 8252 41860 8258 41862
rect 7950 41851 8258 41860
rect 8588 41818 8616 44960
rect 8576 41812 8628 41818
rect 8576 41754 8628 41760
rect 9048 41750 9076 44960
rect 9036 41744 9088 41750
rect 9036 41686 9088 41692
rect 7472 41608 7524 41614
rect 7472 41550 7524 41556
rect 7840 41472 7892 41478
rect 7840 41414 7892 41420
rect 7380 41132 7432 41138
rect 7380 41074 7432 41080
rect 7748 40928 7800 40934
rect 7748 40870 7800 40876
rect 7654 40624 7710 40633
rect 7654 40559 7710 40568
rect 7668 40526 7696 40559
rect 7656 40520 7708 40526
rect 7656 40462 7708 40468
rect 7760 40050 7788 40870
rect 7852 40610 7880 41414
rect 9508 41274 9536 44960
rect 9496 41268 9548 41274
rect 9496 41210 9548 41216
rect 7950 40828 8258 40837
rect 7950 40826 7956 40828
rect 8012 40826 8036 40828
rect 8092 40826 8116 40828
rect 8172 40826 8196 40828
rect 8252 40826 8258 40828
rect 8012 40774 8014 40826
rect 8194 40774 8196 40826
rect 7950 40772 7956 40774
rect 8012 40772 8036 40774
rect 8092 40772 8116 40774
rect 8172 40772 8196 40774
rect 8252 40772 8258 40774
rect 7950 40763 8258 40772
rect 7852 40582 7972 40610
rect 7840 40384 7892 40390
rect 7840 40326 7892 40332
rect 7748 40044 7800 40050
rect 7748 39986 7800 39992
rect 7852 39438 7880 40326
rect 7944 40118 7972 40582
rect 7932 40112 7984 40118
rect 7932 40054 7984 40060
rect 7930 39944 7986 39953
rect 7930 39879 7932 39888
rect 7984 39879 7986 39888
rect 7932 39850 7984 39856
rect 8300 39840 8352 39846
rect 8300 39782 8352 39788
rect 7950 39740 8258 39749
rect 7950 39738 7956 39740
rect 8012 39738 8036 39740
rect 8092 39738 8116 39740
rect 8172 39738 8196 39740
rect 8252 39738 8258 39740
rect 8012 39686 8014 39738
rect 8194 39686 8196 39738
rect 7950 39684 7956 39686
rect 8012 39684 8036 39686
rect 8092 39684 8116 39686
rect 8172 39684 8196 39686
rect 8252 39684 8258 39686
rect 7950 39675 8258 39684
rect 8312 39545 8340 39782
rect 8298 39536 8354 39545
rect 8298 39471 8354 39480
rect 7840 39432 7892 39438
rect 7840 39374 7892 39380
rect 7932 39296 7984 39302
rect 7930 39264 7932 39273
rect 8300 39296 8352 39302
rect 7984 39264 7986 39273
rect 8300 39238 8352 39244
rect 7930 39199 7986 39208
rect 8312 39001 8340 39238
rect 8298 38992 8354 39001
rect 7748 38956 7800 38962
rect 7748 38898 7800 38904
rect 7840 38956 7892 38962
rect 8298 38927 8354 38936
rect 7840 38898 7892 38904
rect 7760 38554 7788 38898
rect 7748 38548 7800 38554
rect 7748 38490 7800 38496
rect 7748 38344 7800 38350
rect 7748 38286 7800 38292
rect 7472 37868 7524 37874
rect 7472 37810 7524 37816
rect 7656 37868 7708 37874
rect 7656 37810 7708 37816
rect 7484 36825 7512 37810
rect 7470 36816 7526 36825
rect 7470 36751 7526 36760
rect 7668 35290 7696 37810
rect 7760 37466 7788 38286
rect 7852 38010 7880 38898
rect 7930 38856 7986 38865
rect 7930 38791 7932 38800
rect 7984 38791 7986 38800
rect 7932 38762 7984 38768
rect 8300 38752 8352 38758
rect 8300 38694 8352 38700
rect 7950 38652 8258 38661
rect 7950 38650 7956 38652
rect 8012 38650 8036 38652
rect 8092 38650 8116 38652
rect 8172 38650 8196 38652
rect 8252 38650 8258 38652
rect 8012 38598 8014 38650
rect 8194 38598 8196 38650
rect 7950 38596 7956 38598
rect 8012 38596 8036 38598
rect 8092 38596 8116 38598
rect 8172 38596 8196 38598
rect 8252 38596 8258 38598
rect 7950 38587 8258 38596
rect 8312 38457 8340 38694
rect 8298 38448 8354 38457
rect 8298 38383 8354 38392
rect 7932 38208 7984 38214
rect 7930 38176 7932 38185
rect 8300 38208 8352 38214
rect 7984 38176 7986 38185
rect 8300 38150 8352 38156
rect 7930 38111 7986 38120
rect 7840 38004 7892 38010
rect 7840 37946 7892 37952
rect 8312 37913 8340 38150
rect 8298 37904 8354 37913
rect 8298 37839 8354 37848
rect 7930 37768 7986 37777
rect 7930 37703 7932 37712
rect 7984 37703 7986 37712
rect 7932 37674 7984 37680
rect 8300 37664 8352 37670
rect 8300 37606 8352 37612
rect 7950 37564 8258 37573
rect 7950 37562 7956 37564
rect 8012 37562 8036 37564
rect 8092 37562 8116 37564
rect 8172 37562 8196 37564
rect 8252 37562 8258 37564
rect 8012 37510 8014 37562
rect 8194 37510 8196 37562
rect 7950 37508 7956 37510
rect 8012 37508 8036 37510
rect 8092 37508 8116 37510
rect 8172 37508 8196 37510
rect 8252 37508 8258 37510
rect 7950 37499 8258 37508
rect 7748 37460 7800 37466
rect 7748 37402 7800 37408
rect 8312 37369 8340 37606
rect 8298 37360 8354 37369
rect 8298 37295 8354 37304
rect 7932 37120 7984 37126
rect 7930 37088 7932 37097
rect 8300 37120 8352 37126
rect 7984 37088 7986 37097
rect 8300 37062 8352 37068
rect 7930 37023 7986 37032
rect 8312 36825 8340 37062
rect 8298 36816 8354 36825
rect 8298 36751 8354 36760
rect 7930 36680 7986 36689
rect 7930 36615 7932 36624
rect 7984 36615 7986 36624
rect 7932 36586 7984 36592
rect 8300 36576 8352 36582
rect 8300 36518 8352 36524
rect 7950 36476 8258 36485
rect 7950 36474 7956 36476
rect 8012 36474 8036 36476
rect 8092 36474 8116 36476
rect 8172 36474 8196 36476
rect 8252 36474 8258 36476
rect 8012 36422 8014 36474
rect 8194 36422 8196 36474
rect 7950 36420 7956 36422
rect 8012 36420 8036 36422
rect 8092 36420 8116 36422
rect 8172 36420 8196 36422
rect 8252 36420 8258 36422
rect 7950 36411 8258 36420
rect 8312 36281 8340 36518
rect 8298 36272 8354 36281
rect 8298 36207 8354 36216
rect 7932 36032 7984 36038
rect 7930 36000 7932 36009
rect 8300 36032 8352 36038
rect 7984 36000 7986 36009
rect 8300 35974 8352 35980
rect 7930 35935 7986 35944
rect 8312 35737 8340 35974
rect 8298 35728 8354 35737
rect 8298 35663 8354 35672
rect 7930 35592 7986 35601
rect 7930 35527 7932 35536
rect 7984 35527 7986 35536
rect 7932 35498 7984 35504
rect 8300 35488 8352 35494
rect 8300 35430 8352 35436
rect 7950 35388 8258 35397
rect 7950 35386 7956 35388
rect 8012 35386 8036 35388
rect 8092 35386 8116 35388
rect 8172 35386 8196 35388
rect 8252 35386 8258 35388
rect 8012 35334 8014 35386
rect 8194 35334 8196 35386
rect 7950 35332 7956 35334
rect 8012 35332 8036 35334
rect 8092 35332 8116 35334
rect 8172 35332 8196 35334
rect 8252 35332 8258 35334
rect 7950 35323 8258 35332
rect 7656 35284 7708 35290
rect 7656 35226 7708 35232
rect 8312 35193 8340 35430
rect 8298 35184 8354 35193
rect 8298 35119 8354 35128
rect 7472 35080 7524 35086
rect 7472 35022 7524 35028
rect 7484 32881 7512 35022
rect 7932 34944 7984 34950
rect 7930 34912 7932 34921
rect 8300 34944 8352 34950
rect 7984 34912 7986 34921
rect 8300 34886 8352 34892
rect 7930 34847 7986 34856
rect 8312 34649 8340 34886
rect 8852 34740 8904 34746
rect 8852 34682 8904 34688
rect 8298 34640 8354 34649
rect 8298 34575 8354 34584
rect 8300 34400 8352 34406
rect 8864 34377 8892 34682
rect 8300 34342 8352 34348
rect 8850 34368 8906 34377
rect 7950 34300 8258 34309
rect 7950 34298 7956 34300
rect 8012 34298 8036 34300
rect 8092 34298 8116 34300
rect 8172 34298 8196 34300
rect 8252 34298 8258 34300
rect 8012 34246 8014 34298
rect 8194 34246 8196 34298
rect 7950 34244 7956 34246
rect 8012 34244 8036 34246
rect 8092 34244 8116 34246
rect 8172 34244 8196 34246
rect 8252 34244 8258 34246
rect 7950 34235 8258 34244
rect 8312 34105 8340 34342
rect 8850 34303 8906 34312
rect 8298 34096 8354 34105
rect 8298 34031 8354 34040
rect 8116 33992 8168 33998
rect 8116 33934 8168 33940
rect 7748 33856 7800 33862
rect 7932 33856 7984 33862
rect 7748 33798 7800 33804
rect 7930 33824 7932 33833
rect 7984 33824 7986 33833
rect 7760 33522 7788 33798
rect 7930 33759 7986 33768
rect 8128 33561 8156 33934
rect 8300 33856 8352 33862
rect 8300 33798 8352 33804
rect 8312 33561 8340 33798
rect 8114 33552 8170 33561
rect 7748 33516 7800 33522
rect 7748 33458 7800 33464
rect 7840 33516 7892 33522
rect 8114 33487 8170 33496
rect 8298 33552 8354 33561
rect 8298 33487 8354 33496
rect 7840 33458 7892 33464
rect 7852 33114 7880 33458
rect 7930 33416 7986 33425
rect 7930 33351 7932 33360
rect 7984 33351 7986 33360
rect 7932 33322 7984 33328
rect 8300 33312 8352 33318
rect 8300 33254 8352 33260
rect 7950 33212 8258 33221
rect 7950 33210 7956 33212
rect 8012 33210 8036 33212
rect 8092 33210 8116 33212
rect 8172 33210 8196 33212
rect 8252 33210 8258 33212
rect 8012 33158 8014 33210
rect 8194 33158 8196 33210
rect 7950 33156 7956 33158
rect 8012 33156 8036 33158
rect 8092 33156 8116 33158
rect 8172 33156 8196 33158
rect 8252 33156 8258 33158
rect 7950 33147 8258 33156
rect 7840 33108 7892 33114
rect 7840 33050 7892 33056
rect 8312 33017 8340 33254
rect 8298 33008 8354 33017
rect 8298 32943 8354 32952
rect 7748 32904 7800 32910
rect 7470 32872 7526 32881
rect 7748 32846 7800 32852
rect 7470 32807 7526 32816
rect 7760 32570 7788 32846
rect 7840 32768 7892 32774
rect 7932 32768 7984 32774
rect 7840 32710 7892 32716
rect 7930 32736 7932 32745
rect 8300 32768 8352 32774
rect 7984 32736 7986 32745
rect 7748 32564 7800 32570
rect 7748 32506 7800 32512
rect 7748 32428 7800 32434
rect 7748 32370 7800 32376
rect 7196 32360 7248 32366
rect 7196 32302 7248 32308
rect 7208 30054 7236 32302
rect 7472 31816 7524 31822
rect 7472 31758 7524 31764
rect 7380 31680 7432 31686
rect 7380 31622 7432 31628
rect 7392 30258 7420 31622
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 7484 30122 7512 31758
rect 7760 31482 7788 32370
rect 7852 31822 7880 32710
rect 8300 32710 8352 32716
rect 7930 32671 7986 32680
rect 8312 32473 8340 32710
rect 8298 32464 8354 32473
rect 8298 32399 8354 32408
rect 7930 32328 7986 32337
rect 7930 32263 7932 32272
rect 7984 32263 7986 32272
rect 7932 32234 7984 32240
rect 8300 32224 8352 32230
rect 8300 32166 8352 32172
rect 7950 32124 8258 32133
rect 7950 32122 7956 32124
rect 8012 32122 8036 32124
rect 8092 32122 8116 32124
rect 8172 32122 8196 32124
rect 8252 32122 8258 32124
rect 8012 32070 8014 32122
rect 8194 32070 8196 32122
rect 7950 32068 7956 32070
rect 8012 32068 8036 32070
rect 8092 32068 8116 32070
rect 8172 32068 8196 32070
rect 8252 32068 8258 32070
rect 7950 32059 8258 32068
rect 8312 31929 8340 32166
rect 8852 31952 8904 31958
rect 8298 31920 8354 31929
rect 8852 31894 8904 31900
rect 8298 31855 8354 31864
rect 7840 31816 7892 31822
rect 7840 31758 7892 31764
rect 8300 31680 8352 31686
rect 8864 31657 8892 31894
rect 8300 31622 8352 31628
rect 8850 31648 8906 31657
rect 7748 31476 7800 31482
rect 7748 31418 7800 31424
rect 8312 31385 8340 31622
rect 8850 31583 8906 31592
rect 8298 31376 8354 31385
rect 7656 31340 7708 31346
rect 8298 31311 8354 31320
rect 7656 31282 7708 31288
rect 7472 30116 7524 30122
rect 7472 30058 7524 30064
rect 7196 30048 7248 30054
rect 7196 29990 7248 29996
rect 7288 28484 7340 28490
rect 7288 28426 7340 28432
rect 7196 27396 7248 27402
rect 7196 27338 7248 27344
rect 7208 26042 7236 27338
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7300 24834 7328 28426
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 7380 26988 7432 26994
rect 7380 26930 7432 26936
rect 7392 26518 7420 26930
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7380 26512 7432 26518
rect 7380 26454 7432 26460
rect 7380 26308 7432 26314
rect 7380 26250 7432 26256
rect 7208 24806 7328 24834
rect 7104 24676 7156 24682
rect 7104 24618 7156 24624
rect 7102 24576 7158 24585
rect 7102 24511 7158 24520
rect 7116 24290 7144 24511
rect 7208 24410 7236 24806
rect 7286 24712 7342 24721
rect 7286 24647 7342 24656
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 7116 24262 7236 24290
rect 7012 24132 7064 24138
rect 7012 24074 7064 24080
rect 7104 24132 7156 24138
rect 7104 24074 7156 24080
rect 7024 24041 7052 24074
rect 7010 24032 7066 24041
rect 7010 23967 7066 23976
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 7024 22658 7052 23802
rect 6932 22630 7052 22658
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6932 21146 6960 22630
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6734 21040 6790 21049
rect 6734 20975 6790 20984
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6748 16153 6776 20878
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6734 16144 6790 16153
rect 6734 16079 6790 16088
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6840 12442 6868 20742
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6932 17218 6960 19994
rect 7024 17338 7052 22442
rect 7116 18426 7144 24074
rect 7208 23866 7236 24262
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7208 20058 7236 22986
rect 7300 22506 7328 24647
rect 7288 22500 7340 22506
rect 7288 22442 7340 22448
rect 7392 22234 7420 26250
rect 7484 24682 7512 26862
rect 7576 26586 7604 27406
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7564 25900 7616 25906
rect 7564 25842 7616 25848
rect 7472 24676 7524 24682
rect 7472 24618 7524 24624
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 7286 22128 7342 22137
rect 7286 22063 7342 22072
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7196 19916 7248 19922
rect 7196 19858 7248 19864
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 7102 17912 7158 17921
rect 7102 17847 7158 17856
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 6932 17190 7052 17218
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6932 14929 6960 17002
rect 6918 14920 6974 14929
rect 6918 14855 6974 14864
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6932 14618 6960 14758
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 7024 10810 7052 17190
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6932 9081 6960 9522
rect 7116 9450 7144 17847
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 6918 9072 6974 9081
rect 6918 9007 6974 9016
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8809 7144 8910
rect 7102 8800 7158 8809
rect 7102 8735 7158 8744
rect 7208 8090 7236 19858
rect 7300 18970 7328 22063
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7392 21690 7420 21966
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7392 18970 7420 21422
rect 7484 19514 7512 24346
rect 7576 20058 7604 25842
rect 7668 24857 7696 31282
rect 7930 31240 7986 31249
rect 7930 31175 7932 31184
rect 7984 31175 7986 31184
rect 7932 31146 7984 31152
rect 8300 31136 8352 31142
rect 8300 31078 8352 31084
rect 7950 31036 8258 31045
rect 7950 31034 7956 31036
rect 8012 31034 8036 31036
rect 8092 31034 8116 31036
rect 8172 31034 8196 31036
rect 8252 31034 8258 31036
rect 8012 30982 8014 31034
rect 8194 30982 8196 31034
rect 7950 30980 7956 30982
rect 8012 30980 8036 30982
rect 8092 30980 8116 30982
rect 8172 30980 8196 30982
rect 8252 30980 8258 30982
rect 7950 30971 8258 30980
rect 8312 30841 8340 31078
rect 8298 30832 8354 30841
rect 8298 30767 8354 30776
rect 7840 30592 7892 30598
rect 7932 30592 7984 30598
rect 7840 30534 7892 30540
rect 7930 30560 7932 30569
rect 8300 30592 8352 30598
rect 7984 30560 7986 30569
rect 7852 30258 7880 30534
rect 8300 30534 8352 30540
rect 7930 30495 7986 30504
rect 8312 30297 8340 30534
rect 8298 30288 8354 30297
rect 7840 30252 7892 30258
rect 8298 30223 8354 30232
rect 7840 30194 7892 30200
rect 9128 30184 9180 30190
rect 7930 30152 7986 30161
rect 9128 30126 9180 30132
rect 7930 30087 7932 30096
rect 7984 30087 7986 30096
rect 7932 30058 7984 30064
rect 7748 30048 7800 30054
rect 7748 29990 7800 29996
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 7760 29646 7788 29990
rect 7950 29948 8258 29957
rect 7950 29946 7956 29948
rect 8012 29946 8036 29948
rect 8092 29946 8116 29948
rect 8172 29946 8196 29948
rect 8252 29946 8258 29948
rect 8012 29894 8014 29946
rect 8194 29894 8196 29946
rect 7950 29892 7956 29894
rect 8012 29892 8036 29894
rect 8092 29892 8116 29894
rect 8172 29892 8196 29894
rect 8252 29892 8258 29894
rect 7950 29883 8258 29892
rect 8312 29753 8340 29990
rect 8298 29744 8354 29753
rect 8298 29679 8354 29688
rect 7748 29640 7800 29646
rect 7748 29582 7800 29588
rect 7932 29504 7984 29510
rect 7930 29472 7932 29481
rect 8300 29504 8352 29510
rect 7984 29472 7986 29481
rect 8300 29446 8352 29452
rect 7930 29407 7986 29416
rect 8312 29209 8340 29446
rect 8298 29200 8354 29209
rect 7840 29164 7892 29170
rect 8298 29135 8354 29144
rect 7840 29106 7892 29112
rect 7852 28762 7880 29106
rect 8944 29028 8996 29034
rect 8944 28970 8996 28976
rect 8300 28960 8352 28966
rect 8956 28937 8984 28970
rect 8300 28902 8352 28908
rect 8942 28928 8998 28937
rect 7950 28860 8258 28869
rect 7950 28858 7956 28860
rect 8012 28858 8036 28860
rect 8092 28858 8116 28860
rect 8172 28858 8196 28860
rect 8252 28858 8258 28860
rect 8012 28806 8014 28858
rect 8194 28806 8196 28858
rect 7950 28804 7956 28806
rect 8012 28804 8036 28806
rect 8092 28804 8116 28806
rect 8172 28804 8196 28806
rect 8252 28804 8258 28806
rect 7950 28795 8258 28804
rect 7840 28756 7892 28762
rect 7840 28698 7892 28704
rect 8312 28665 8340 28902
rect 8942 28863 8998 28872
rect 8298 28656 8354 28665
rect 8298 28591 8354 28600
rect 8668 28620 8720 28626
rect 8668 28562 8720 28568
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 7932 28416 7984 28422
rect 7930 28384 7932 28393
rect 7984 28384 7986 28393
rect 7930 28319 7986 28328
rect 8128 28218 8156 28494
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8116 28212 8168 28218
rect 8116 28154 8168 28160
rect 8312 28121 8340 28358
rect 8298 28112 8354 28121
rect 7748 28076 7800 28082
rect 7748 28018 7800 28024
rect 7840 28076 7892 28082
rect 8298 28047 8354 28056
rect 7840 28018 7892 28024
rect 7760 27674 7788 28018
rect 7748 27668 7800 27674
rect 7748 27610 7800 27616
rect 7852 27130 7880 28018
rect 7930 27976 7986 27985
rect 7930 27911 7932 27920
rect 7984 27911 7986 27920
rect 7932 27882 7984 27888
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 7950 27772 8258 27781
rect 7950 27770 7956 27772
rect 8012 27770 8036 27772
rect 8092 27770 8116 27772
rect 8172 27770 8196 27772
rect 8252 27770 8258 27772
rect 8012 27718 8014 27770
rect 8194 27718 8196 27770
rect 7950 27716 7956 27718
rect 8012 27716 8036 27718
rect 8092 27716 8116 27718
rect 8172 27716 8196 27718
rect 8252 27716 8258 27718
rect 7950 27707 8258 27716
rect 8312 27577 8340 27814
rect 8298 27568 8354 27577
rect 8298 27503 8354 27512
rect 7932 27328 7984 27334
rect 7930 27296 7932 27305
rect 8300 27328 8352 27334
rect 7984 27296 7986 27305
rect 8300 27270 8352 27276
rect 7930 27231 7986 27240
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 8312 27033 8340 27270
rect 8298 27024 8354 27033
rect 7748 26988 7800 26994
rect 8298 26959 8354 26968
rect 7748 26930 7800 26936
rect 7760 25498 7788 26930
rect 7930 26888 7986 26897
rect 7930 26823 7932 26832
rect 7984 26823 7986 26832
rect 7932 26794 7984 26800
rect 8300 26784 8352 26790
rect 8300 26726 8352 26732
rect 7950 26684 8258 26693
rect 7950 26682 7956 26684
rect 8012 26682 8036 26684
rect 8092 26682 8116 26684
rect 8172 26682 8196 26684
rect 8252 26682 8258 26684
rect 8012 26630 8014 26682
rect 8194 26630 8196 26682
rect 7950 26628 7956 26630
rect 8012 26628 8036 26630
rect 8092 26628 8116 26630
rect 8172 26628 8196 26630
rect 8252 26628 8258 26630
rect 7950 26619 8258 26628
rect 8312 26489 8340 26726
rect 8298 26480 8354 26489
rect 8298 26415 8354 26424
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8024 26376 8076 26382
rect 8022 26344 8024 26353
rect 8076 26344 8078 26353
rect 8022 26279 8078 26288
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8312 25945 8340 26182
rect 8484 25968 8536 25974
rect 8298 25936 8354 25945
rect 8484 25910 8536 25916
rect 8298 25871 8354 25880
rect 7930 25800 7986 25809
rect 7930 25735 7932 25744
rect 7984 25735 7986 25744
rect 7932 25706 7984 25712
rect 8300 25696 8352 25702
rect 8300 25638 8352 25644
rect 7950 25596 8258 25605
rect 7950 25594 7956 25596
rect 8012 25594 8036 25596
rect 8092 25594 8116 25596
rect 8172 25594 8196 25596
rect 8252 25594 8258 25596
rect 8012 25542 8014 25594
rect 8194 25542 8196 25594
rect 7950 25540 7956 25542
rect 8012 25540 8036 25542
rect 8092 25540 8116 25542
rect 8172 25540 8196 25542
rect 8252 25540 8258 25542
rect 7950 25531 8258 25540
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 8312 25401 8340 25638
rect 8298 25392 8354 25401
rect 8298 25327 8354 25336
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 7654 24848 7710 24857
rect 7654 24783 7710 24792
rect 7656 24744 7708 24750
rect 7656 24686 7708 24692
rect 7668 24410 7696 24686
rect 7656 24404 7708 24410
rect 7656 24346 7708 24352
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7668 22817 7696 23054
rect 7654 22808 7710 22817
rect 7654 22743 7656 22752
rect 7708 22743 7710 22752
rect 7656 22714 7708 22720
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7668 22166 7696 22578
rect 7656 22160 7708 22166
rect 7656 22102 7708 22108
rect 7760 21026 7788 25230
rect 7932 25152 7984 25158
rect 7930 25120 7932 25129
rect 8300 25152 8352 25158
rect 7984 25120 7986 25129
rect 8300 25094 8352 25100
rect 7930 25055 7986 25064
rect 8312 24857 8340 25094
rect 8298 24848 8354 24857
rect 7840 24812 7892 24818
rect 8298 24783 8354 24792
rect 7840 24754 7892 24760
rect 7852 24721 7880 24754
rect 7838 24712 7894 24721
rect 7838 24647 7894 24656
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7852 24313 7880 24550
rect 7950 24508 8258 24517
rect 7950 24506 7956 24508
rect 8012 24506 8036 24508
rect 8092 24506 8116 24508
rect 8172 24506 8196 24508
rect 8252 24506 8258 24508
rect 8012 24454 8014 24506
rect 8194 24454 8196 24506
rect 7950 24452 7956 24454
rect 8012 24452 8036 24454
rect 8092 24452 8116 24454
rect 8172 24452 8196 24454
rect 8252 24452 8258 24454
rect 7950 24443 8258 24452
rect 7838 24304 7894 24313
rect 7838 24239 7894 24248
rect 7932 24064 7984 24070
rect 8300 24064 8352 24070
rect 7932 24006 7984 24012
rect 8298 24032 8300 24041
rect 8352 24032 8354 24041
rect 7944 23769 7972 24006
rect 8298 23967 8354 23976
rect 7930 23760 7986 23769
rect 7840 23724 7892 23730
rect 7930 23695 7986 23704
rect 7840 23666 7892 23672
rect 7852 23322 7880 23666
rect 7950 23420 8258 23429
rect 7950 23418 7956 23420
rect 8012 23418 8036 23420
rect 8092 23418 8116 23420
rect 8172 23418 8196 23420
rect 8252 23418 8258 23420
rect 8012 23366 8014 23418
rect 8194 23366 8196 23418
rect 7950 23364 7956 23366
rect 8012 23364 8036 23366
rect 8092 23364 8116 23366
rect 8172 23364 8196 23366
rect 8252 23364 8258 23366
rect 7950 23355 8258 23364
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 7932 22976 7984 22982
rect 7932 22918 7984 22924
rect 7944 22681 7972 22918
rect 7930 22672 7986 22681
rect 7930 22607 7986 22616
rect 8128 22545 8156 23054
rect 8300 22976 8352 22982
rect 8298 22944 8300 22953
rect 8352 22944 8354 22953
rect 8298 22879 8354 22888
rect 8114 22536 8170 22545
rect 8114 22471 8170 22480
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7852 22137 7880 22374
rect 7950 22332 8258 22341
rect 7950 22330 7956 22332
rect 8012 22330 8036 22332
rect 8092 22330 8116 22332
rect 8172 22330 8196 22332
rect 8252 22330 8258 22332
rect 8012 22278 8014 22330
rect 8194 22278 8196 22330
rect 7950 22276 7956 22278
rect 8012 22276 8036 22278
rect 8092 22276 8116 22278
rect 8172 22276 8196 22278
rect 8252 22276 8258 22278
rect 7950 22267 8258 22276
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 8208 22160 8260 22166
rect 7838 22128 7894 22137
rect 8208 22102 8260 22108
rect 7838 22063 7894 22072
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7944 21593 7972 21830
rect 7930 21584 7986 21593
rect 7930 21519 7986 21528
rect 8036 21457 8064 21966
rect 8022 21448 8078 21457
rect 8220 21434 8248 22102
rect 8300 21888 8352 21894
rect 8298 21856 8300 21865
rect 8352 21856 8354 21865
rect 8298 21791 8354 21800
rect 8220 21406 8340 21434
rect 8022 21383 8078 21392
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7852 21049 7880 21286
rect 7950 21244 8258 21253
rect 7950 21242 7956 21244
rect 8012 21242 8036 21244
rect 8092 21242 8116 21244
rect 8172 21242 8196 21244
rect 8252 21242 8258 21244
rect 8012 21190 8014 21242
rect 8194 21190 8196 21242
rect 7950 21188 7956 21190
rect 8012 21188 8036 21190
rect 8092 21188 8116 21190
rect 8172 21188 8196 21190
rect 8252 21188 8258 21190
rect 7950 21179 8258 21188
rect 7668 20998 7788 21026
rect 7838 21040 7894 21049
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7576 19378 7604 19654
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7668 19258 7696 20998
rect 8312 21026 8340 21406
rect 7838 20975 7894 20984
rect 8220 20998 8340 21026
rect 7748 20936 7800 20942
rect 8116 20936 8168 20942
rect 7748 20878 7800 20884
rect 8114 20904 8116 20913
rect 8168 20904 8170 20913
rect 7760 20777 7788 20878
rect 8114 20839 8170 20848
rect 7746 20768 7802 20777
rect 7746 20703 7802 20712
rect 8220 20505 8248 20998
rect 8300 20800 8352 20806
rect 8298 20768 8300 20777
rect 8352 20768 8354 20777
rect 8298 20703 8354 20712
rect 8206 20496 8262 20505
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 8116 20460 8168 20466
rect 8206 20431 8262 20440
rect 8116 20402 8168 20408
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 7576 19230 7696 19258
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7300 18358 7328 18702
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7378 15464 7434 15473
rect 7378 15399 7434 15408
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7010 7984 7066 7993
rect 7010 7919 7066 7928
rect 7024 7886 7052 7919
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7194 7440 7250 7449
rect 7194 7375 7250 7384
rect 6734 6896 6790 6905
rect 6734 6831 6790 6840
rect 6366 5808 6422 5817
rect 6366 5743 6422 5752
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6380 3058 6408 5743
rect 6748 4622 6776 6831
rect 7208 6322 7236 7375
rect 7286 6624 7342 6633
rect 7286 6559 7342 6568
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 7300 4146 7328 6559
rect 7392 6458 7420 15399
rect 7484 14618 7512 19178
rect 7576 16250 7604 19230
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7562 14920 7618 14929
rect 7562 14855 7618 14864
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7576 14249 7604 14855
rect 7668 14521 7696 17614
rect 7654 14512 7710 14521
rect 7654 14447 7710 14456
rect 7562 14240 7618 14249
rect 7562 14175 7618 14184
rect 7654 9480 7710 9489
rect 7654 9415 7710 9424
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 5736 2094 5856 2122
rect 5828 56 5856 2094
rect 6276 468 6328 474
rect 6276 410 6328 416
rect 6288 56 6316 410
rect 6748 56 6776 3402
rect 7194 1184 7250 1193
rect 7194 1119 7250 1128
rect 7208 56 7236 1119
rect 7668 354 7696 9415
rect 7760 6662 7788 20402
rect 8128 20369 8156 20402
rect 8114 20360 8170 20369
rect 8404 20346 8432 22170
rect 8114 20295 8170 20304
rect 8312 20318 8432 20346
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7852 19961 7880 20198
rect 7950 20156 8258 20165
rect 7950 20154 7956 20156
rect 8012 20154 8036 20156
rect 8092 20154 8116 20156
rect 8172 20154 8196 20156
rect 8252 20154 8258 20156
rect 8012 20102 8014 20154
rect 8194 20102 8196 20154
rect 7950 20100 7956 20102
rect 8012 20100 8036 20102
rect 8092 20100 8116 20102
rect 8172 20100 8196 20102
rect 8252 20100 8258 20102
rect 7950 20091 8258 20100
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7838 19952 7894 19961
rect 7838 19887 7894 19896
rect 7944 19802 7972 19994
rect 8312 19938 8340 20318
rect 7852 19774 7972 19802
rect 8220 19910 8340 19938
rect 7852 15586 7880 19774
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7944 19417 7972 19654
rect 7930 19408 7986 19417
rect 7930 19343 7986 19352
rect 8220 19242 8248 19910
rect 8300 19712 8352 19718
rect 8298 19680 8300 19689
rect 8352 19680 8354 19689
rect 8298 19615 8354 19624
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 7950 19068 8258 19077
rect 7950 19066 7956 19068
rect 8012 19066 8036 19068
rect 8092 19066 8116 19068
rect 8172 19066 8196 19068
rect 8252 19066 8258 19068
rect 8012 19014 8014 19066
rect 8194 19014 8196 19066
rect 7950 19012 7956 19014
rect 8012 19012 8036 19014
rect 8092 19012 8116 19014
rect 8172 19012 8196 19014
rect 8252 19012 8258 19014
rect 7950 19003 8258 19012
rect 7932 18624 7984 18630
rect 8300 18624 8352 18630
rect 7932 18566 7984 18572
rect 8298 18592 8300 18601
rect 8352 18592 8354 18601
rect 7944 18329 7972 18566
rect 8298 18527 8354 18536
rect 7930 18320 7986 18329
rect 7930 18255 7986 18264
rect 7950 17980 8258 17989
rect 7950 17978 7956 17980
rect 8012 17978 8036 17980
rect 8092 17978 8116 17980
rect 8172 17978 8196 17980
rect 8252 17978 8258 17980
rect 8012 17926 8014 17978
rect 8194 17926 8196 17978
rect 7950 17924 7956 17926
rect 8012 17924 8036 17926
rect 8092 17924 8116 17926
rect 8172 17924 8196 17926
rect 8252 17924 8258 17926
rect 7950 17915 8258 17924
rect 8404 17785 8432 19246
rect 8390 17776 8446 17785
rect 8390 17711 8446 17720
rect 8390 17640 8446 17649
rect 8390 17575 8446 17584
rect 7950 16892 8258 16901
rect 7950 16890 7956 16892
rect 8012 16890 8036 16892
rect 8092 16890 8116 16892
rect 8172 16890 8196 16892
rect 8252 16890 8258 16892
rect 8012 16838 8014 16890
rect 8194 16838 8196 16890
rect 7950 16836 7956 16838
rect 8012 16836 8036 16838
rect 8092 16836 8116 16838
rect 8172 16836 8196 16838
rect 8252 16836 8258 16838
rect 7950 16827 8258 16836
rect 7950 15804 8258 15813
rect 7950 15802 7956 15804
rect 8012 15802 8036 15804
rect 8092 15802 8116 15804
rect 8172 15802 8196 15804
rect 8252 15802 8258 15804
rect 8012 15750 8014 15802
rect 8194 15750 8196 15802
rect 7950 15748 7956 15750
rect 8012 15748 8036 15750
rect 8092 15748 8116 15750
rect 8172 15748 8196 15750
rect 8252 15748 8258 15750
rect 7950 15739 8258 15748
rect 7852 15558 7972 15586
rect 7838 15464 7894 15473
rect 7838 15399 7894 15408
rect 7852 13530 7880 15399
rect 7944 14822 7972 15558
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7950 14716 8258 14725
rect 7950 14714 7956 14716
rect 8012 14714 8036 14716
rect 8092 14714 8116 14716
rect 8172 14714 8196 14716
rect 8252 14714 8258 14716
rect 8012 14662 8014 14714
rect 8194 14662 8196 14714
rect 7950 14660 7956 14662
rect 8012 14660 8036 14662
rect 8092 14660 8116 14662
rect 8172 14660 8196 14662
rect 8252 14660 8258 14662
rect 7950 14651 8258 14660
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 7950 13628 8258 13637
rect 7950 13626 7956 13628
rect 8012 13626 8036 13628
rect 8092 13626 8116 13628
rect 8172 13626 8196 13628
rect 8252 13626 8258 13628
rect 8012 13574 8014 13626
rect 8194 13574 8196 13626
rect 7950 13572 7956 13574
rect 8012 13572 8036 13574
rect 8092 13572 8116 13574
rect 8172 13572 8196 13574
rect 8252 13572 8258 13574
rect 7950 13563 8258 13572
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 8312 12889 8340 14282
rect 8298 12880 8354 12889
rect 8298 12815 8354 12824
rect 7950 12540 8258 12549
rect 7950 12538 7956 12540
rect 8012 12538 8036 12540
rect 8092 12538 8116 12540
rect 8172 12538 8196 12540
rect 8252 12538 8258 12540
rect 8012 12486 8014 12538
rect 8194 12486 8196 12538
rect 7950 12484 7956 12486
rect 8012 12484 8036 12486
rect 8092 12484 8116 12486
rect 8172 12484 8196 12486
rect 8252 12484 8258 12486
rect 7950 12475 8258 12484
rect 8404 11898 8432 17575
rect 8496 16574 8524 25910
rect 8588 20641 8616 26386
rect 8574 20632 8630 20641
rect 8574 20567 8630 20576
rect 8680 17513 8708 28562
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 8760 26512 8812 26518
rect 8760 26454 8812 26460
rect 8772 26217 8800 26454
rect 8758 26208 8814 26217
rect 8758 26143 8814 26152
rect 8852 23588 8904 23594
rect 8852 23530 8904 23536
rect 8864 23225 8892 23530
rect 8850 23216 8906 23225
rect 8850 23151 8906 23160
rect 8852 21072 8904 21078
rect 8852 21014 8904 21020
rect 8864 20505 8892 21014
rect 8850 20496 8906 20505
rect 8850 20431 8906 20440
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8772 18873 8800 19382
rect 8758 18864 8814 18873
rect 8758 18799 8814 18808
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8666 17504 8722 17513
rect 8666 17439 8722 17448
rect 8772 16574 8800 18226
rect 8956 18057 8984 27950
rect 9036 24608 9088 24614
rect 9034 24576 9036 24585
rect 9088 24576 9090 24585
rect 9034 24511 9090 24520
rect 9036 23520 9088 23526
rect 9034 23488 9036 23497
rect 9088 23488 9090 23497
rect 9034 23423 9090 23432
rect 9036 22432 9088 22438
rect 9034 22400 9036 22409
rect 9088 22400 9090 22409
rect 9034 22335 9090 22344
rect 9036 21344 9088 21350
rect 9034 21312 9036 21321
rect 9088 21312 9090 21321
rect 9034 21247 9090 21256
rect 9036 20256 9088 20262
rect 9034 20224 9036 20233
rect 9088 20224 9090 20233
rect 9034 20159 9090 20168
rect 9036 19508 9088 19514
rect 9036 19450 9088 19456
rect 9048 19145 9076 19450
rect 9034 19136 9090 19145
rect 9034 19071 9090 19080
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 8942 18048 8998 18057
rect 8942 17983 8998 17992
rect 8496 16546 8708 16574
rect 8772 16546 8892 16574
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8496 13161 8524 14962
rect 8588 13705 8616 15982
rect 8574 13696 8630 13705
rect 8574 13631 8630 13640
rect 8482 13152 8538 13161
rect 8482 13087 8538 13096
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 7950 11452 8258 11461
rect 7950 11450 7956 11452
rect 8012 11450 8036 11452
rect 8092 11450 8116 11452
rect 8172 11450 8196 11452
rect 8252 11450 8258 11452
rect 8012 11398 8014 11450
rect 8194 11398 8196 11450
rect 7950 11396 7956 11398
rect 8012 11396 8036 11398
rect 8092 11396 8116 11398
rect 8172 11396 8196 11398
rect 8252 11396 8258 11398
rect 7950 11387 8258 11396
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 7950 10364 8258 10373
rect 7950 10362 7956 10364
rect 8012 10362 8036 10364
rect 8092 10362 8116 10364
rect 8172 10362 8196 10364
rect 8252 10362 8258 10364
rect 8012 10310 8014 10362
rect 8194 10310 8196 10362
rect 7950 10308 7956 10310
rect 8012 10308 8036 10310
rect 8092 10308 8116 10310
rect 8172 10308 8196 10310
rect 8252 10308 8258 10310
rect 7950 10299 8258 10308
rect 8312 9625 8340 11086
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8298 9616 8354 9625
rect 8298 9551 8354 9560
rect 8404 9353 8432 10610
rect 8496 9897 8524 12106
rect 8680 11529 8708 16546
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8772 13433 8800 16050
rect 8864 14793 8892 16546
rect 9048 15065 9076 18294
rect 9140 16697 9168 30126
rect 9220 29708 9272 29714
rect 9220 29650 9272 29656
rect 9232 22094 9260 29650
rect 9496 29096 9548 29102
rect 9496 29038 9548 29044
rect 9312 25356 9364 25362
rect 9312 25298 9364 25304
rect 9324 22545 9352 25298
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 9310 22536 9366 22545
rect 9310 22471 9366 22480
rect 9232 22066 9352 22094
rect 9324 16969 9352 22066
rect 9310 16960 9366 16969
rect 9310 16895 9366 16904
rect 9126 16688 9182 16697
rect 9126 16623 9182 16632
rect 9034 15056 9090 15065
rect 9034 14991 9090 15000
rect 8850 14784 8906 14793
rect 8850 14719 8906 14728
rect 9416 13977 9444 24210
rect 9508 17241 9536 29038
rect 9588 24676 9640 24682
rect 9588 24618 9640 24624
rect 9494 17232 9550 17241
rect 9494 17167 9550 17176
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9402 13968 9458 13977
rect 9402 13903 9458 13912
rect 8758 13424 8814 13433
rect 8758 13359 8814 13368
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8772 12345 8800 13262
rect 9508 12617 9536 14350
rect 9494 12608 9550 12617
rect 9494 12543 9550 12552
rect 8758 12336 8814 12345
rect 8758 12271 8814 12280
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8666 11520 8722 11529
rect 8666 11455 8722 11464
rect 8772 10169 8800 12174
rect 9600 12073 9628 24618
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9586 12064 9642 12073
rect 9586 11999 9642 12008
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8956 10441 8984 11698
rect 8942 10432 8998 10441
rect 8942 10367 8998 10376
rect 8758 10160 8814 10169
rect 8758 10095 8814 10104
rect 8482 9888 8538 9897
rect 8482 9823 8538 9832
rect 8390 9344 8446 9353
rect 7950 9276 8258 9285
rect 8390 9279 8446 9288
rect 7950 9274 7956 9276
rect 8012 9274 8036 9276
rect 8092 9274 8116 9276
rect 8172 9274 8196 9276
rect 8252 9274 8258 9276
rect 8012 9222 8014 9274
rect 8194 9222 8196 9274
rect 7950 9220 7956 9222
rect 8012 9220 8036 9222
rect 8092 9220 8116 9222
rect 8172 9220 8196 9222
rect 8252 9220 8258 9222
rect 7950 9211 8258 9220
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 8265 8432 8434
rect 8390 8256 8446 8265
rect 7950 8188 8258 8197
rect 8390 8191 8446 8200
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 7838 7712 7894 7721
rect 7838 7647 7894 7656
rect 7852 6798 7880 7647
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 9692 6361 9720 18634
rect 9678 6352 9734 6361
rect 9678 6287 9734 6296
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7838 5536 7894 5545
rect 7838 5471 7894 5480
rect 7746 5264 7802 5273
rect 7746 5199 7802 5208
rect 7760 3058 7788 5199
rect 7852 3534 7880 5471
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 7668 326 7788 354
rect 7654 96 7710 105
rect 1596 54 1730 56
rect 1596 42 1624 54
rect 1412 14 1624 42
rect 1674 0 1730 54
rect 2134 0 2190 56
rect 2594 0 2650 56
rect 3054 0 3110 56
rect 3514 0 3570 56
rect 3974 0 4030 56
rect 4434 0 4490 56
rect 4894 0 4950 56
rect 5354 0 5410 56
rect 5814 0 5870 56
rect 6274 0 6330 56
rect 6734 0 6790 56
rect 7194 0 7250 56
rect 7654 0 7710 40
rect 7760 42 7788 326
rect 8036 56 8156 82
rect 8588 56 8616 2586
rect 9494 1320 9550 1329
rect 9494 1255 9550 1264
rect 9034 1048 9090 1057
rect 9034 983 9090 992
rect 9048 56 9076 983
rect 9508 56 9536 1255
rect 8036 54 8170 56
rect 8036 42 8064 54
rect 7760 14 8064 42
rect 8114 0 8170 54
rect 8574 0 8630 56
rect 9034 0 9090 56
rect 9494 0 9550 56
<< via2 >>
rect 3016 42458 3072 42460
rect 3096 42458 3152 42460
rect 3176 42458 3232 42460
rect 3256 42458 3312 42460
rect 3016 42406 3062 42458
rect 3062 42406 3072 42458
rect 3096 42406 3126 42458
rect 3126 42406 3138 42458
rect 3138 42406 3152 42458
rect 3176 42406 3190 42458
rect 3190 42406 3202 42458
rect 3202 42406 3232 42458
rect 3256 42406 3266 42458
rect 3266 42406 3312 42458
rect 3016 42404 3072 42406
rect 3096 42404 3152 42406
rect 3176 42404 3232 42406
rect 3256 42404 3312 42406
rect 7378 43560 7434 43616
rect 202 34040 258 34096
rect 110 31320 166 31376
rect 294 23160 350 23216
rect 202 5480 258 5536
rect 110 2760 166 2816
rect 1306 29960 1362 30016
rect 1306 28600 1362 28656
rect 1214 25880 1270 25936
rect 846 24520 902 24576
rect 938 20440 994 20496
rect 754 19080 810 19136
rect 1122 17720 1178 17776
rect 846 16360 902 16416
rect 754 15000 810 15056
rect 754 12280 810 12336
rect 1030 13640 1086 13696
rect 938 10920 994 10976
rect 570 9560 626 9616
rect 478 8200 534 8256
rect 386 4120 442 4176
rect 662 1400 718 1456
rect 1956 41914 2012 41916
rect 2036 41914 2092 41916
rect 2116 41914 2172 41916
rect 2196 41914 2252 41916
rect 1956 41862 2002 41914
rect 2002 41862 2012 41914
rect 2036 41862 2066 41914
rect 2066 41862 2078 41914
rect 2078 41862 2092 41914
rect 2116 41862 2130 41914
rect 2130 41862 2142 41914
rect 2142 41862 2172 41914
rect 2196 41862 2206 41914
rect 2206 41862 2252 41914
rect 1956 41860 2012 41862
rect 2036 41860 2092 41862
rect 2116 41860 2172 41862
rect 2196 41860 2252 41862
rect 1674 41656 1730 41712
rect 1674 41384 1730 41440
rect 1490 21800 1546 21856
rect 1956 40826 2012 40828
rect 2036 40826 2092 40828
rect 2116 40826 2172 40828
rect 2196 40826 2252 40828
rect 1956 40774 2002 40826
rect 2002 40774 2012 40826
rect 2036 40774 2066 40826
rect 2066 40774 2078 40826
rect 2078 40774 2092 40826
rect 2116 40774 2130 40826
rect 2130 40774 2142 40826
rect 2142 40774 2172 40826
rect 2196 40774 2206 40826
rect 2206 40774 2252 40826
rect 1956 40772 2012 40774
rect 2036 40772 2092 40774
rect 2116 40772 2172 40774
rect 2196 40772 2252 40774
rect 1956 39738 2012 39740
rect 2036 39738 2092 39740
rect 2116 39738 2172 39740
rect 2196 39738 2252 39740
rect 1956 39686 2002 39738
rect 2002 39686 2012 39738
rect 2036 39686 2066 39738
rect 2066 39686 2078 39738
rect 2078 39686 2092 39738
rect 2116 39686 2130 39738
rect 2130 39686 2142 39738
rect 2142 39686 2172 39738
rect 2196 39686 2206 39738
rect 2206 39686 2252 39738
rect 1956 39684 2012 39686
rect 2036 39684 2092 39686
rect 2116 39684 2172 39686
rect 2196 39684 2252 39686
rect 1956 38650 2012 38652
rect 2036 38650 2092 38652
rect 2116 38650 2172 38652
rect 2196 38650 2252 38652
rect 1956 38598 2002 38650
rect 2002 38598 2012 38650
rect 2036 38598 2066 38650
rect 2066 38598 2078 38650
rect 2078 38598 2092 38650
rect 2116 38598 2130 38650
rect 2130 38598 2142 38650
rect 2142 38598 2172 38650
rect 2196 38598 2206 38650
rect 2206 38598 2252 38650
rect 1956 38596 2012 38598
rect 2036 38596 2092 38598
rect 2116 38596 2172 38598
rect 2196 38596 2252 38598
rect 1956 37562 2012 37564
rect 2036 37562 2092 37564
rect 2116 37562 2172 37564
rect 2196 37562 2252 37564
rect 1956 37510 2002 37562
rect 2002 37510 2012 37562
rect 2036 37510 2066 37562
rect 2066 37510 2078 37562
rect 2078 37510 2092 37562
rect 2116 37510 2130 37562
rect 2130 37510 2142 37562
rect 2142 37510 2172 37562
rect 2196 37510 2206 37562
rect 2206 37510 2252 37562
rect 1956 37508 2012 37510
rect 2036 37508 2092 37510
rect 2116 37508 2172 37510
rect 2196 37508 2252 37510
rect 1956 36474 2012 36476
rect 2036 36474 2092 36476
rect 2116 36474 2172 36476
rect 2196 36474 2252 36476
rect 1956 36422 2002 36474
rect 2002 36422 2012 36474
rect 2036 36422 2066 36474
rect 2066 36422 2078 36474
rect 2078 36422 2092 36474
rect 2116 36422 2130 36474
rect 2130 36422 2142 36474
rect 2142 36422 2172 36474
rect 2196 36422 2206 36474
rect 2206 36422 2252 36474
rect 1956 36420 2012 36422
rect 2036 36420 2092 36422
rect 2116 36420 2172 36422
rect 2196 36420 2252 36422
rect 1956 35386 2012 35388
rect 2036 35386 2092 35388
rect 2116 35386 2172 35388
rect 2196 35386 2252 35388
rect 1956 35334 2002 35386
rect 2002 35334 2012 35386
rect 2036 35334 2066 35386
rect 2066 35334 2078 35386
rect 2078 35334 2092 35386
rect 2116 35334 2130 35386
rect 2130 35334 2142 35386
rect 2142 35334 2172 35386
rect 2196 35334 2206 35386
rect 2206 35334 2252 35386
rect 1956 35332 2012 35334
rect 2036 35332 2092 35334
rect 2116 35332 2172 35334
rect 2196 35332 2252 35334
rect 1956 34298 2012 34300
rect 2036 34298 2092 34300
rect 2116 34298 2172 34300
rect 2196 34298 2252 34300
rect 1956 34246 2002 34298
rect 2002 34246 2012 34298
rect 2036 34246 2066 34298
rect 2066 34246 2078 34298
rect 2078 34246 2092 34298
rect 2116 34246 2130 34298
rect 2130 34246 2142 34298
rect 2142 34246 2172 34298
rect 2196 34246 2206 34298
rect 2206 34246 2252 34298
rect 1956 34244 2012 34246
rect 2036 34244 2092 34246
rect 2116 34244 2172 34246
rect 2196 34244 2252 34246
rect 1956 33210 2012 33212
rect 2036 33210 2092 33212
rect 2116 33210 2172 33212
rect 2196 33210 2252 33212
rect 1956 33158 2002 33210
rect 2002 33158 2012 33210
rect 2036 33158 2066 33210
rect 2066 33158 2078 33210
rect 2078 33158 2092 33210
rect 2116 33158 2130 33210
rect 2130 33158 2142 33210
rect 2142 33158 2172 33210
rect 2196 33158 2206 33210
rect 2206 33158 2252 33210
rect 1956 33156 2012 33158
rect 2036 33156 2092 33158
rect 2116 33156 2172 33158
rect 2196 33156 2252 33158
rect 1956 32122 2012 32124
rect 2036 32122 2092 32124
rect 2116 32122 2172 32124
rect 2196 32122 2252 32124
rect 1956 32070 2002 32122
rect 2002 32070 2012 32122
rect 2036 32070 2066 32122
rect 2066 32070 2078 32122
rect 2078 32070 2092 32122
rect 2116 32070 2130 32122
rect 2130 32070 2142 32122
rect 2142 32070 2172 32122
rect 2196 32070 2206 32122
rect 2206 32070 2252 32122
rect 1956 32068 2012 32070
rect 2036 32068 2092 32070
rect 2116 32068 2172 32070
rect 2196 32068 2252 32070
rect 1956 31034 2012 31036
rect 2036 31034 2092 31036
rect 2116 31034 2172 31036
rect 2196 31034 2252 31036
rect 1956 30982 2002 31034
rect 2002 30982 2012 31034
rect 2036 30982 2066 31034
rect 2066 30982 2078 31034
rect 2078 30982 2092 31034
rect 2116 30982 2130 31034
rect 2130 30982 2142 31034
rect 2142 30982 2172 31034
rect 2196 30982 2206 31034
rect 2206 30982 2252 31034
rect 1956 30980 2012 30982
rect 2036 30980 2092 30982
rect 2116 30980 2172 30982
rect 2196 30980 2252 30982
rect 1956 29946 2012 29948
rect 2036 29946 2092 29948
rect 2116 29946 2172 29948
rect 2196 29946 2252 29948
rect 1956 29894 2002 29946
rect 2002 29894 2012 29946
rect 2036 29894 2066 29946
rect 2066 29894 2078 29946
rect 2078 29894 2092 29946
rect 2116 29894 2130 29946
rect 2130 29894 2142 29946
rect 2142 29894 2172 29946
rect 2196 29894 2206 29946
rect 2206 29894 2252 29946
rect 1956 29892 2012 29894
rect 2036 29892 2092 29894
rect 2116 29892 2172 29894
rect 2196 29892 2252 29894
rect 1956 28858 2012 28860
rect 2036 28858 2092 28860
rect 2116 28858 2172 28860
rect 2196 28858 2252 28860
rect 1956 28806 2002 28858
rect 2002 28806 2012 28858
rect 2036 28806 2066 28858
rect 2066 28806 2078 28858
rect 2078 28806 2092 28858
rect 2116 28806 2130 28858
rect 2130 28806 2142 28858
rect 2142 28806 2172 28858
rect 2196 28806 2206 28858
rect 2206 28806 2252 28858
rect 1956 28804 2012 28806
rect 2036 28804 2092 28806
rect 2116 28804 2172 28806
rect 2196 28804 2252 28806
rect 1956 27770 2012 27772
rect 2036 27770 2092 27772
rect 2116 27770 2172 27772
rect 2196 27770 2252 27772
rect 1956 27718 2002 27770
rect 2002 27718 2012 27770
rect 2036 27718 2066 27770
rect 2066 27718 2078 27770
rect 2078 27718 2092 27770
rect 2116 27718 2130 27770
rect 2130 27718 2142 27770
rect 2142 27718 2172 27770
rect 2196 27718 2206 27770
rect 2206 27718 2252 27770
rect 1956 27716 2012 27718
rect 2036 27716 2092 27718
rect 2116 27716 2172 27718
rect 2196 27716 2252 27718
rect 1956 26682 2012 26684
rect 2036 26682 2092 26684
rect 2116 26682 2172 26684
rect 2196 26682 2252 26684
rect 1956 26630 2002 26682
rect 2002 26630 2012 26682
rect 2036 26630 2066 26682
rect 2066 26630 2078 26682
rect 2078 26630 2092 26682
rect 2116 26630 2130 26682
rect 2130 26630 2142 26682
rect 2142 26630 2172 26682
rect 2196 26630 2206 26682
rect 2206 26630 2252 26682
rect 1956 26628 2012 26630
rect 2036 26628 2092 26630
rect 2116 26628 2172 26630
rect 2196 26628 2252 26630
rect 1956 25594 2012 25596
rect 2036 25594 2092 25596
rect 2116 25594 2172 25596
rect 2196 25594 2252 25596
rect 1956 25542 2002 25594
rect 2002 25542 2012 25594
rect 2036 25542 2066 25594
rect 2066 25542 2078 25594
rect 2078 25542 2092 25594
rect 2116 25542 2130 25594
rect 2130 25542 2142 25594
rect 2142 25542 2172 25594
rect 2196 25542 2206 25594
rect 2206 25542 2252 25594
rect 1956 25540 2012 25542
rect 2036 25540 2092 25542
rect 2116 25540 2172 25542
rect 2196 25540 2252 25542
rect 1956 24506 2012 24508
rect 2036 24506 2092 24508
rect 2116 24506 2172 24508
rect 2196 24506 2252 24508
rect 1956 24454 2002 24506
rect 2002 24454 2012 24506
rect 2036 24454 2066 24506
rect 2066 24454 2078 24506
rect 2078 24454 2092 24506
rect 2116 24454 2130 24506
rect 2130 24454 2142 24506
rect 2142 24454 2172 24506
rect 2196 24454 2206 24506
rect 2206 24454 2252 24506
rect 1956 24452 2012 24454
rect 2036 24452 2092 24454
rect 2116 24452 2172 24454
rect 2196 24452 2252 24454
rect 1956 23418 2012 23420
rect 2036 23418 2092 23420
rect 2116 23418 2172 23420
rect 2196 23418 2252 23420
rect 1956 23366 2002 23418
rect 2002 23366 2012 23418
rect 2036 23366 2066 23418
rect 2066 23366 2078 23418
rect 2078 23366 2092 23418
rect 2116 23366 2130 23418
rect 2130 23366 2142 23418
rect 2142 23366 2172 23418
rect 2196 23366 2206 23418
rect 2206 23366 2252 23418
rect 1956 23364 2012 23366
rect 2036 23364 2092 23366
rect 2116 23364 2172 23366
rect 2196 23364 2252 23366
rect 1956 22330 2012 22332
rect 2036 22330 2092 22332
rect 2116 22330 2172 22332
rect 2196 22330 2252 22332
rect 1956 22278 2002 22330
rect 2002 22278 2012 22330
rect 2036 22278 2066 22330
rect 2066 22278 2078 22330
rect 2078 22278 2092 22330
rect 2116 22278 2130 22330
rect 2130 22278 2142 22330
rect 2142 22278 2172 22330
rect 2196 22278 2206 22330
rect 2206 22278 2252 22330
rect 1956 22276 2012 22278
rect 2036 22276 2092 22278
rect 2116 22276 2172 22278
rect 2196 22276 2252 22278
rect 1956 21242 2012 21244
rect 2036 21242 2092 21244
rect 2116 21242 2172 21244
rect 2196 21242 2252 21244
rect 1956 21190 2002 21242
rect 2002 21190 2012 21242
rect 2036 21190 2066 21242
rect 2066 21190 2078 21242
rect 2078 21190 2092 21242
rect 2116 21190 2130 21242
rect 2130 21190 2142 21242
rect 2142 21190 2172 21242
rect 2196 21190 2206 21242
rect 2206 21190 2252 21242
rect 1956 21188 2012 21190
rect 2036 21188 2092 21190
rect 2116 21188 2172 21190
rect 2196 21188 2252 21190
rect 1956 20154 2012 20156
rect 2036 20154 2092 20156
rect 2116 20154 2172 20156
rect 2196 20154 2252 20156
rect 1956 20102 2002 20154
rect 2002 20102 2012 20154
rect 2036 20102 2066 20154
rect 2066 20102 2078 20154
rect 2078 20102 2092 20154
rect 2116 20102 2130 20154
rect 2130 20102 2142 20154
rect 2142 20102 2172 20154
rect 2196 20102 2206 20154
rect 2206 20102 2252 20154
rect 1956 20100 2012 20102
rect 2036 20100 2092 20102
rect 2116 20100 2172 20102
rect 2196 20100 2252 20102
rect 1956 19066 2012 19068
rect 2036 19066 2092 19068
rect 2116 19066 2172 19068
rect 2196 19066 2252 19068
rect 1956 19014 2002 19066
rect 2002 19014 2012 19066
rect 2036 19014 2066 19066
rect 2066 19014 2078 19066
rect 2078 19014 2092 19066
rect 2116 19014 2130 19066
rect 2130 19014 2142 19066
rect 2142 19014 2172 19066
rect 2196 19014 2206 19066
rect 2206 19014 2252 19066
rect 1956 19012 2012 19014
rect 2036 19012 2092 19014
rect 2116 19012 2172 19014
rect 2196 19012 2252 19014
rect 1956 17978 2012 17980
rect 2036 17978 2092 17980
rect 2116 17978 2172 17980
rect 2196 17978 2252 17980
rect 1956 17926 2002 17978
rect 2002 17926 2012 17978
rect 2036 17926 2066 17978
rect 2066 17926 2078 17978
rect 2078 17926 2092 17978
rect 2116 17926 2130 17978
rect 2130 17926 2142 17978
rect 2142 17926 2172 17978
rect 2196 17926 2206 17978
rect 2206 17926 2252 17978
rect 1956 17924 2012 17926
rect 2036 17924 2092 17926
rect 2116 17924 2172 17926
rect 2196 17924 2252 17926
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 1858 16244 1914 16280
rect 1858 16224 1860 16244
rect 1860 16224 1912 16244
rect 1912 16224 1914 16244
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 2410 27240 2466 27296
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 1858 13776 1914 13832
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 1858 11600 1914 11656
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 3016 41370 3072 41372
rect 3096 41370 3152 41372
rect 3176 41370 3232 41372
rect 3256 41370 3312 41372
rect 3016 41318 3062 41370
rect 3062 41318 3072 41370
rect 3096 41318 3126 41370
rect 3126 41318 3138 41370
rect 3138 41318 3152 41370
rect 3176 41318 3190 41370
rect 3190 41318 3202 41370
rect 3202 41318 3232 41370
rect 3256 41318 3266 41370
rect 3266 41318 3312 41370
rect 3016 41316 3072 41318
rect 3096 41316 3152 41318
rect 3176 41316 3232 41318
rect 3256 41316 3312 41318
rect 3016 40282 3072 40284
rect 3096 40282 3152 40284
rect 3176 40282 3232 40284
rect 3256 40282 3312 40284
rect 3016 40230 3062 40282
rect 3062 40230 3072 40282
rect 3096 40230 3126 40282
rect 3126 40230 3138 40282
rect 3138 40230 3152 40282
rect 3176 40230 3190 40282
rect 3190 40230 3202 40282
rect 3202 40230 3232 40282
rect 3256 40230 3266 40282
rect 3266 40230 3312 40282
rect 3016 40228 3072 40230
rect 3096 40228 3152 40230
rect 3176 40228 3232 40230
rect 3256 40228 3312 40230
rect 3016 39194 3072 39196
rect 3096 39194 3152 39196
rect 3176 39194 3232 39196
rect 3256 39194 3312 39196
rect 3016 39142 3062 39194
rect 3062 39142 3072 39194
rect 3096 39142 3126 39194
rect 3126 39142 3138 39194
rect 3138 39142 3152 39194
rect 3176 39142 3190 39194
rect 3190 39142 3202 39194
rect 3202 39142 3232 39194
rect 3256 39142 3266 39194
rect 3266 39142 3312 39194
rect 3016 39140 3072 39142
rect 3096 39140 3152 39142
rect 3176 39140 3232 39142
rect 3256 39140 3312 39142
rect 3016 38106 3072 38108
rect 3096 38106 3152 38108
rect 3176 38106 3232 38108
rect 3256 38106 3312 38108
rect 3016 38054 3062 38106
rect 3062 38054 3072 38106
rect 3096 38054 3126 38106
rect 3126 38054 3138 38106
rect 3138 38054 3152 38106
rect 3176 38054 3190 38106
rect 3190 38054 3202 38106
rect 3202 38054 3232 38106
rect 3256 38054 3266 38106
rect 3266 38054 3312 38106
rect 3016 38052 3072 38054
rect 3096 38052 3152 38054
rect 3176 38052 3232 38054
rect 3256 38052 3312 38054
rect 3016 37018 3072 37020
rect 3096 37018 3152 37020
rect 3176 37018 3232 37020
rect 3256 37018 3312 37020
rect 3016 36966 3062 37018
rect 3062 36966 3072 37018
rect 3096 36966 3126 37018
rect 3126 36966 3138 37018
rect 3138 36966 3152 37018
rect 3176 36966 3190 37018
rect 3190 36966 3202 37018
rect 3202 36966 3232 37018
rect 3256 36966 3266 37018
rect 3266 36966 3312 37018
rect 3016 36964 3072 36966
rect 3096 36964 3152 36966
rect 3176 36964 3232 36966
rect 3256 36964 3312 36966
rect 3016 35930 3072 35932
rect 3096 35930 3152 35932
rect 3176 35930 3232 35932
rect 3256 35930 3312 35932
rect 3016 35878 3062 35930
rect 3062 35878 3072 35930
rect 3096 35878 3126 35930
rect 3126 35878 3138 35930
rect 3138 35878 3152 35930
rect 3176 35878 3190 35930
rect 3190 35878 3202 35930
rect 3202 35878 3232 35930
rect 3256 35878 3266 35930
rect 3266 35878 3312 35930
rect 3016 35876 3072 35878
rect 3096 35876 3152 35878
rect 3176 35876 3232 35878
rect 3256 35876 3312 35878
rect 3016 34842 3072 34844
rect 3096 34842 3152 34844
rect 3176 34842 3232 34844
rect 3256 34842 3312 34844
rect 3016 34790 3062 34842
rect 3062 34790 3072 34842
rect 3096 34790 3126 34842
rect 3126 34790 3138 34842
rect 3138 34790 3152 34842
rect 3176 34790 3190 34842
rect 3190 34790 3202 34842
rect 3202 34790 3232 34842
rect 3256 34790 3266 34842
rect 3266 34790 3312 34842
rect 3016 34788 3072 34790
rect 3096 34788 3152 34790
rect 3176 34788 3232 34790
rect 3256 34788 3312 34790
rect 3016 33754 3072 33756
rect 3096 33754 3152 33756
rect 3176 33754 3232 33756
rect 3256 33754 3312 33756
rect 3016 33702 3062 33754
rect 3062 33702 3072 33754
rect 3096 33702 3126 33754
rect 3126 33702 3138 33754
rect 3138 33702 3152 33754
rect 3176 33702 3190 33754
rect 3190 33702 3202 33754
rect 3202 33702 3232 33754
rect 3256 33702 3266 33754
rect 3266 33702 3312 33754
rect 3016 33700 3072 33702
rect 3096 33700 3152 33702
rect 3176 33700 3232 33702
rect 3256 33700 3312 33702
rect 3016 32666 3072 32668
rect 3096 32666 3152 32668
rect 3176 32666 3232 32668
rect 3256 32666 3312 32668
rect 3016 32614 3062 32666
rect 3062 32614 3072 32666
rect 3096 32614 3126 32666
rect 3126 32614 3138 32666
rect 3138 32614 3152 32666
rect 3176 32614 3190 32666
rect 3190 32614 3202 32666
rect 3202 32614 3232 32666
rect 3256 32614 3266 32666
rect 3266 32614 3312 32666
rect 3016 32612 3072 32614
rect 3096 32612 3152 32614
rect 3176 32612 3232 32614
rect 3256 32612 3312 32614
rect 3016 31578 3072 31580
rect 3096 31578 3152 31580
rect 3176 31578 3232 31580
rect 3256 31578 3312 31580
rect 3016 31526 3062 31578
rect 3062 31526 3072 31578
rect 3096 31526 3126 31578
rect 3126 31526 3138 31578
rect 3138 31526 3152 31578
rect 3176 31526 3190 31578
rect 3190 31526 3202 31578
rect 3202 31526 3232 31578
rect 3256 31526 3266 31578
rect 3266 31526 3312 31578
rect 3016 31524 3072 31526
rect 3096 31524 3152 31526
rect 3176 31524 3232 31526
rect 3256 31524 3312 31526
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3016 30490 3072 30492
rect 3096 30490 3152 30492
rect 3176 30490 3232 30492
rect 3256 30490 3312 30492
rect 3016 30438 3062 30490
rect 3062 30438 3072 30490
rect 3096 30438 3126 30490
rect 3126 30438 3138 30490
rect 3138 30438 3152 30490
rect 3176 30438 3190 30490
rect 3190 30438 3202 30490
rect 3202 30438 3232 30490
rect 3256 30438 3266 30490
rect 3266 30438 3312 30490
rect 3016 30436 3072 30438
rect 3096 30436 3152 30438
rect 3176 30436 3232 30438
rect 3256 30436 3312 30438
rect 3016 29402 3072 29404
rect 3096 29402 3152 29404
rect 3176 29402 3232 29404
rect 3256 29402 3312 29404
rect 3016 29350 3062 29402
rect 3062 29350 3072 29402
rect 3096 29350 3126 29402
rect 3126 29350 3138 29402
rect 3138 29350 3152 29402
rect 3176 29350 3190 29402
rect 3190 29350 3202 29402
rect 3202 29350 3232 29402
rect 3256 29350 3266 29402
rect 3266 29350 3312 29402
rect 3016 29348 3072 29350
rect 3096 29348 3152 29350
rect 3176 29348 3232 29350
rect 3256 29348 3312 29350
rect 3016 28314 3072 28316
rect 3096 28314 3152 28316
rect 3176 28314 3232 28316
rect 3256 28314 3312 28316
rect 3016 28262 3062 28314
rect 3062 28262 3072 28314
rect 3096 28262 3126 28314
rect 3126 28262 3138 28314
rect 3138 28262 3152 28314
rect 3176 28262 3190 28314
rect 3190 28262 3202 28314
rect 3202 28262 3232 28314
rect 3256 28262 3266 28314
rect 3266 28262 3312 28314
rect 3016 28260 3072 28262
rect 3096 28260 3152 28262
rect 3176 28260 3232 28262
rect 3256 28260 3312 28262
rect 3016 27226 3072 27228
rect 3096 27226 3152 27228
rect 3176 27226 3232 27228
rect 3256 27226 3312 27228
rect 3016 27174 3062 27226
rect 3062 27174 3072 27226
rect 3096 27174 3126 27226
rect 3126 27174 3138 27226
rect 3138 27174 3152 27226
rect 3176 27174 3190 27226
rect 3190 27174 3202 27226
rect 3202 27174 3232 27226
rect 3256 27174 3266 27226
rect 3266 27174 3312 27226
rect 3016 27172 3072 27174
rect 3096 27172 3152 27174
rect 3176 27172 3232 27174
rect 3256 27172 3312 27174
rect 3016 26138 3072 26140
rect 3096 26138 3152 26140
rect 3176 26138 3232 26140
rect 3256 26138 3312 26140
rect 3016 26086 3062 26138
rect 3062 26086 3072 26138
rect 3096 26086 3126 26138
rect 3126 26086 3138 26138
rect 3138 26086 3152 26138
rect 3176 26086 3190 26138
rect 3190 26086 3202 26138
rect 3202 26086 3232 26138
rect 3256 26086 3266 26138
rect 3266 26086 3312 26138
rect 3016 26084 3072 26086
rect 3096 26084 3152 26086
rect 3176 26084 3232 26086
rect 3256 26084 3312 26086
rect 3054 25220 3110 25256
rect 3054 25200 3056 25220
rect 3056 25200 3108 25220
rect 3108 25200 3110 25220
rect 3016 25050 3072 25052
rect 3096 25050 3152 25052
rect 3176 25050 3232 25052
rect 3256 25050 3312 25052
rect 3016 24998 3062 25050
rect 3062 24998 3072 25050
rect 3096 24998 3126 25050
rect 3126 24998 3138 25050
rect 3138 24998 3152 25050
rect 3176 24998 3190 25050
rect 3190 24998 3202 25050
rect 3202 24998 3232 25050
rect 3256 24998 3266 25050
rect 3266 24998 3312 25050
rect 3016 24996 3072 24998
rect 3096 24996 3152 24998
rect 3176 24996 3232 24998
rect 3256 24996 3312 24998
rect 3016 23962 3072 23964
rect 3096 23962 3152 23964
rect 3176 23962 3232 23964
rect 3256 23962 3312 23964
rect 3016 23910 3062 23962
rect 3062 23910 3072 23962
rect 3096 23910 3126 23962
rect 3126 23910 3138 23962
rect 3138 23910 3152 23962
rect 3176 23910 3190 23962
rect 3190 23910 3202 23962
rect 3202 23910 3232 23962
rect 3256 23910 3266 23962
rect 3266 23910 3312 23962
rect 3016 23908 3072 23910
rect 3096 23908 3152 23910
rect 3176 23908 3232 23910
rect 3256 23908 3312 23910
rect 3016 22874 3072 22876
rect 3096 22874 3152 22876
rect 3176 22874 3232 22876
rect 3256 22874 3312 22876
rect 3016 22822 3062 22874
rect 3062 22822 3072 22874
rect 3096 22822 3126 22874
rect 3126 22822 3138 22874
rect 3138 22822 3152 22874
rect 3176 22822 3190 22874
rect 3190 22822 3202 22874
rect 3202 22822 3232 22874
rect 3256 22822 3266 22874
rect 3266 22822 3312 22874
rect 3016 22820 3072 22822
rect 3096 22820 3152 22822
rect 3176 22820 3232 22822
rect 3256 22820 3312 22822
rect 3016 21786 3072 21788
rect 3096 21786 3152 21788
rect 3176 21786 3232 21788
rect 3256 21786 3312 21788
rect 3016 21734 3062 21786
rect 3062 21734 3072 21786
rect 3096 21734 3126 21786
rect 3126 21734 3138 21786
rect 3138 21734 3152 21786
rect 3176 21734 3190 21786
rect 3190 21734 3202 21786
rect 3202 21734 3232 21786
rect 3256 21734 3266 21786
rect 3266 21734 3312 21786
rect 3016 21732 3072 21734
rect 3096 21732 3152 21734
rect 3176 21732 3232 21734
rect 3256 21732 3312 21734
rect 3016 20698 3072 20700
rect 3096 20698 3152 20700
rect 3176 20698 3232 20700
rect 3256 20698 3312 20700
rect 3016 20646 3062 20698
rect 3062 20646 3072 20698
rect 3096 20646 3126 20698
rect 3126 20646 3138 20698
rect 3138 20646 3152 20698
rect 3176 20646 3190 20698
rect 3190 20646 3202 20698
rect 3202 20646 3232 20698
rect 3256 20646 3266 20698
rect 3266 20646 3312 20698
rect 3016 20644 3072 20646
rect 3096 20644 3152 20646
rect 3176 20644 3232 20646
rect 3256 20644 3312 20646
rect 3016 19610 3072 19612
rect 3096 19610 3152 19612
rect 3176 19610 3232 19612
rect 3256 19610 3312 19612
rect 3016 19558 3062 19610
rect 3062 19558 3072 19610
rect 3096 19558 3126 19610
rect 3126 19558 3138 19610
rect 3138 19558 3152 19610
rect 3176 19558 3190 19610
rect 3190 19558 3202 19610
rect 3202 19558 3232 19610
rect 3256 19558 3266 19610
rect 3266 19558 3312 19610
rect 3016 19556 3072 19558
rect 3096 19556 3152 19558
rect 3176 19556 3232 19558
rect 3256 19556 3312 19558
rect 3514 19508 3570 19544
rect 3698 31728 3754 31784
rect 3698 23432 3754 23488
rect 3882 31728 3938 31784
rect 3514 19488 3516 19508
rect 3516 19488 3568 19508
rect 3568 19488 3570 19508
rect 3016 18522 3072 18524
rect 3096 18522 3152 18524
rect 3176 18522 3232 18524
rect 3256 18522 3312 18524
rect 3016 18470 3062 18522
rect 3062 18470 3072 18522
rect 3096 18470 3126 18522
rect 3126 18470 3138 18522
rect 3138 18470 3152 18522
rect 3176 18470 3190 18522
rect 3190 18470 3202 18522
rect 3202 18470 3232 18522
rect 3256 18470 3266 18522
rect 3266 18470 3312 18522
rect 3016 18468 3072 18470
rect 3096 18468 3152 18470
rect 3176 18468 3232 18470
rect 3256 18468 3312 18470
rect 3016 17434 3072 17436
rect 3096 17434 3152 17436
rect 3176 17434 3232 17436
rect 3256 17434 3312 17436
rect 3016 17382 3062 17434
rect 3062 17382 3072 17434
rect 3096 17382 3126 17434
rect 3126 17382 3138 17434
rect 3138 17382 3152 17434
rect 3176 17382 3190 17434
rect 3190 17382 3202 17434
rect 3202 17382 3232 17434
rect 3256 17382 3266 17434
rect 3266 17382 3312 17434
rect 3016 17380 3072 17382
rect 3096 17380 3152 17382
rect 3176 17380 3232 17382
rect 3256 17380 3312 17382
rect 3016 16346 3072 16348
rect 3096 16346 3152 16348
rect 3176 16346 3232 16348
rect 3256 16346 3312 16348
rect 3016 16294 3062 16346
rect 3062 16294 3072 16346
rect 3096 16294 3126 16346
rect 3126 16294 3138 16346
rect 3138 16294 3152 16346
rect 3176 16294 3190 16346
rect 3190 16294 3202 16346
rect 3202 16294 3232 16346
rect 3256 16294 3266 16346
rect 3266 16294 3312 16346
rect 3016 16292 3072 16294
rect 3096 16292 3152 16294
rect 3176 16292 3232 16294
rect 3256 16292 3312 16294
rect 3016 15258 3072 15260
rect 3096 15258 3152 15260
rect 3176 15258 3232 15260
rect 3256 15258 3312 15260
rect 3016 15206 3062 15258
rect 3062 15206 3072 15258
rect 3096 15206 3126 15258
rect 3126 15206 3138 15258
rect 3138 15206 3152 15258
rect 3176 15206 3190 15258
rect 3190 15206 3202 15258
rect 3202 15206 3232 15258
rect 3256 15206 3266 15258
rect 3266 15206 3312 15258
rect 3016 15204 3072 15206
rect 3096 15204 3152 15206
rect 3176 15204 3232 15206
rect 3256 15204 3312 15206
rect 3016 14170 3072 14172
rect 3096 14170 3152 14172
rect 3176 14170 3232 14172
rect 3256 14170 3312 14172
rect 3016 14118 3062 14170
rect 3062 14118 3072 14170
rect 3096 14118 3126 14170
rect 3126 14118 3138 14170
rect 3138 14118 3152 14170
rect 3176 14118 3190 14170
rect 3190 14118 3202 14170
rect 3202 14118 3232 14170
rect 3256 14118 3266 14170
rect 3266 14118 3312 14170
rect 3016 14116 3072 14118
rect 3096 14116 3152 14118
rect 3176 14116 3232 14118
rect 3256 14116 3312 14118
rect 3016 13082 3072 13084
rect 3096 13082 3152 13084
rect 3176 13082 3232 13084
rect 3256 13082 3312 13084
rect 3016 13030 3062 13082
rect 3062 13030 3072 13082
rect 3096 13030 3126 13082
rect 3126 13030 3138 13082
rect 3138 13030 3152 13082
rect 3176 13030 3190 13082
rect 3190 13030 3202 13082
rect 3202 13030 3232 13082
rect 3256 13030 3266 13082
rect 3266 13030 3312 13082
rect 3016 13028 3072 13030
rect 3096 13028 3152 13030
rect 3176 13028 3232 13030
rect 3256 13028 3312 13030
rect 3016 11994 3072 11996
rect 3096 11994 3152 11996
rect 3176 11994 3232 11996
rect 3256 11994 3312 11996
rect 3016 11942 3062 11994
rect 3062 11942 3072 11994
rect 3096 11942 3126 11994
rect 3126 11942 3138 11994
rect 3138 11942 3152 11994
rect 3176 11942 3190 11994
rect 3190 11942 3202 11994
rect 3202 11942 3232 11994
rect 3256 11942 3266 11994
rect 3266 11942 3312 11994
rect 3016 11940 3072 11942
rect 3096 11940 3152 11942
rect 3176 11940 3232 11942
rect 3256 11940 3312 11942
rect 2870 11056 2926 11112
rect 3016 10906 3072 10908
rect 3096 10906 3152 10908
rect 3176 10906 3232 10908
rect 3256 10906 3312 10908
rect 3016 10854 3062 10906
rect 3062 10854 3072 10906
rect 3096 10854 3126 10906
rect 3126 10854 3138 10906
rect 3138 10854 3152 10906
rect 3176 10854 3190 10906
rect 3190 10854 3202 10906
rect 3202 10854 3232 10906
rect 3256 10854 3266 10906
rect 3266 10854 3312 10906
rect 3016 10852 3072 10854
rect 3096 10852 3152 10854
rect 3176 10852 3232 10854
rect 3256 10852 3312 10854
rect 3016 9818 3072 9820
rect 3096 9818 3152 9820
rect 3176 9818 3232 9820
rect 3256 9818 3312 9820
rect 3016 9766 3062 9818
rect 3062 9766 3072 9818
rect 3096 9766 3126 9818
rect 3126 9766 3138 9818
rect 3138 9766 3152 9818
rect 3176 9766 3190 9818
rect 3190 9766 3202 9818
rect 3202 9766 3232 9818
rect 3256 9766 3266 9818
rect 3266 9766 3312 9818
rect 3016 9764 3072 9766
rect 3096 9764 3152 9766
rect 3176 9764 3232 9766
rect 3256 9764 3312 9766
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 2778 6840 2834 6896
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 3054 1264 3110 1320
rect 4526 29008 4582 29064
rect 4066 16088 4122 16144
rect 4986 41384 5042 41440
rect 4986 23468 4988 23488
rect 4988 23468 5040 23488
rect 5040 23468 5042 23488
rect 4986 23432 5042 23468
rect 4986 16360 5042 16416
rect 4894 16244 4950 16280
rect 4894 16224 4896 16244
rect 4896 16224 4948 16244
rect 4948 16224 4950 16244
rect 4618 8200 4674 8256
rect 5078 15544 5134 15600
rect 5538 39480 5594 39536
rect 5538 38292 5540 38312
rect 5540 38292 5592 38312
rect 5592 38292 5594 38312
rect 5538 38256 5594 38292
rect 6918 35536 6974 35592
rect 5998 11600 6054 11656
rect 5722 8200 5778 8256
rect 5814 7248 5870 7304
rect 5906 6160 5962 6216
rect 6182 13776 6238 13832
rect 6458 15408 6514 15464
rect 6734 23432 6790 23488
rect 7010 24928 7066 24984
rect 7470 42200 7526 42256
rect 7956 41914 8012 41916
rect 8036 41914 8092 41916
rect 8116 41914 8172 41916
rect 8196 41914 8252 41916
rect 7956 41862 8002 41914
rect 8002 41862 8012 41914
rect 8036 41862 8066 41914
rect 8066 41862 8078 41914
rect 8078 41862 8092 41914
rect 8116 41862 8130 41914
rect 8130 41862 8142 41914
rect 8142 41862 8172 41914
rect 8196 41862 8206 41914
rect 8206 41862 8252 41914
rect 7956 41860 8012 41862
rect 8036 41860 8092 41862
rect 8116 41860 8172 41862
rect 8196 41860 8252 41862
rect 7654 40568 7710 40624
rect 7956 40826 8012 40828
rect 8036 40826 8092 40828
rect 8116 40826 8172 40828
rect 8196 40826 8252 40828
rect 7956 40774 8002 40826
rect 8002 40774 8012 40826
rect 8036 40774 8066 40826
rect 8066 40774 8078 40826
rect 8078 40774 8092 40826
rect 8116 40774 8130 40826
rect 8130 40774 8142 40826
rect 8142 40774 8172 40826
rect 8196 40774 8206 40826
rect 8206 40774 8252 40826
rect 7956 40772 8012 40774
rect 8036 40772 8092 40774
rect 8116 40772 8172 40774
rect 8196 40772 8252 40774
rect 7930 39908 7986 39944
rect 7930 39888 7932 39908
rect 7932 39888 7984 39908
rect 7984 39888 7986 39908
rect 7956 39738 8012 39740
rect 8036 39738 8092 39740
rect 8116 39738 8172 39740
rect 8196 39738 8252 39740
rect 7956 39686 8002 39738
rect 8002 39686 8012 39738
rect 8036 39686 8066 39738
rect 8066 39686 8078 39738
rect 8078 39686 8092 39738
rect 8116 39686 8130 39738
rect 8130 39686 8142 39738
rect 8142 39686 8172 39738
rect 8196 39686 8206 39738
rect 8206 39686 8252 39738
rect 7956 39684 8012 39686
rect 8036 39684 8092 39686
rect 8116 39684 8172 39686
rect 8196 39684 8252 39686
rect 8298 39480 8354 39536
rect 7930 39244 7932 39264
rect 7932 39244 7984 39264
rect 7984 39244 7986 39264
rect 7930 39208 7986 39244
rect 8298 38936 8354 38992
rect 7470 36760 7526 36816
rect 7930 38820 7986 38856
rect 7930 38800 7932 38820
rect 7932 38800 7984 38820
rect 7984 38800 7986 38820
rect 7956 38650 8012 38652
rect 8036 38650 8092 38652
rect 8116 38650 8172 38652
rect 8196 38650 8252 38652
rect 7956 38598 8002 38650
rect 8002 38598 8012 38650
rect 8036 38598 8066 38650
rect 8066 38598 8078 38650
rect 8078 38598 8092 38650
rect 8116 38598 8130 38650
rect 8130 38598 8142 38650
rect 8142 38598 8172 38650
rect 8196 38598 8206 38650
rect 8206 38598 8252 38650
rect 7956 38596 8012 38598
rect 8036 38596 8092 38598
rect 8116 38596 8172 38598
rect 8196 38596 8252 38598
rect 8298 38392 8354 38448
rect 7930 38156 7932 38176
rect 7932 38156 7984 38176
rect 7984 38156 7986 38176
rect 7930 38120 7986 38156
rect 8298 37848 8354 37904
rect 7930 37732 7986 37768
rect 7930 37712 7932 37732
rect 7932 37712 7984 37732
rect 7984 37712 7986 37732
rect 7956 37562 8012 37564
rect 8036 37562 8092 37564
rect 8116 37562 8172 37564
rect 8196 37562 8252 37564
rect 7956 37510 8002 37562
rect 8002 37510 8012 37562
rect 8036 37510 8066 37562
rect 8066 37510 8078 37562
rect 8078 37510 8092 37562
rect 8116 37510 8130 37562
rect 8130 37510 8142 37562
rect 8142 37510 8172 37562
rect 8196 37510 8206 37562
rect 8206 37510 8252 37562
rect 7956 37508 8012 37510
rect 8036 37508 8092 37510
rect 8116 37508 8172 37510
rect 8196 37508 8252 37510
rect 8298 37304 8354 37360
rect 7930 37068 7932 37088
rect 7932 37068 7984 37088
rect 7984 37068 7986 37088
rect 7930 37032 7986 37068
rect 8298 36760 8354 36816
rect 7930 36644 7986 36680
rect 7930 36624 7932 36644
rect 7932 36624 7984 36644
rect 7984 36624 7986 36644
rect 7956 36474 8012 36476
rect 8036 36474 8092 36476
rect 8116 36474 8172 36476
rect 8196 36474 8252 36476
rect 7956 36422 8002 36474
rect 8002 36422 8012 36474
rect 8036 36422 8066 36474
rect 8066 36422 8078 36474
rect 8078 36422 8092 36474
rect 8116 36422 8130 36474
rect 8130 36422 8142 36474
rect 8142 36422 8172 36474
rect 8196 36422 8206 36474
rect 8206 36422 8252 36474
rect 7956 36420 8012 36422
rect 8036 36420 8092 36422
rect 8116 36420 8172 36422
rect 8196 36420 8252 36422
rect 8298 36216 8354 36272
rect 7930 35980 7932 36000
rect 7932 35980 7984 36000
rect 7984 35980 7986 36000
rect 7930 35944 7986 35980
rect 8298 35672 8354 35728
rect 7930 35556 7986 35592
rect 7930 35536 7932 35556
rect 7932 35536 7984 35556
rect 7984 35536 7986 35556
rect 7956 35386 8012 35388
rect 8036 35386 8092 35388
rect 8116 35386 8172 35388
rect 8196 35386 8252 35388
rect 7956 35334 8002 35386
rect 8002 35334 8012 35386
rect 8036 35334 8066 35386
rect 8066 35334 8078 35386
rect 8078 35334 8092 35386
rect 8116 35334 8130 35386
rect 8130 35334 8142 35386
rect 8142 35334 8172 35386
rect 8196 35334 8206 35386
rect 8206 35334 8252 35386
rect 7956 35332 8012 35334
rect 8036 35332 8092 35334
rect 8116 35332 8172 35334
rect 8196 35332 8252 35334
rect 8298 35128 8354 35184
rect 7930 34892 7932 34912
rect 7932 34892 7984 34912
rect 7984 34892 7986 34912
rect 7930 34856 7986 34892
rect 8298 34584 8354 34640
rect 7956 34298 8012 34300
rect 8036 34298 8092 34300
rect 8116 34298 8172 34300
rect 8196 34298 8252 34300
rect 7956 34246 8002 34298
rect 8002 34246 8012 34298
rect 8036 34246 8066 34298
rect 8066 34246 8078 34298
rect 8078 34246 8092 34298
rect 8116 34246 8130 34298
rect 8130 34246 8142 34298
rect 8142 34246 8172 34298
rect 8196 34246 8206 34298
rect 8206 34246 8252 34298
rect 7956 34244 8012 34246
rect 8036 34244 8092 34246
rect 8116 34244 8172 34246
rect 8196 34244 8252 34246
rect 8850 34312 8906 34368
rect 8298 34040 8354 34096
rect 7930 33804 7932 33824
rect 7932 33804 7984 33824
rect 7984 33804 7986 33824
rect 7930 33768 7986 33804
rect 8114 33496 8170 33552
rect 8298 33496 8354 33552
rect 7930 33380 7986 33416
rect 7930 33360 7932 33380
rect 7932 33360 7984 33380
rect 7984 33360 7986 33380
rect 7956 33210 8012 33212
rect 8036 33210 8092 33212
rect 8116 33210 8172 33212
rect 8196 33210 8252 33212
rect 7956 33158 8002 33210
rect 8002 33158 8012 33210
rect 8036 33158 8066 33210
rect 8066 33158 8078 33210
rect 8078 33158 8092 33210
rect 8116 33158 8130 33210
rect 8130 33158 8142 33210
rect 8142 33158 8172 33210
rect 8196 33158 8206 33210
rect 8206 33158 8252 33210
rect 7956 33156 8012 33158
rect 8036 33156 8092 33158
rect 8116 33156 8172 33158
rect 8196 33156 8252 33158
rect 8298 32952 8354 33008
rect 7470 32816 7526 32872
rect 7930 32716 7932 32736
rect 7932 32716 7984 32736
rect 7984 32716 7986 32736
rect 7930 32680 7986 32716
rect 8298 32408 8354 32464
rect 7930 32292 7986 32328
rect 7930 32272 7932 32292
rect 7932 32272 7984 32292
rect 7984 32272 7986 32292
rect 7956 32122 8012 32124
rect 8036 32122 8092 32124
rect 8116 32122 8172 32124
rect 8196 32122 8252 32124
rect 7956 32070 8002 32122
rect 8002 32070 8012 32122
rect 8036 32070 8066 32122
rect 8066 32070 8078 32122
rect 8078 32070 8092 32122
rect 8116 32070 8130 32122
rect 8130 32070 8142 32122
rect 8142 32070 8172 32122
rect 8196 32070 8206 32122
rect 8206 32070 8252 32122
rect 7956 32068 8012 32070
rect 8036 32068 8092 32070
rect 8116 32068 8172 32070
rect 8196 32068 8252 32070
rect 8298 31864 8354 31920
rect 8850 31592 8906 31648
rect 8298 31320 8354 31376
rect 7102 24520 7158 24576
rect 7286 24656 7342 24712
rect 7010 23976 7066 24032
rect 6734 20984 6790 21040
rect 6734 16088 6790 16144
rect 7286 22072 7342 22128
rect 7102 17856 7158 17912
rect 6918 14864 6974 14920
rect 6918 9016 6974 9072
rect 7102 8744 7158 8800
rect 7930 31204 7986 31240
rect 7930 31184 7932 31204
rect 7932 31184 7984 31204
rect 7984 31184 7986 31204
rect 7956 31034 8012 31036
rect 8036 31034 8092 31036
rect 8116 31034 8172 31036
rect 8196 31034 8252 31036
rect 7956 30982 8002 31034
rect 8002 30982 8012 31034
rect 8036 30982 8066 31034
rect 8066 30982 8078 31034
rect 8078 30982 8092 31034
rect 8116 30982 8130 31034
rect 8130 30982 8142 31034
rect 8142 30982 8172 31034
rect 8196 30982 8206 31034
rect 8206 30982 8252 31034
rect 7956 30980 8012 30982
rect 8036 30980 8092 30982
rect 8116 30980 8172 30982
rect 8196 30980 8252 30982
rect 8298 30776 8354 30832
rect 7930 30540 7932 30560
rect 7932 30540 7984 30560
rect 7984 30540 7986 30560
rect 7930 30504 7986 30540
rect 8298 30232 8354 30288
rect 7930 30116 7986 30152
rect 7930 30096 7932 30116
rect 7932 30096 7984 30116
rect 7984 30096 7986 30116
rect 7956 29946 8012 29948
rect 8036 29946 8092 29948
rect 8116 29946 8172 29948
rect 8196 29946 8252 29948
rect 7956 29894 8002 29946
rect 8002 29894 8012 29946
rect 8036 29894 8066 29946
rect 8066 29894 8078 29946
rect 8078 29894 8092 29946
rect 8116 29894 8130 29946
rect 8130 29894 8142 29946
rect 8142 29894 8172 29946
rect 8196 29894 8206 29946
rect 8206 29894 8252 29946
rect 7956 29892 8012 29894
rect 8036 29892 8092 29894
rect 8116 29892 8172 29894
rect 8196 29892 8252 29894
rect 8298 29688 8354 29744
rect 7930 29452 7932 29472
rect 7932 29452 7984 29472
rect 7984 29452 7986 29472
rect 7930 29416 7986 29452
rect 8298 29144 8354 29200
rect 7956 28858 8012 28860
rect 8036 28858 8092 28860
rect 8116 28858 8172 28860
rect 8196 28858 8252 28860
rect 7956 28806 8002 28858
rect 8002 28806 8012 28858
rect 8036 28806 8066 28858
rect 8066 28806 8078 28858
rect 8078 28806 8092 28858
rect 8116 28806 8130 28858
rect 8130 28806 8142 28858
rect 8142 28806 8172 28858
rect 8196 28806 8206 28858
rect 8206 28806 8252 28858
rect 7956 28804 8012 28806
rect 8036 28804 8092 28806
rect 8116 28804 8172 28806
rect 8196 28804 8252 28806
rect 8942 28872 8998 28928
rect 8298 28600 8354 28656
rect 7930 28364 7932 28384
rect 7932 28364 7984 28384
rect 7984 28364 7986 28384
rect 7930 28328 7986 28364
rect 8298 28056 8354 28112
rect 7930 27940 7986 27976
rect 7930 27920 7932 27940
rect 7932 27920 7984 27940
rect 7984 27920 7986 27940
rect 7956 27770 8012 27772
rect 8036 27770 8092 27772
rect 8116 27770 8172 27772
rect 8196 27770 8252 27772
rect 7956 27718 8002 27770
rect 8002 27718 8012 27770
rect 8036 27718 8066 27770
rect 8066 27718 8078 27770
rect 8078 27718 8092 27770
rect 8116 27718 8130 27770
rect 8130 27718 8142 27770
rect 8142 27718 8172 27770
rect 8196 27718 8206 27770
rect 8206 27718 8252 27770
rect 7956 27716 8012 27718
rect 8036 27716 8092 27718
rect 8116 27716 8172 27718
rect 8196 27716 8252 27718
rect 8298 27512 8354 27568
rect 7930 27276 7932 27296
rect 7932 27276 7984 27296
rect 7984 27276 7986 27296
rect 7930 27240 7986 27276
rect 8298 26968 8354 27024
rect 7930 26852 7986 26888
rect 7930 26832 7932 26852
rect 7932 26832 7984 26852
rect 7984 26832 7986 26852
rect 7956 26682 8012 26684
rect 8036 26682 8092 26684
rect 8116 26682 8172 26684
rect 8196 26682 8252 26684
rect 7956 26630 8002 26682
rect 8002 26630 8012 26682
rect 8036 26630 8066 26682
rect 8066 26630 8078 26682
rect 8078 26630 8092 26682
rect 8116 26630 8130 26682
rect 8130 26630 8142 26682
rect 8142 26630 8172 26682
rect 8196 26630 8206 26682
rect 8206 26630 8252 26682
rect 7956 26628 8012 26630
rect 8036 26628 8092 26630
rect 8116 26628 8172 26630
rect 8196 26628 8252 26630
rect 8298 26424 8354 26480
rect 8022 26324 8024 26344
rect 8024 26324 8076 26344
rect 8076 26324 8078 26344
rect 8022 26288 8078 26324
rect 8298 25880 8354 25936
rect 7930 25764 7986 25800
rect 7930 25744 7932 25764
rect 7932 25744 7984 25764
rect 7984 25744 7986 25764
rect 7956 25594 8012 25596
rect 8036 25594 8092 25596
rect 8116 25594 8172 25596
rect 8196 25594 8252 25596
rect 7956 25542 8002 25594
rect 8002 25542 8012 25594
rect 8036 25542 8066 25594
rect 8066 25542 8078 25594
rect 8078 25542 8092 25594
rect 8116 25542 8130 25594
rect 8130 25542 8142 25594
rect 8142 25542 8172 25594
rect 8196 25542 8206 25594
rect 8206 25542 8252 25594
rect 7956 25540 8012 25542
rect 8036 25540 8092 25542
rect 8116 25540 8172 25542
rect 8196 25540 8252 25542
rect 8298 25336 8354 25392
rect 7654 24792 7710 24848
rect 7654 22772 7710 22808
rect 7654 22752 7656 22772
rect 7656 22752 7708 22772
rect 7708 22752 7710 22772
rect 7930 25100 7932 25120
rect 7932 25100 7984 25120
rect 7984 25100 7986 25120
rect 7930 25064 7986 25100
rect 8298 24792 8354 24848
rect 7838 24656 7894 24712
rect 7956 24506 8012 24508
rect 8036 24506 8092 24508
rect 8116 24506 8172 24508
rect 8196 24506 8252 24508
rect 7956 24454 8002 24506
rect 8002 24454 8012 24506
rect 8036 24454 8066 24506
rect 8066 24454 8078 24506
rect 8078 24454 8092 24506
rect 8116 24454 8130 24506
rect 8130 24454 8142 24506
rect 8142 24454 8172 24506
rect 8196 24454 8206 24506
rect 8206 24454 8252 24506
rect 7956 24452 8012 24454
rect 8036 24452 8092 24454
rect 8116 24452 8172 24454
rect 8196 24452 8252 24454
rect 7838 24248 7894 24304
rect 8298 24012 8300 24032
rect 8300 24012 8352 24032
rect 8352 24012 8354 24032
rect 8298 23976 8354 24012
rect 7930 23704 7986 23760
rect 7956 23418 8012 23420
rect 8036 23418 8092 23420
rect 8116 23418 8172 23420
rect 8196 23418 8252 23420
rect 7956 23366 8002 23418
rect 8002 23366 8012 23418
rect 8036 23366 8066 23418
rect 8066 23366 8078 23418
rect 8078 23366 8092 23418
rect 8116 23366 8130 23418
rect 8130 23366 8142 23418
rect 8142 23366 8172 23418
rect 8196 23366 8206 23418
rect 8206 23366 8252 23418
rect 7956 23364 8012 23366
rect 8036 23364 8092 23366
rect 8116 23364 8172 23366
rect 8196 23364 8252 23366
rect 7930 22616 7986 22672
rect 8298 22924 8300 22944
rect 8300 22924 8352 22944
rect 8352 22924 8354 22944
rect 8298 22888 8354 22924
rect 8114 22480 8170 22536
rect 7956 22330 8012 22332
rect 8036 22330 8092 22332
rect 8116 22330 8172 22332
rect 8196 22330 8252 22332
rect 7956 22278 8002 22330
rect 8002 22278 8012 22330
rect 8036 22278 8066 22330
rect 8066 22278 8078 22330
rect 8078 22278 8092 22330
rect 8116 22278 8130 22330
rect 8130 22278 8142 22330
rect 8142 22278 8172 22330
rect 8196 22278 8206 22330
rect 8206 22278 8252 22330
rect 7956 22276 8012 22278
rect 8036 22276 8092 22278
rect 8116 22276 8172 22278
rect 8196 22276 8252 22278
rect 7838 22072 7894 22128
rect 7930 21528 7986 21584
rect 8022 21392 8078 21448
rect 8298 21836 8300 21856
rect 8300 21836 8352 21856
rect 8352 21836 8354 21856
rect 8298 21800 8354 21836
rect 7956 21242 8012 21244
rect 8036 21242 8092 21244
rect 8116 21242 8172 21244
rect 8196 21242 8252 21244
rect 7956 21190 8002 21242
rect 8002 21190 8012 21242
rect 8036 21190 8066 21242
rect 8066 21190 8078 21242
rect 8078 21190 8092 21242
rect 8116 21190 8130 21242
rect 8130 21190 8142 21242
rect 8142 21190 8172 21242
rect 8196 21190 8206 21242
rect 8206 21190 8252 21242
rect 7956 21188 8012 21190
rect 8036 21188 8092 21190
rect 8116 21188 8172 21190
rect 8196 21188 8252 21190
rect 7838 20984 7894 21040
rect 8114 20884 8116 20904
rect 8116 20884 8168 20904
rect 8168 20884 8170 20904
rect 8114 20848 8170 20884
rect 7746 20712 7802 20768
rect 8298 20748 8300 20768
rect 8300 20748 8352 20768
rect 8352 20748 8354 20768
rect 8298 20712 8354 20748
rect 8206 20440 8262 20496
rect 7378 15408 7434 15464
rect 7010 7928 7066 7984
rect 7194 7384 7250 7440
rect 6734 6840 6790 6896
rect 6366 5752 6422 5808
rect 7286 6568 7342 6624
rect 7562 14864 7618 14920
rect 7654 14456 7710 14512
rect 7562 14184 7618 14240
rect 7654 9424 7710 9480
rect 7194 1128 7250 1184
rect 8114 20304 8170 20360
rect 7956 20154 8012 20156
rect 8036 20154 8092 20156
rect 8116 20154 8172 20156
rect 8196 20154 8252 20156
rect 7956 20102 8002 20154
rect 8002 20102 8012 20154
rect 8036 20102 8066 20154
rect 8066 20102 8078 20154
rect 8078 20102 8092 20154
rect 8116 20102 8130 20154
rect 8130 20102 8142 20154
rect 8142 20102 8172 20154
rect 8196 20102 8206 20154
rect 8206 20102 8252 20154
rect 7956 20100 8012 20102
rect 8036 20100 8092 20102
rect 8116 20100 8172 20102
rect 8196 20100 8252 20102
rect 7838 19896 7894 19952
rect 7930 19352 7986 19408
rect 8298 19660 8300 19680
rect 8300 19660 8352 19680
rect 8352 19660 8354 19680
rect 8298 19624 8354 19660
rect 7956 19066 8012 19068
rect 8036 19066 8092 19068
rect 8116 19066 8172 19068
rect 8196 19066 8252 19068
rect 7956 19014 8002 19066
rect 8002 19014 8012 19066
rect 8036 19014 8066 19066
rect 8066 19014 8078 19066
rect 8078 19014 8092 19066
rect 8116 19014 8130 19066
rect 8130 19014 8142 19066
rect 8142 19014 8172 19066
rect 8196 19014 8206 19066
rect 8206 19014 8252 19066
rect 7956 19012 8012 19014
rect 8036 19012 8092 19014
rect 8116 19012 8172 19014
rect 8196 19012 8252 19014
rect 8298 18572 8300 18592
rect 8300 18572 8352 18592
rect 8352 18572 8354 18592
rect 8298 18536 8354 18572
rect 7930 18264 7986 18320
rect 7956 17978 8012 17980
rect 8036 17978 8092 17980
rect 8116 17978 8172 17980
rect 8196 17978 8252 17980
rect 7956 17926 8002 17978
rect 8002 17926 8012 17978
rect 8036 17926 8066 17978
rect 8066 17926 8078 17978
rect 8078 17926 8092 17978
rect 8116 17926 8130 17978
rect 8130 17926 8142 17978
rect 8142 17926 8172 17978
rect 8196 17926 8206 17978
rect 8206 17926 8252 17978
rect 7956 17924 8012 17926
rect 8036 17924 8092 17926
rect 8116 17924 8172 17926
rect 8196 17924 8252 17926
rect 8390 17720 8446 17776
rect 8390 17584 8446 17640
rect 7956 16890 8012 16892
rect 8036 16890 8092 16892
rect 8116 16890 8172 16892
rect 8196 16890 8252 16892
rect 7956 16838 8002 16890
rect 8002 16838 8012 16890
rect 8036 16838 8066 16890
rect 8066 16838 8078 16890
rect 8078 16838 8092 16890
rect 8116 16838 8130 16890
rect 8130 16838 8142 16890
rect 8142 16838 8172 16890
rect 8196 16838 8206 16890
rect 8206 16838 8252 16890
rect 7956 16836 8012 16838
rect 8036 16836 8092 16838
rect 8116 16836 8172 16838
rect 8196 16836 8252 16838
rect 7956 15802 8012 15804
rect 8036 15802 8092 15804
rect 8116 15802 8172 15804
rect 8196 15802 8252 15804
rect 7956 15750 8002 15802
rect 8002 15750 8012 15802
rect 8036 15750 8066 15802
rect 8066 15750 8078 15802
rect 8078 15750 8092 15802
rect 8116 15750 8130 15802
rect 8130 15750 8142 15802
rect 8142 15750 8172 15802
rect 8196 15750 8206 15802
rect 8206 15750 8252 15802
rect 7956 15748 8012 15750
rect 8036 15748 8092 15750
rect 8116 15748 8172 15750
rect 8196 15748 8252 15750
rect 7838 15408 7894 15464
rect 7956 14714 8012 14716
rect 8036 14714 8092 14716
rect 8116 14714 8172 14716
rect 8196 14714 8252 14716
rect 7956 14662 8002 14714
rect 8002 14662 8012 14714
rect 8036 14662 8066 14714
rect 8066 14662 8078 14714
rect 8078 14662 8092 14714
rect 8116 14662 8130 14714
rect 8130 14662 8142 14714
rect 8142 14662 8172 14714
rect 8196 14662 8206 14714
rect 8206 14662 8252 14714
rect 7956 14660 8012 14662
rect 8036 14660 8092 14662
rect 8116 14660 8172 14662
rect 8196 14660 8252 14662
rect 7956 13626 8012 13628
rect 8036 13626 8092 13628
rect 8116 13626 8172 13628
rect 8196 13626 8252 13628
rect 7956 13574 8002 13626
rect 8002 13574 8012 13626
rect 8036 13574 8066 13626
rect 8066 13574 8078 13626
rect 8078 13574 8092 13626
rect 8116 13574 8130 13626
rect 8130 13574 8142 13626
rect 8142 13574 8172 13626
rect 8196 13574 8206 13626
rect 8206 13574 8252 13626
rect 7956 13572 8012 13574
rect 8036 13572 8092 13574
rect 8116 13572 8172 13574
rect 8196 13572 8252 13574
rect 8298 12824 8354 12880
rect 7956 12538 8012 12540
rect 8036 12538 8092 12540
rect 8116 12538 8172 12540
rect 8196 12538 8252 12540
rect 7956 12486 8002 12538
rect 8002 12486 8012 12538
rect 8036 12486 8066 12538
rect 8066 12486 8078 12538
rect 8078 12486 8092 12538
rect 8116 12486 8130 12538
rect 8130 12486 8142 12538
rect 8142 12486 8172 12538
rect 8196 12486 8206 12538
rect 8206 12486 8252 12538
rect 7956 12484 8012 12486
rect 8036 12484 8092 12486
rect 8116 12484 8172 12486
rect 8196 12484 8252 12486
rect 8574 20576 8630 20632
rect 8758 26152 8814 26208
rect 8850 23160 8906 23216
rect 8850 20440 8906 20496
rect 8758 18808 8814 18864
rect 8666 17448 8722 17504
rect 9034 24556 9036 24576
rect 9036 24556 9088 24576
rect 9088 24556 9090 24576
rect 9034 24520 9090 24556
rect 9034 23468 9036 23488
rect 9036 23468 9088 23488
rect 9088 23468 9090 23488
rect 9034 23432 9090 23468
rect 9034 22380 9036 22400
rect 9036 22380 9088 22400
rect 9088 22380 9090 22400
rect 9034 22344 9090 22380
rect 9034 21292 9036 21312
rect 9036 21292 9088 21312
rect 9088 21292 9090 21312
rect 9034 21256 9090 21292
rect 9034 20204 9036 20224
rect 9036 20204 9088 20224
rect 9088 20204 9090 20224
rect 9034 20168 9090 20204
rect 9034 19080 9090 19136
rect 8942 17992 8998 18048
rect 8574 13640 8630 13696
rect 8482 13096 8538 13152
rect 7956 11450 8012 11452
rect 8036 11450 8092 11452
rect 8116 11450 8172 11452
rect 8196 11450 8252 11452
rect 7956 11398 8002 11450
rect 8002 11398 8012 11450
rect 8036 11398 8066 11450
rect 8066 11398 8078 11450
rect 8078 11398 8092 11450
rect 8116 11398 8130 11450
rect 8130 11398 8142 11450
rect 8142 11398 8172 11450
rect 8196 11398 8206 11450
rect 8206 11398 8252 11450
rect 7956 11396 8012 11398
rect 8036 11396 8092 11398
rect 8116 11396 8172 11398
rect 8196 11396 8252 11398
rect 7956 10362 8012 10364
rect 8036 10362 8092 10364
rect 8116 10362 8172 10364
rect 8196 10362 8252 10364
rect 7956 10310 8002 10362
rect 8002 10310 8012 10362
rect 8036 10310 8066 10362
rect 8066 10310 8078 10362
rect 8078 10310 8092 10362
rect 8116 10310 8130 10362
rect 8130 10310 8142 10362
rect 8142 10310 8172 10362
rect 8196 10310 8206 10362
rect 8206 10310 8252 10362
rect 7956 10308 8012 10310
rect 8036 10308 8092 10310
rect 8116 10308 8172 10310
rect 8196 10308 8252 10310
rect 8298 9560 8354 9616
rect 9310 22480 9366 22536
rect 9310 16904 9366 16960
rect 9126 16632 9182 16688
rect 9034 15000 9090 15056
rect 8850 14728 8906 14784
rect 9494 17176 9550 17232
rect 9402 13912 9458 13968
rect 8758 13368 8814 13424
rect 9494 12552 9550 12608
rect 8758 12280 8814 12336
rect 8666 11464 8722 11520
rect 9586 12008 9642 12064
rect 8942 10376 8998 10432
rect 8758 10104 8814 10160
rect 8482 9832 8538 9888
rect 8390 9288 8446 9344
rect 7956 9274 8012 9276
rect 8036 9274 8092 9276
rect 8116 9274 8172 9276
rect 8196 9274 8252 9276
rect 7956 9222 8002 9274
rect 8002 9222 8012 9274
rect 8036 9222 8066 9274
rect 8066 9222 8078 9274
rect 8078 9222 8092 9274
rect 8116 9222 8130 9274
rect 8130 9222 8142 9274
rect 8142 9222 8172 9274
rect 8196 9222 8206 9274
rect 8206 9222 8252 9274
rect 7956 9220 8012 9222
rect 8036 9220 8092 9222
rect 8116 9220 8172 9222
rect 8196 9220 8252 9222
rect 8390 8200 8446 8256
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7838 7656 7894 7712
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 9678 6296 9734 6352
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 7838 5480 7894 5536
rect 7746 5208 7802 5264
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 7654 40 7710 96
rect 9494 1264 9550 1320
rect 9034 992 9090 1048
<< metal3 >>
rect 0 43618 120 43648
rect 7373 43618 7439 43621
rect 0 43616 7439 43618
rect 0 43560 7378 43616
rect 7434 43560 7439 43616
rect 0 43558 7439 43560
rect 0 43528 120 43558
rect 7373 43555 7439 43558
rect 3006 42464 3322 42465
rect 3006 42400 3012 42464
rect 3076 42400 3092 42464
rect 3156 42400 3172 42464
rect 3236 42400 3252 42464
rect 3316 42400 3322 42464
rect 3006 42399 3322 42400
rect 0 42258 120 42288
rect 7465 42258 7531 42261
rect 0 42256 7531 42258
rect 0 42200 7470 42256
rect 7526 42200 7531 42256
rect 0 42198 7531 42200
rect 0 42168 120 42198
rect 7465 42195 7531 42198
rect 1946 41920 2262 41921
rect 1946 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2262 41920
rect 1946 41855 2262 41856
rect 7946 41920 8262 41921
rect 7946 41856 7952 41920
rect 8016 41856 8032 41920
rect 8096 41856 8112 41920
rect 8176 41856 8192 41920
rect 8256 41856 8262 41920
rect 7946 41855 8262 41856
rect 1526 41652 1532 41716
rect 1596 41714 1602 41716
rect 1669 41714 1735 41717
rect 1596 41712 1735 41714
rect 1596 41656 1674 41712
rect 1730 41656 1735 41712
rect 1596 41654 1735 41656
rect 1596 41652 1602 41654
rect 1669 41651 1735 41654
rect 1669 41444 1735 41445
rect 4981 41444 5047 41445
rect 1669 41440 1716 41444
rect 1780 41442 1786 41444
rect 1669 41384 1674 41440
rect 1669 41380 1716 41384
rect 1780 41382 1826 41442
rect 4981 41440 5028 41444
rect 5092 41442 5098 41444
rect 4981 41384 4986 41440
rect 1780 41380 1786 41382
rect 4981 41380 5028 41384
rect 5092 41382 5138 41442
rect 5092 41380 5098 41382
rect 1669 41379 1735 41380
rect 4981 41379 5047 41380
rect 3006 41376 3322 41377
rect 3006 41312 3012 41376
rect 3076 41312 3092 41376
rect 3156 41312 3172 41376
rect 3236 41312 3252 41376
rect 3316 41312 3322 41376
rect 3006 41311 3322 41312
rect 0 40898 120 40928
rect 0 40838 1778 40898
rect 0 40808 120 40838
rect 1718 40626 1778 40838
rect 1946 40832 2262 40833
rect 1946 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2262 40832
rect 1946 40767 2262 40768
rect 7946 40832 8262 40833
rect 7946 40768 7952 40832
rect 8016 40768 8032 40832
rect 8096 40768 8112 40832
rect 8176 40768 8192 40832
rect 8256 40768 8262 40832
rect 7946 40767 8262 40768
rect 7649 40626 7715 40629
rect 1718 40624 7715 40626
rect 1718 40568 7654 40624
rect 7710 40568 7715 40624
rect 1718 40566 7715 40568
rect 7649 40563 7715 40566
rect 3006 40288 3322 40289
rect 3006 40224 3012 40288
rect 3076 40224 3092 40288
rect 3156 40224 3172 40288
rect 3236 40224 3252 40288
rect 3316 40224 3322 40288
rect 3006 40223 3322 40224
rect 7925 39946 7991 39949
rect 7925 39944 8908 39946
rect 7925 39888 7930 39944
rect 7986 39888 8908 39944
rect 7925 39886 8908 39888
rect 7925 39883 7991 39886
rect 8848 39810 8908 39886
rect 9724 39810 9844 39840
rect 8848 39750 9844 39810
rect 1946 39744 2262 39745
rect 1946 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2262 39744
rect 1946 39679 2262 39680
rect 7946 39744 8262 39745
rect 7946 39680 7952 39744
rect 8016 39680 8032 39744
rect 8096 39680 8112 39744
rect 8176 39680 8192 39744
rect 8256 39680 8262 39744
rect 9724 39720 9844 39750
rect 7946 39679 8262 39680
rect 0 39538 120 39568
rect 5533 39538 5599 39541
rect 0 39536 5599 39538
rect 0 39480 5538 39536
rect 5594 39480 5599 39536
rect 0 39478 5599 39480
rect 0 39448 120 39478
rect 5533 39475 5599 39478
rect 8293 39538 8359 39541
rect 9724 39538 9844 39568
rect 8293 39536 9844 39538
rect 8293 39480 8298 39536
rect 8354 39480 9844 39536
rect 8293 39478 9844 39480
rect 8293 39475 8359 39478
rect 9724 39448 9844 39478
rect 7925 39266 7991 39269
rect 9724 39266 9844 39296
rect 7925 39264 9844 39266
rect 7925 39208 7930 39264
rect 7986 39208 9844 39264
rect 7925 39206 9844 39208
rect 7925 39203 7991 39206
rect 3006 39200 3322 39201
rect 3006 39136 3012 39200
rect 3076 39136 3092 39200
rect 3156 39136 3172 39200
rect 3236 39136 3252 39200
rect 3316 39136 3322 39200
rect 9724 39176 9844 39206
rect 3006 39135 3322 39136
rect 8293 38994 8359 38997
rect 9724 38994 9844 39024
rect 8293 38992 9844 38994
rect 8293 38936 8298 38992
rect 8354 38936 9844 38992
rect 8293 38934 9844 38936
rect 8293 38931 8359 38934
rect 9724 38904 9844 38934
rect 7925 38858 7991 38861
rect 7925 38856 8908 38858
rect 7925 38800 7930 38856
rect 7986 38800 8908 38856
rect 7925 38798 8908 38800
rect 7925 38795 7991 38798
rect 8848 38722 8908 38798
rect 9724 38722 9844 38752
rect 8848 38662 9844 38722
rect 1946 38656 2262 38657
rect 1946 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2262 38656
rect 1946 38591 2262 38592
rect 7946 38656 8262 38657
rect 7946 38592 7952 38656
rect 8016 38592 8032 38656
rect 8096 38592 8112 38656
rect 8176 38592 8192 38656
rect 8256 38592 8262 38656
rect 9724 38632 9844 38662
rect 7946 38591 8262 38592
rect 8293 38450 8359 38453
rect 9724 38450 9844 38480
rect 8293 38448 9844 38450
rect 8293 38392 8298 38448
rect 8354 38392 9844 38448
rect 8293 38390 9844 38392
rect 8293 38387 8359 38390
rect 9724 38360 9844 38390
rect 5533 38314 5599 38317
rect 2730 38312 5599 38314
rect 2730 38256 5538 38312
rect 5594 38256 5599 38312
rect 2730 38254 5599 38256
rect 0 38178 120 38208
rect 2730 38178 2790 38254
rect 5533 38251 5599 38254
rect 0 38118 2790 38178
rect 7925 38178 7991 38181
rect 9724 38178 9844 38208
rect 7925 38176 9844 38178
rect 7925 38120 7930 38176
rect 7986 38120 9844 38176
rect 7925 38118 9844 38120
rect 0 38088 120 38118
rect 7925 38115 7991 38118
rect 3006 38112 3322 38113
rect 3006 38048 3012 38112
rect 3076 38048 3092 38112
rect 3156 38048 3172 38112
rect 3236 38048 3252 38112
rect 3316 38048 3322 38112
rect 9724 38088 9844 38118
rect 3006 38047 3322 38048
rect 8293 37906 8359 37909
rect 9724 37906 9844 37936
rect 8293 37904 9844 37906
rect 8293 37848 8298 37904
rect 8354 37848 9844 37904
rect 8293 37846 9844 37848
rect 8293 37843 8359 37846
rect 9724 37816 9844 37846
rect 7925 37770 7991 37773
rect 7925 37768 8908 37770
rect 7925 37712 7930 37768
rect 7986 37712 8908 37768
rect 7925 37710 8908 37712
rect 7925 37707 7991 37710
rect 8848 37634 8908 37710
rect 9724 37634 9844 37664
rect 8848 37574 9844 37634
rect 1946 37568 2262 37569
rect 1946 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2262 37568
rect 1946 37503 2262 37504
rect 7946 37568 8262 37569
rect 7946 37504 7952 37568
rect 8016 37504 8032 37568
rect 8096 37504 8112 37568
rect 8176 37504 8192 37568
rect 8256 37504 8262 37568
rect 9724 37544 9844 37574
rect 7946 37503 8262 37504
rect 8293 37362 8359 37365
rect 9724 37362 9844 37392
rect 8293 37360 9844 37362
rect 8293 37304 8298 37360
rect 8354 37304 9844 37360
rect 8293 37302 9844 37304
rect 8293 37299 8359 37302
rect 9724 37272 9844 37302
rect 7925 37090 7991 37093
rect 9724 37090 9844 37120
rect 7925 37088 9844 37090
rect 7925 37032 7930 37088
rect 7986 37032 9844 37088
rect 7925 37030 9844 37032
rect 7925 37027 7991 37030
rect 3006 37024 3322 37025
rect 3006 36960 3012 37024
rect 3076 36960 3092 37024
rect 3156 36960 3172 37024
rect 3236 36960 3252 37024
rect 3316 36960 3322 37024
rect 9724 37000 9844 37030
rect 3006 36959 3322 36960
rect 0 36818 120 36848
rect 7465 36818 7531 36821
rect 0 36816 7531 36818
rect 0 36760 7470 36816
rect 7526 36760 7531 36816
rect 0 36758 7531 36760
rect 0 36728 120 36758
rect 7465 36755 7531 36758
rect 8293 36818 8359 36821
rect 9724 36818 9844 36848
rect 8293 36816 9844 36818
rect 8293 36760 8298 36816
rect 8354 36760 9844 36816
rect 8293 36758 9844 36760
rect 8293 36755 8359 36758
rect 9724 36728 9844 36758
rect 7925 36682 7991 36685
rect 7925 36680 8908 36682
rect 7925 36624 7930 36680
rect 7986 36624 8908 36680
rect 7925 36622 8908 36624
rect 7925 36619 7991 36622
rect 8848 36546 8908 36622
rect 9724 36546 9844 36576
rect 8848 36486 9844 36546
rect 1946 36480 2262 36481
rect 1946 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2262 36480
rect 1946 36415 2262 36416
rect 7946 36480 8262 36481
rect 7946 36416 7952 36480
rect 8016 36416 8032 36480
rect 8096 36416 8112 36480
rect 8176 36416 8192 36480
rect 8256 36416 8262 36480
rect 9724 36456 9844 36486
rect 7946 36415 8262 36416
rect 8293 36274 8359 36277
rect 9724 36274 9844 36304
rect 8293 36272 9844 36274
rect 8293 36216 8298 36272
rect 8354 36216 9844 36272
rect 8293 36214 9844 36216
rect 8293 36211 8359 36214
rect 9724 36184 9844 36214
rect 7925 36002 7991 36005
rect 9724 36002 9844 36032
rect 7925 36000 9844 36002
rect 7925 35944 7930 36000
rect 7986 35944 9844 36000
rect 7925 35942 9844 35944
rect 7925 35939 7991 35942
rect 3006 35936 3322 35937
rect 3006 35872 3012 35936
rect 3076 35872 3092 35936
rect 3156 35872 3172 35936
rect 3236 35872 3252 35936
rect 3316 35872 3322 35936
rect 9724 35912 9844 35942
rect 3006 35871 3322 35872
rect 8293 35730 8359 35733
rect 9724 35730 9844 35760
rect 8293 35728 9844 35730
rect 8293 35672 8298 35728
rect 8354 35672 9844 35728
rect 8293 35670 9844 35672
rect 8293 35667 8359 35670
rect 9724 35640 9844 35670
rect 6913 35594 6979 35597
rect 1718 35592 6979 35594
rect 1718 35536 6918 35592
rect 6974 35536 6979 35592
rect 1718 35534 6979 35536
rect 0 35458 120 35488
rect 1718 35458 1778 35534
rect 6913 35531 6979 35534
rect 7925 35594 7991 35597
rect 7925 35592 8908 35594
rect 7925 35536 7930 35592
rect 7986 35536 8908 35592
rect 7925 35534 8908 35536
rect 7925 35531 7991 35534
rect 0 35398 1778 35458
rect 8848 35458 8908 35534
rect 9724 35458 9844 35488
rect 8848 35398 9844 35458
rect 0 35368 120 35398
rect 1946 35392 2262 35393
rect 1946 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2262 35392
rect 1946 35327 2262 35328
rect 7946 35392 8262 35393
rect 7946 35328 7952 35392
rect 8016 35328 8032 35392
rect 8096 35328 8112 35392
rect 8176 35328 8192 35392
rect 8256 35328 8262 35392
rect 9724 35368 9844 35398
rect 7946 35327 8262 35328
rect 8293 35186 8359 35189
rect 9724 35186 9844 35216
rect 8293 35184 9844 35186
rect 8293 35128 8298 35184
rect 8354 35128 9844 35184
rect 8293 35126 9844 35128
rect 8293 35123 8359 35126
rect 9724 35096 9844 35126
rect 7925 34914 7991 34917
rect 9724 34914 9844 34944
rect 7925 34912 9844 34914
rect 7925 34856 7930 34912
rect 7986 34856 9844 34912
rect 7925 34854 9844 34856
rect 7925 34851 7991 34854
rect 3006 34848 3322 34849
rect 3006 34784 3012 34848
rect 3076 34784 3092 34848
rect 3156 34784 3172 34848
rect 3236 34784 3252 34848
rect 3316 34784 3322 34848
rect 9724 34824 9844 34854
rect 3006 34783 3322 34784
rect 8293 34642 8359 34645
rect 9724 34642 9844 34672
rect 8293 34640 9844 34642
rect 8293 34584 8298 34640
rect 8354 34584 9844 34640
rect 8293 34582 9844 34584
rect 8293 34579 8359 34582
rect 9724 34552 9844 34582
rect 8845 34370 8911 34373
rect 9724 34370 9844 34400
rect 8845 34368 9844 34370
rect 8845 34312 8850 34368
rect 8906 34312 9844 34368
rect 8845 34310 9844 34312
rect 8845 34307 8911 34310
rect 1946 34304 2262 34305
rect 1946 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2262 34304
rect 1946 34239 2262 34240
rect 7946 34304 8262 34305
rect 7946 34240 7952 34304
rect 8016 34240 8032 34304
rect 8096 34240 8112 34304
rect 8176 34240 8192 34304
rect 8256 34240 8262 34304
rect 9724 34280 9844 34310
rect 7946 34239 8262 34240
rect 0 34098 120 34128
rect 197 34098 263 34101
rect 0 34096 263 34098
rect 0 34040 202 34096
rect 258 34040 263 34096
rect 0 34038 263 34040
rect 0 34008 120 34038
rect 197 34035 263 34038
rect 8293 34098 8359 34101
rect 9724 34098 9844 34128
rect 8293 34096 9844 34098
rect 8293 34040 8298 34096
rect 8354 34040 9844 34096
rect 8293 34038 9844 34040
rect 8293 34035 8359 34038
rect 9724 34008 9844 34038
rect 7925 33826 7991 33829
rect 9724 33826 9844 33856
rect 7925 33824 9844 33826
rect 7925 33768 7930 33824
rect 7986 33768 9844 33824
rect 7925 33766 9844 33768
rect 7925 33763 7991 33766
rect 3006 33760 3322 33761
rect 3006 33696 3012 33760
rect 3076 33696 3092 33760
rect 3156 33696 3172 33760
rect 3236 33696 3252 33760
rect 3316 33696 3322 33760
rect 9724 33736 9844 33766
rect 3006 33695 3322 33696
rect 4654 33492 4660 33556
rect 4724 33554 4730 33556
rect 8109 33554 8175 33557
rect 4724 33552 8175 33554
rect 4724 33496 8114 33552
rect 8170 33496 8175 33552
rect 4724 33494 8175 33496
rect 4724 33492 4730 33494
rect 8109 33491 8175 33494
rect 8293 33554 8359 33557
rect 9724 33554 9844 33584
rect 8293 33552 9844 33554
rect 8293 33496 8298 33552
rect 8354 33496 9844 33552
rect 8293 33494 9844 33496
rect 8293 33491 8359 33494
rect 9724 33464 9844 33494
rect 7925 33418 7991 33421
rect 7925 33416 8908 33418
rect 7925 33360 7930 33416
rect 7986 33360 8908 33416
rect 7925 33358 8908 33360
rect 7925 33355 7991 33358
rect 8848 33282 8908 33358
rect 9724 33282 9844 33312
rect 8848 33222 9844 33282
rect 1946 33216 2262 33217
rect 1946 33152 1952 33216
rect 2016 33152 2032 33216
rect 2096 33152 2112 33216
rect 2176 33152 2192 33216
rect 2256 33152 2262 33216
rect 1946 33151 2262 33152
rect 7946 33216 8262 33217
rect 7946 33152 7952 33216
rect 8016 33152 8032 33216
rect 8096 33152 8112 33216
rect 8176 33152 8192 33216
rect 8256 33152 8262 33216
rect 9724 33192 9844 33222
rect 7946 33151 8262 33152
rect 8293 33010 8359 33013
rect 9724 33010 9844 33040
rect 8293 33008 9844 33010
rect 8293 32952 8298 33008
rect 8354 32952 9844 33008
rect 8293 32950 9844 32952
rect 8293 32947 8359 32950
rect 9724 32920 9844 32950
rect 7465 32874 7531 32877
rect 2730 32872 7531 32874
rect 2730 32816 7470 32872
rect 7526 32816 7531 32872
rect 2730 32814 7531 32816
rect 0 32738 120 32768
rect 2730 32738 2790 32814
rect 7465 32811 7531 32814
rect 0 32678 2790 32738
rect 7925 32738 7991 32741
rect 9724 32738 9844 32768
rect 7925 32736 9844 32738
rect 7925 32680 7930 32736
rect 7986 32680 9844 32736
rect 7925 32678 9844 32680
rect 0 32648 120 32678
rect 7925 32675 7991 32678
rect 3006 32672 3322 32673
rect 3006 32608 3012 32672
rect 3076 32608 3092 32672
rect 3156 32608 3172 32672
rect 3236 32608 3252 32672
rect 3316 32608 3322 32672
rect 9724 32648 9844 32678
rect 3006 32607 3322 32608
rect 8293 32466 8359 32469
rect 9724 32466 9844 32496
rect 8293 32464 9844 32466
rect 8293 32408 8298 32464
rect 8354 32408 9844 32464
rect 8293 32406 9844 32408
rect 8293 32403 8359 32406
rect 9724 32376 9844 32406
rect 7925 32330 7991 32333
rect 7925 32328 8908 32330
rect 7925 32272 7930 32328
rect 7986 32272 8908 32328
rect 7925 32270 8908 32272
rect 7925 32267 7991 32270
rect 8848 32194 8908 32270
rect 9724 32194 9844 32224
rect 8848 32134 9844 32194
rect 1946 32128 2262 32129
rect 1946 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2262 32128
rect 1946 32063 2262 32064
rect 7946 32128 8262 32129
rect 7946 32064 7952 32128
rect 8016 32064 8032 32128
rect 8096 32064 8112 32128
rect 8176 32064 8192 32128
rect 8256 32064 8262 32128
rect 9724 32104 9844 32134
rect 7946 32063 8262 32064
rect 8293 31922 8359 31925
rect 9724 31922 9844 31952
rect 8293 31920 9844 31922
rect 8293 31864 8298 31920
rect 8354 31864 9844 31920
rect 8293 31862 9844 31864
rect 8293 31859 8359 31862
rect 9724 31832 9844 31862
rect 3693 31786 3759 31789
rect 3877 31786 3943 31789
rect 3693 31784 3943 31786
rect 3693 31728 3698 31784
rect 3754 31728 3882 31784
rect 3938 31728 3943 31784
rect 3693 31726 3943 31728
rect 3693 31723 3759 31726
rect 3877 31723 3943 31726
rect 8845 31650 8911 31653
rect 9724 31650 9844 31680
rect 8845 31648 9844 31650
rect 8845 31592 8850 31648
rect 8906 31592 9844 31648
rect 8845 31590 9844 31592
rect 8845 31587 8911 31590
rect 3006 31584 3322 31585
rect 3006 31520 3012 31584
rect 3076 31520 3092 31584
rect 3156 31520 3172 31584
rect 3236 31520 3252 31584
rect 3316 31520 3322 31584
rect 9724 31560 9844 31590
rect 3006 31519 3322 31520
rect 0 31381 120 31408
rect 0 31376 171 31381
rect 0 31320 110 31376
rect 166 31320 171 31376
rect 0 31315 171 31320
rect 8293 31378 8359 31381
rect 9724 31378 9844 31408
rect 8293 31376 9844 31378
rect 8293 31320 8298 31376
rect 8354 31320 9844 31376
rect 8293 31318 9844 31320
rect 8293 31315 8359 31318
rect 0 31288 120 31315
rect 9724 31288 9844 31318
rect 7925 31242 7991 31245
rect 7925 31240 8908 31242
rect 7925 31184 7930 31240
rect 7986 31184 8908 31240
rect 7925 31182 8908 31184
rect 7925 31179 7991 31182
rect 8848 31106 8908 31182
rect 9724 31106 9844 31136
rect 8848 31046 9844 31106
rect 1946 31040 2262 31041
rect 1946 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2262 31040
rect 1946 30975 2262 30976
rect 7946 31040 8262 31041
rect 7946 30976 7952 31040
rect 8016 30976 8032 31040
rect 8096 30976 8112 31040
rect 8176 30976 8192 31040
rect 8256 30976 8262 31040
rect 9724 31016 9844 31046
rect 7946 30975 8262 30976
rect 8293 30834 8359 30837
rect 9724 30834 9844 30864
rect 8293 30832 9844 30834
rect 8293 30776 8298 30832
rect 8354 30776 9844 30832
rect 8293 30774 9844 30776
rect 8293 30771 8359 30774
rect 9724 30744 9844 30774
rect 7925 30562 7991 30565
rect 9724 30562 9844 30592
rect 7925 30560 9844 30562
rect 7925 30504 7930 30560
rect 7986 30504 9844 30560
rect 7925 30502 9844 30504
rect 7925 30499 7991 30502
rect 3006 30496 3322 30497
rect 3006 30432 3012 30496
rect 3076 30432 3092 30496
rect 3156 30432 3172 30496
rect 3236 30432 3252 30496
rect 3316 30432 3322 30496
rect 9724 30472 9844 30502
rect 3006 30431 3322 30432
rect 8293 30290 8359 30293
rect 9724 30290 9844 30320
rect 8293 30288 9844 30290
rect 8293 30232 8298 30288
rect 8354 30232 9844 30288
rect 8293 30230 9844 30232
rect 8293 30227 8359 30230
rect 9724 30200 9844 30230
rect 7925 30154 7991 30157
rect 7925 30152 8908 30154
rect 7925 30096 7930 30152
rect 7986 30096 8908 30152
rect 7925 30094 8908 30096
rect 7925 30091 7991 30094
rect 0 30018 120 30048
rect 1301 30018 1367 30021
rect 0 30016 1367 30018
rect 0 29960 1306 30016
rect 1362 29960 1367 30016
rect 0 29958 1367 29960
rect 8848 30018 8908 30094
rect 9724 30018 9844 30048
rect 8848 29958 9844 30018
rect 0 29928 120 29958
rect 1301 29955 1367 29958
rect 1946 29952 2262 29953
rect 1946 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2262 29952
rect 1946 29887 2262 29888
rect 7946 29952 8262 29953
rect 7946 29888 7952 29952
rect 8016 29888 8032 29952
rect 8096 29888 8112 29952
rect 8176 29888 8192 29952
rect 8256 29888 8262 29952
rect 9724 29928 9844 29958
rect 7946 29887 8262 29888
rect 8293 29746 8359 29749
rect 9724 29746 9844 29776
rect 8293 29744 9844 29746
rect 8293 29688 8298 29744
rect 8354 29688 9844 29744
rect 8293 29686 9844 29688
rect 8293 29683 8359 29686
rect 9724 29656 9844 29686
rect 7925 29474 7991 29477
rect 9724 29474 9844 29504
rect 7925 29472 9844 29474
rect 7925 29416 7930 29472
rect 7986 29416 9844 29472
rect 7925 29414 9844 29416
rect 7925 29411 7991 29414
rect 3006 29408 3322 29409
rect 3006 29344 3012 29408
rect 3076 29344 3092 29408
rect 3156 29344 3172 29408
rect 3236 29344 3252 29408
rect 3316 29344 3322 29408
rect 9724 29384 9844 29414
rect 3006 29343 3322 29344
rect 8293 29202 8359 29205
rect 9724 29202 9844 29232
rect 8293 29200 9844 29202
rect 8293 29144 8298 29200
rect 8354 29144 9844 29200
rect 8293 29142 9844 29144
rect 8293 29139 8359 29142
rect 9724 29112 9844 29142
rect 3918 29004 3924 29068
rect 3988 29066 3994 29068
rect 4521 29066 4587 29069
rect 3988 29064 4587 29066
rect 3988 29008 4526 29064
rect 4582 29008 4587 29064
rect 3988 29006 4587 29008
rect 3988 29004 3994 29006
rect 4521 29003 4587 29006
rect 8937 28930 9003 28933
rect 9724 28930 9844 28960
rect 8937 28928 9844 28930
rect 8937 28872 8942 28928
rect 8998 28872 9844 28928
rect 8937 28870 9844 28872
rect 8937 28867 9003 28870
rect 1946 28864 2262 28865
rect 1946 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2262 28864
rect 1946 28799 2262 28800
rect 7946 28864 8262 28865
rect 7946 28800 7952 28864
rect 8016 28800 8032 28864
rect 8096 28800 8112 28864
rect 8176 28800 8192 28864
rect 8256 28800 8262 28864
rect 9724 28840 9844 28870
rect 7946 28799 8262 28800
rect 0 28658 120 28688
rect 1301 28658 1367 28661
rect 0 28656 1367 28658
rect 0 28600 1306 28656
rect 1362 28600 1367 28656
rect 0 28598 1367 28600
rect 0 28568 120 28598
rect 1301 28595 1367 28598
rect 8293 28658 8359 28661
rect 9724 28658 9844 28688
rect 8293 28656 9844 28658
rect 8293 28600 8298 28656
rect 8354 28600 9844 28656
rect 8293 28598 9844 28600
rect 8293 28595 8359 28598
rect 9724 28568 9844 28598
rect 7925 28386 7991 28389
rect 9724 28386 9844 28416
rect 7925 28384 9844 28386
rect 7925 28328 7930 28384
rect 7986 28328 9844 28384
rect 7925 28326 9844 28328
rect 7925 28323 7991 28326
rect 3006 28320 3322 28321
rect 3006 28256 3012 28320
rect 3076 28256 3092 28320
rect 3156 28256 3172 28320
rect 3236 28256 3252 28320
rect 3316 28256 3322 28320
rect 9724 28296 9844 28326
rect 3006 28255 3322 28256
rect 8293 28114 8359 28117
rect 9724 28114 9844 28144
rect 8293 28112 9844 28114
rect 8293 28056 8298 28112
rect 8354 28056 9844 28112
rect 8293 28054 9844 28056
rect 8293 28051 8359 28054
rect 9724 28024 9844 28054
rect 7925 27978 7991 27981
rect 7925 27976 8908 27978
rect 7925 27920 7930 27976
rect 7986 27920 8908 27976
rect 7925 27918 8908 27920
rect 7925 27915 7991 27918
rect 8848 27842 8908 27918
rect 9724 27842 9844 27872
rect 8848 27782 9844 27842
rect 1946 27776 2262 27777
rect 1946 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2262 27776
rect 1946 27711 2262 27712
rect 7946 27776 8262 27777
rect 7946 27712 7952 27776
rect 8016 27712 8032 27776
rect 8096 27712 8112 27776
rect 8176 27712 8192 27776
rect 8256 27712 8262 27776
rect 9724 27752 9844 27782
rect 7946 27711 8262 27712
rect 8293 27570 8359 27573
rect 9724 27570 9844 27600
rect 8293 27568 9844 27570
rect 8293 27512 8298 27568
rect 8354 27512 9844 27568
rect 8293 27510 9844 27512
rect 8293 27507 8359 27510
rect 9724 27480 9844 27510
rect 0 27298 120 27328
rect 2405 27298 2471 27301
rect 0 27296 2471 27298
rect 0 27240 2410 27296
rect 2466 27240 2471 27296
rect 0 27238 2471 27240
rect 0 27208 120 27238
rect 2405 27235 2471 27238
rect 7925 27298 7991 27301
rect 9724 27298 9844 27328
rect 7925 27296 9844 27298
rect 7925 27240 7930 27296
rect 7986 27240 9844 27296
rect 7925 27238 9844 27240
rect 7925 27235 7991 27238
rect 3006 27232 3322 27233
rect 3006 27168 3012 27232
rect 3076 27168 3092 27232
rect 3156 27168 3172 27232
rect 3236 27168 3252 27232
rect 3316 27168 3322 27232
rect 9724 27208 9844 27238
rect 3006 27167 3322 27168
rect 8293 27026 8359 27029
rect 9724 27026 9844 27056
rect 8293 27024 9844 27026
rect 8293 26968 8298 27024
rect 8354 26968 9844 27024
rect 8293 26966 9844 26968
rect 8293 26963 8359 26966
rect 9724 26936 9844 26966
rect 7925 26890 7991 26893
rect 7925 26888 8908 26890
rect 7925 26832 7930 26888
rect 7986 26832 8908 26888
rect 7925 26830 8908 26832
rect 7925 26827 7991 26830
rect 8848 26754 8908 26830
rect 9724 26754 9844 26784
rect 8848 26694 9844 26754
rect 1946 26688 2262 26689
rect 1946 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2262 26688
rect 1946 26623 2262 26624
rect 7946 26688 8262 26689
rect 7946 26624 7952 26688
rect 8016 26624 8032 26688
rect 8096 26624 8112 26688
rect 8176 26624 8192 26688
rect 8256 26624 8262 26688
rect 9724 26664 9844 26694
rect 7946 26623 8262 26624
rect 8293 26482 8359 26485
rect 9724 26482 9844 26512
rect 8293 26480 9844 26482
rect 8293 26424 8298 26480
rect 8354 26424 9844 26480
rect 8293 26422 9844 26424
rect 8293 26419 8359 26422
rect 9724 26392 9844 26422
rect 7598 26284 7604 26348
rect 7668 26346 7674 26348
rect 8017 26346 8083 26349
rect 7668 26344 8083 26346
rect 7668 26288 8022 26344
rect 8078 26288 8083 26344
rect 7668 26286 8083 26288
rect 7668 26284 7674 26286
rect 8017 26283 8083 26286
rect 8753 26210 8819 26213
rect 9724 26210 9844 26240
rect 8753 26208 9844 26210
rect 8753 26152 8758 26208
rect 8814 26152 9844 26208
rect 8753 26150 9844 26152
rect 8753 26147 8819 26150
rect 3006 26144 3322 26145
rect 3006 26080 3012 26144
rect 3076 26080 3092 26144
rect 3156 26080 3172 26144
rect 3236 26080 3252 26144
rect 3316 26080 3322 26144
rect 9724 26120 9844 26150
rect 3006 26079 3322 26080
rect 0 25938 120 25968
rect 1209 25938 1275 25941
rect 0 25936 1275 25938
rect 0 25880 1214 25936
rect 1270 25880 1275 25936
rect 0 25878 1275 25880
rect 0 25848 120 25878
rect 1209 25875 1275 25878
rect 8293 25938 8359 25941
rect 9724 25938 9844 25968
rect 8293 25936 9844 25938
rect 8293 25880 8298 25936
rect 8354 25880 9844 25936
rect 8293 25878 9844 25880
rect 8293 25875 8359 25878
rect 9724 25848 9844 25878
rect 7925 25802 7991 25805
rect 7925 25800 9138 25802
rect 7925 25744 7930 25800
rect 7986 25744 9138 25800
rect 7925 25742 9138 25744
rect 7925 25739 7991 25742
rect 9078 25666 9138 25742
rect 9724 25666 9844 25696
rect 9078 25606 9844 25666
rect 1946 25600 2262 25601
rect 1946 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2262 25600
rect 1946 25535 2262 25536
rect 7946 25600 8262 25601
rect 7946 25536 7952 25600
rect 8016 25536 8032 25600
rect 8096 25536 8112 25600
rect 8176 25536 8192 25600
rect 8256 25536 8262 25600
rect 9724 25576 9844 25606
rect 7946 25535 8262 25536
rect 8293 25394 8359 25397
rect 9724 25394 9844 25424
rect 8293 25392 9844 25394
rect 8293 25336 8298 25392
rect 8354 25336 9844 25392
rect 8293 25334 9844 25336
rect 8293 25331 8359 25334
rect 9724 25304 9844 25334
rect 3049 25258 3115 25261
rect 3550 25258 3556 25260
rect 3049 25256 3556 25258
rect 3049 25200 3054 25256
rect 3110 25200 3556 25256
rect 3049 25198 3556 25200
rect 3049 25195 3115 25198
rect 3550 25196 3556 25198
rect 3620 25196 3626 25260
rect 7925 25122 7991 25125
rect 9724 25122 9844 25152
rect 7925 25120 9844 25122
rect 7925 25064 7930 25120
rect 7986 25064 9844 25120
rect 7925 25062 9844 25064
rect 7925 25059 7991 25062
rect 3006 25056 3322 25057
rect 3006 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3172 25056
rect 3236 24992 3252 25056
rect 3316 24992 3322 25056
rect 9724 25032 9844 25062
rect 3006 24991 3322 24992
rect 7005 24986 7071 24989
rect 7005 24984 7114 24986
rect 7005 24928 7010 24984
rect 7066 24928 7114 24984
rect 7005 24923 7114 24928
rect 0 24578 120 24608
rect 7054 24581 7114 24923
rect 7230 24788 7236 24852
rect 7300 24850 7306 24852
rect 7649 24850 7715 24853
rect 7300 24848 7715 24850
rect 7300 24792 7654 24848
rect 7710 24792 7715 24848
rect 7300 24790 7715 24792
rect 7300 24788 7306 24790
rect 7649 24787 7715 24790
rect 8293 24850 8359 24853
rect 9724 24850 9844 24880
rect 8293 24848 9844 24850
rect 8293 24792 8298 24848
rect 8354 24792 9844 24848
rect 8293 24790 9844 24792
rect 8293 24787 8359 24790
rect 9724 24760 9844 24790
rect 7281 24714 7347 24717
rect 7833 24714 7899 24717
rect 7281 24712 7899 24714
rect 7281 24656 7286 24712
rect 7342 24656 7838 24712
rect 7894 24656 7899 24712
rect 7281 24654 7899 24656
rect 7281 24651 7347 24654
rect 7833 24651 7899 24654
rect 841 24578 907 24581
rect 0 24576 907 24578
rect 0 24520 846 24576
rect 902 24520 907 24576
rect 0 24518 907 24520
rect 7054 24576 7163 24581
rect 7054 24520 7102 24576
rect 7158 24520 7163 24576
rect 7054 24518 7163 24520
rect 0 24488 120 24518
rect 841 24515 907 24518
rect 7097 24515 7163 24518
rect 9029 24578 9095 24581
rect 9724 24578 9844 24608
rect 9029 24576 9844 24578
rect 9029 24520 9034 24576
rect 9090 24520 9844 24576
rect 9029 24518 9844 24520
rect 9029 24515 9095 24518
rect 1946 24512 2262 24513
rect 1946 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2262 24512
rect 1946 24447 2262 24448
rect 7946 24512 8262 24513
rect 7946 24448 7952 24512
rect 8016 24448 8032 24512
rect 8096 24448 8112 24512
rect 8176 24448 8192 24512
rect 8256 24448 8262 24512
rect 9724 24488 9844 24518
rect 7946 24447 8262 24448
rect 7833 24306 7899 24309
rect 9724 24306 9844 24336
rect 7833 24304 9844 24306
rect 7833 24248 7838 24304
rect 7894 24248 9844 24304
rect 7833 24246 9844 24248
rect 7833 24243 7899 24246
rect 9724 24216 9844 24246
rect 5390 23972 5396 24036
rect 5460 24034 5466 24036
rect 7005 24034 7071 24037
rect 5460 24032 7071 24034
rect 5460 23976 7010 24032
rect 7066 23976 7071 24032
rect 5460 23974 7071 23976
rect 5460 23972 5466 23974
rect 7005 23971 7071 23974
rect 8293 24034 8359 24037
rect 9724 24034 9844 24064
rect 8293 24032 9844 24034
rect 8293 23976 8298 24032
rect 8354 23976 9844 24032
rect 8293 23974 9844 23976
rect 8293 23971 8359 23974
rect 3006 23968 3322 23969
rect 3006 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3172 23968
rect 3236 23904 3252 23968
rect 3316 23904 3322 23968
rect 9724 23944 9844 23974
rect 3006 23903 3322 23904
rect 7925 23762 7991 23765
rect 9724 23762 9844 23792
rect 7925 23760 9844 23762
rect 7925 23704 7930 23760
rect 7986 23704 9844 23760
rect 7925 23702 9844 23704
rect 7925 23699 7991 23702
rect 9724 23672 9844 23702
rect 3693 23492 3759 23493
rect 3693 23488 3740 23492
rect 3804 23490 3810 23492
rect 4981 23490 5047 23493
rect 5206 23490 5212 23492
rect 3693 23432 3698 23488
rect 3693 23428 3740 23432
rect 3804 23430 3850 23490
rect 4981 23488 5212 23490
rect 4981 23432 4986 23488
rect 5042 23432 5212 23488
rect 4981 23430 5212 23432
rect 3804 23428 3810 23430
rect 3693 23427 3759 23428
rect 4981 23427 5047 23430
rect 5206 23428 5212 23430
rect 5276 23428 5282 23492
rect 6494 23428 6500 23492
rect 6564 23490 6570 23492
rect 6729 23490 6795 23493
rect 6564 23488 6795 23490
rect 6564 23432 6734 23488
rect 6790 23432 6795 23488
rect 6564 23430 6795 23432
rect 6564 23428 6570 23430
rect 6729 23427 6795 23430
rect 9029 23490 9095 23493
rect 9724 23490 9844 23520
rect 9029 23488 9844 23490
rect 9029 23432 9034 23488
rect 9090 23432 9844 23488
rect 9029 23430 9844 23432
rect 9029 23427 9095 23430
rect 1946 23424 2262 23425
rect 1946 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2262 23424
rect 1946 23359 2262 23360
rect 7946 23424 8262 23425
rect 7946 23360 7952 23424
rect 8016 23360 8032 23424
rect 8096 23360 8112 23424
rect 8176 23360 8192 23424
rect 8256 23360 8262 23424
rect 9724 23400 9844 23430
rect 7946 23359 8262 23360
rect 0 23218 120 23248
rect 289 23218 355 23221
rect 0 23216 355 23218
rect 0 23160 294 23216
rect 350 23160 355 23216
rect 0 23158 355 23160
rect 0 23128 120 23158
rect 289 23155 355 23158
rect 8845 23218 8911 23221
rect 9724 23218 9844 23248
rect 8845 23216 9844 23218
rect 8845 23160 8850 23216
rect 8906 23160 9844 23216
rect 8845 23158 9844 23160
rect 8845 23155 8911 23158
rect 9724 23128 9844 23158
rect 8293 22946 8359 22949
rect 9724 22946 9844 22976
rect 8293 22944 9844 22946
rect 8293 22888 8298 22944
rect 8354 22888 9844 22944
rect 8293 22886 9844 22888
rect 8293 22883 8359 22886
rect 3006 22880 3322 22881
rect 3006 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3172 22880
rect 3236 22816 3252 22880
rect 3316 22816 3322 22880
rect 9724 22856 9844 22886
rect 3006 22815 3322 22816
rect 7649 22810 7715 22813
rect 9438 22810 9444 22812
rect 7649 22808 9444 22810
rect 7649 22752 7654 22808
rect 7710 22752 9444 22808
rect 7649 22750 9444 22752
rect 7649 22747 7715 22750
rect 9438 22748 9444 22750
rect 9508 22748 9514 22812
rect 7925 22674 7991 22677
rect 9724 22674 9844 22704
rect 7925 22672 9844 22674
rect 7925 22616 7930 22672
rect 7986 22616 9844 22672
rect 7925 22614 9844 22616
rect 7925 22611 7991 22614
rect 9724 22584 9844 22614
rect 7414 22476 7420 22540
rect 7484 22538 7490 22540
rect 8109 22538 8175 22541
rect 7484 22536 8175 22538
rect 7484 22480 8114 22536
rect 8170 22480 8175 22536
rect 7484 22478 8175 22480
rect 7484 22476 7490 22478
rect 8109 22475 8175 22478
rect 9305 22538 9371 22541
rect 9438 22538 9444 22540
rect 9305 22536 9444 22538
rect 9305 22480 9310 22536
rect 9366 22480 9444 22536
rect 9305 22478 9444 22480
rect 9305 22475 9371 22478
rect 9438 22476 9444 22478
rect 9508 22476 9514 22540
rect 9029 22402 9095 22405
rect 9724 22402 9844 22432
rect 9029 22400 9844 22402
rect 9029 22344 9034 22400
rect 9090 22344 9844 22400
rect 9029 22342 9844 22344
rect 9029 22339 9095 22342
rect 1946 22336 2262 22337
rect 1946 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2262 22336
rect 1946 22271 2262 22272
rect 7946 22336 8262 22337
rect 7946 22272 7952 22336
rect 8016 22272 8032 22336
rect 8096 22272 8112 22336
rect 8176 22272 8192 22336
rect 8256 22272 8262 22336
rect 9724 22312 9844 22342
rect 7946 22271 8262 22272
rect 7281 22132 7347 22133
rect 7230 22068 7236 22132
rect 7300 22130 7347 22132
rect 7833 22130 7899 22133
rect 9724 22130 9844 22160
rect 7300 22128 7392 22130
rect 7342 22072 7392 22128
rect 7300 22070 7392 22072
rect 7833 22128 9844 22130
rect 7833 22072 7838 22128
rect 7894 22072 9844 22128
rect 7833 22070 9844 22072
rect 7300 22068 7347 22070
rect 7281 22067 7347 22068
rect 7833 22067 7899 22070
rect 9724 22040 9844 22070
rect 0 21858 120 21888
rect 1485 21858 1551 21861
rect 0 21856 1551 21858
rect 0 21800 1490 21856
rect 1546 21800 1551 21856
rect 0 21798 1551 21800
rect 0 21768 120 21798
rect 1485 21795 1551 21798
rect 8293 21858 8359 21861
rect 9724 21858 9844 21888
rect 8293 21856 9844 21858
rect 8293 21800 8298 21856
rect 8354 21800 9844 21856
rect 8293 21798 9844 21800
rect 8293 21795 8359 21798
rect 3006 21792 3322 21793
rect 3006 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3172 21792
rect 3236 21728 3252 21792
rect 3316 21728 3322 21792
rect 9724 21768 9844 21798
rect 3006 21727 3322 21728
rect 7925 21586 7991 21589
rect 9724 21586 9844 21616
rect 7925 21584 9844 21586
rect 7925 21528 7930 21584
rect 7986 21528 9844 21584
rect 7925 21526 9844 21528
rect 7925 21523 7991 21526
rect 9724 21496 9844 21526
rect 8017 21450 8083 21453
rect 8334 21450 8340 21452
rect 8017 21448 8340 21450
rect 8017 21392 8022 21448
rect 8078 21392 8340 21448
rect 8017 21390 8340 21392
rect 8017 21387 8083 21390
rect 8334 21388 8340 21390
rect 8404 21388 8410 21452
rect 9029 21314 9095 21317
rect 9724 21314 9844 21344
rect 9029 21312 9844 21314
rect 9029 21256 9034 21312
rect 9090 21256 9844 21312
rect 9029 21254 9844 21256
rect 9029 21251 9095 21254
rect 1946 21248 2262 21249
rect 1946 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2262 21248
rect 1946 21183 2262 21184
rect 7946 21248 8262 21249
rect 7946 21184 7952 21248
rect 8016 21184 8032 21248
rect 8096 21184 8112 21248
rect 8176 21184 8192 21248
rect 8256 21184 8262 21248
rect 9724 21224 9844 21254
rect 7946 21183 8262 21184
rect 6729 21044 6795 21045
rect 6678 21042 6684 21044
rect 6638 20982 6684 21042
rect 6748 21040 6795 21044
rect 6790 20984 6795 21040
rect 6678 20980 6684 20982
rect 6748 20980 6795 20984
rect 6729 20979 6795 20980
rect 7833 21042 7899 21045
rect 9724 21042 9844 21072
rect 7833 21040 9844 21042
rect 7833 20984 7838 21040
rect 7894 20984 9844 21040
rect 7833 20982 9844 20984
rect 7833 20979 7899 20982
rect 9724 20952 9844 20982
rect 6126 20844 6132 20908
rect 6196 20906 6202 20908
rect 8109 20906 8175 20909
rect 6196 20904 8175 20906
rect 6196 20848 8114 20904
rect 8170 20848 8175 20904
rect 6196 20846 8175 20848
rect 6196 20844 6202 20846
rect 8109 20843 8175 20846
rect 6310 20708 6316 20772
rect 6380 20770 6386 20772
rect 7741 20770 7807 20773
rect 6380 20768 7807 20770
rect 6380 20712 7746 20768
rect 7802 20712 7807 20768
rect 6380 20710 7807 20712
rect 6380 20708 6386 20710
rect 7741 20707 7807 20710
rect 8293 20770 8359 20773
rect 9724 20770 9844 20800
rect 8293 20768 9844 20770
rect 8293 20712 8298 20768
rect 8354 20712 9844 20768
rect 8293 20710 9844 20712
rect 8293 20707 8359 20710
rect 3006 20704 3322 20705
rect 3006 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3172 20704
rect 3236 20640 3252 20704
rect 3316 20640 3322 20704
rect 9724 20680 9844 20710
rect 3006 20639 3322 20640
rect 8569 20634 8635 20637
rect 9254 20634 9260 20636
rect 8569 20632 9260 20634
rect 8569 20576 8574 20632
rect 8630 20576 9260 20632
rect 8569 20574 9260 20576
rect 8569 20571 8635 20574
rect 9254 20572 9260 20574
rect 9324 20572 9330 20636
rect 0 20498 120 20528
rect 933 20498 999 20501
rect 0 20496 999 20498
rect 0 20440 938 20496
rect 994 20440 999 20496
rect 0 20438 999 20440
rect 0 20408 120 20438
rect 933 20435 999 20438
rect 8201 20498 8267 20501
rect 8702 20498 8708 20500
rect 8201 20496 8708 20498
rect 8201 20440 8206 20496
rect 8262 20440 8708 20496
rect 8201 20438 8708 20440
rect 8201 20435 8267 20438
rect 8702 20436 8708 20438
rect 8772 20436 8778 20500
rect 8845 20498 8911 20501
rect 9724 20498 9844 20528
rect 8845 20496 9844 20498
rect 8845 20440 8850 20496
rect 8906 20440 9844 20496
rect 8845 20438 9844 20440
rect 8845 20435 8911 20438
rect 9724 20408 9844 20438
rect 7230 20300 7236 20364
rect 7300 20362 7306 20364
rect 8109 20362 8175 20365
rect 7300 20360 8175 20362
rect 7300 20304 8114 20360
rect 8170 20304 8175 20360
rect 7300 20302 8175 20304
rect 7300 20300 7306 20302
rect 8109 20299 8175 20302
rect 9029 20226 9095 20229
rect 9724 20226 9844 20256
rect 9029 20224 9844 20226
rect 9029 20168 9034 20224
rect 9090 20168 9844 20224
rect 9029 20166 9844 20168
rect 9029 20163 9095 20166
rect 1946 20160 2262 20161
rect 1946 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2262 20160
rect 1946 20095 2262 20096
rect 7946 20160 8262 20161
rect 7946 20096 7952 20160
rect 8016 20096 8032 20160
rect 8096 20096 8112 20160
rect 8176 20096 8192 20160
rect 8256 20096 8262 20160
rect 9724 20136 9844 20166
rect 7946 20095 8262 20096
rect 7833 19954 7899 19957
rect 9724 19954 9844 19984
rect 7833 19952 9844 19954
rect 7833 19896 7838 19952
rect 7894 19896 9844 19952
rect 7833 19894 9844 19896
rect 7833 19891 7899 19894
rect 9724 19864 9844 19894
rect 8293 19682 8359 19685
rect 9724 19682 9844 19712
rect 8293 19680 9844 19682
rect 8293 19624 8298 19680
rect 8354 19624 9844 19680
rect 8293 19622 9844 19624
rect 8293 19619 8359 19622
rect 3006 19616 3322 19617
rect 3006 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3322 19616
rect 9724 19592 9844 19622
rect 3006 19551 3322 19552
rect 3509 19546 3575 19549
rect 3918 19546 3924 19548
rect 3509 19544 3924 19546
rect 3509 19488 3514 19544
rect 3570 19488 3924 19544
rect 3509 19486 3924 19488
rect 3509 19483 3575 19486
rect 3918 19484 3924 19486
rect 3988 19484 3994 19548
rect 7925 19410 7991 19413
rect 9724 19410 9844 19440
rect 7925 19408 9844 19410
rect 7925 19352 7930 19408
rect 7986 19352 9844 19408
rect 7925 19350 9844 19352
rect 7925 19347 7991 19350
rect 9724 19320 9844 19350
rect 0 19138 120 19168
rect 749 19138 815 19141
rect 0 19136 815 19138
rect 0 19080 754 19136
rect 810 19080 815 19136
rect 0 19078 815 19080
rect 0 19048 120 19078
rect 749 19075 815 19078
rect 9029 19138 9095 19141
rect 9724 19138 9844 19168
rect 9029 19136 9844 19138
rect 9029 19080 9034 19136
rect 9090 19080 9844 19136
rect 9029 19078 9844 19080
rect 9029 19075 9095 19078
rect 1946 19072 2262 19073
rect 1946 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2262 19072
rect 1946 19007 2262 19008
rect 7946 19072 8262 19073
rect 7946 19008 7952 19072
rect 8016 19008 8032 19072
rect 8096 19008 8112 19072
rect 8176 19008 8192 19072
rect 8256 19008 8262 19072
rect 9724 19048 9844 19078
rect 7946 19007 8262 19008
rect 8753 18866 8819 18869
rect 9724 18866 9844 18896
rect 8753 18864 9844 18866
rect 8753 18808 8758 18864
rect 8814 18808 9844 18864
rect 8753 18806 9844 18808
rect 8753 18803 8819 18806
rect 9724 18776 9844 18806
rect 8293 18594 8359 18597
rect 9724 18594 9844 18624
rect 8293 18592 9844 18594
rect 8293 18536 8298 18592
rect 8354 18536 9844 18592
rect 8293 18534 9844 18536
rect 8293 18531 8359 18534
rect 3006 18528 3322 18529
rect 3006 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3322 18528
rect 9724 18504 9844 18534
rect 3006 18463 3322 18464
rect 7925 18322 7991 18325
rect 9724 18322 9844 18352
rect 7925 18320 9844 18322
rect 7925 18264 7930 18320
rect 7986 18264 9844 18320
rect 7925 18262 9844 18264
rect 7925 18259 7991 18262
rect 9724 18232 9844 18262
rect 8937 18050 9003 18053
rect 9724 18050 9844 18080
rect 8937 18048 9844 18050
rect 8937 17992 8942 18048
rect 8998 17992 9844 18048
rect 8937 17990 9844 17992
rect 8937 17987 9003 17990
rect 1946 17984 2262 17985
rect 1946 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2262 17984
rect 1946 17919 2262 17920
rect 7946 17984 8262 17985
rect 7946 17920 7952 17984
rect 8016 17920 8032 17984
rect 8096 17920 8112 17984
rect 8176 17920 8192 17984
rect 8256 17920 8262 17984
rect 9724 17960 9844 17990
rect 7946 17919 8262 17920
rect 7097 17914 7163 17917
rect 7414 17914 7420 17916
rect 7097 17912 7420 17914
rect 7097 17856 7102 17912
rect 7158 17856 7420 17912
rect 7097 17854 7420 17856
rect 7097 17851 7163 17854
rect 7414 17852 7420 17854
rect 7484 17852 7490 17916
rect 0 17778 120 17808
rect 1117 17778 1183 17781
rect 0 17776 1183 17778
rect 0 17720 1122 17776
rect 1178 17720 1183 17776
rect 0 17718 1183 17720
rect 0 17688 120 17718
rect 1117 17715 1183 17718
rect 8385 17778 8451 17781
rect 9724 17778 9844 17808
rect 8385 17776 9844 17778
rect 8385 17720 8390 17776
rect 8446 17720 9844 17776
rect 8385 17718 9844 17720
rect 8385 17715 8451 17718
rect 9724 17688 9844 17718
rect 8385 17644 8451 17645
rect 8334 17580 8340 17644
rect 8404 17642 8451 17644
rect 8404 17640 8496 17642
rect 8446 17584 8496 17640
rect 8404 17582 8496 17584
rect 8404 17580 8451 17582
rect 8385 17579 8451 17580
rect 8661 17506 8727 17509
rect 9724 17506 9844 17536
rect 8661 17504 9844 17506
rect 8661 17448 8666 17504
rect 8722 17448 9844 17504
rect 8661 17446 9844 17448
rect 8661 17443 8727 17446
rect 3006 17440 3322 17441
rect 3006 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3322 17440
rect 9724 17416 9844 17446
rect 3006 17375 3322 17376
rect 9489 17234 9555 17237
rect 9724 17234 9844 17264
rect 9489 17232 9844 17234
rect 9489 17176 9494 17232
rect 9550 17176 9844 17232
rect 9489 17174 9844 17176
rect 9489 17171 9555 17174
rect 9724 17144 9844 17174
rect 9305 16962 9371 16965
rect 9724 16962 9844 16992
rect 9305 16960 9844 16962
rect 9305 16904 9310 16960
rect 9366 16904 9844 16960
rect 9305 16902 9844 16904
rect 9305 16899 9371 16902
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 7946 16896 8262 16897
rect 7946 16832 7952 16896
rect 8016 16832 8032 16896
rect 8096 16832 8112 16896
rect 8176 16832 8192 16896
rect 8256 16832 8262 16896
rect 9724 16872 9844 16902
rect 7946 16831 8262 16832
rect 9121 16690 9187 16693
rect 9724 16690 9844 16720
rect 9121 16688 9844 16690
rect 9121 16632 9126 16688
rect 9182 16632 9844 16688
rect 9121 16630 9844 16632
rect 9121 16627 9187 16630
rect 9724 16600 9844 16630
rect 0 16418 120 16448
rect 841 16418 907 16421
rect 0 16416 907 16418
rect 0 16360 846 16416
rect 902 16360 907 16416
rect 0 16358 907 16360
rect 0 16328 120 16358
rect 841 16355 907 16358
rect 4981 16418 5047 16421
rect 9724 16418 9844 16448
rect 4981 16416 9844 16418
rect 4981 16360 4986 16416
rect 5042 16360 9844 16416
rect 4981 16358 9844 16360
rect 4981 16355 5047 16358
rect 3006 16352 3322 16353
rect 3006 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3322 16352
rect 9724 16328 9844 16358
rect 3006 16287 3322 16288
rect 1526 16220 1532 16284
rect 1596 16282 1602 16284
rect 1853 16282 1919 16285
rect 1596 16280 1919 16282
rect 1596 16224 1858 16280
rect 1914 16224 1919 16280
rect 1596 16222 1919 16224
rect 1596 16220 1602 16222
rect 1853 16219 1919 16222
rect 4889 16282 4955 16285
rect 5022 16282 5028 16284
rect 4889 16280 5028 16282
rect 4889 16224 4894 16280
rect 4950 16224 5028 16280
rect 4889 16222 5028 16224
rect 4889 16219 4955 16222
rect 5022 16220 5028 16222
rect 5092 16220 5098 16284
rect 5214 16222 8402 16282
rect 4061 16146 4127 16149
rect 5214 16146 5274 16222
rect 4061 16144 5274 16146
rect 4061 16088 4066 16144
rect 4122 16088 5274 16144
rect 4061 16086 5274 16088
rect 6729 16146 6795 16149
rect 8342 16146 8402 16222
rect 9724 16146 9844 16176
rect 6729 16144 6930 16146
rect 6729 16088 6734 16144
rect 6790 16088 6930 16144
rect 6729 16086 6930 16088
rect 8342 16086 9844 16146
rect 4061 16083 4127 16086
rect 6729 16083 6795 16086
rect 6870 16010 6930 16086
rect 9724 16056 9844 16086
rect 6870 15950 8402 16010
rect 8342 15874 8402 15950
rect 9724 15874 9844 15904
rect 8342 15814 9844 15874
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 7946 15808 8262 15809
rect 7946 15744 7952 15808
rect 8016 15744 8032 15808
rect 8096 15744 8112 15808
rect 8176 15744 8192 15808
rect 8256 15744 8262 15808
rect 9724 15784 9844 15814
rect 7946 15743 8262 15744
rect 5073 15602 5139 15605
rect 9724 15602 9844 15632
rect 5073 15600 9844 15602
rect 5073 15544 5078 15600
rect 5134 15544 9844 15600
rect 5073 15542 9844 15544
rect 5073 15539 5139 15542
rect 9724 15512 9844 15542
rect 6453 15466 6519 15469
rect 6453 15464 6930 15466
rect 6453 15408 6458 15464
rect 6514 15408 6930 15464
rect 6453 15406 6930 15408
rect 6453 15403 6519 15406
rect 6870 15330 6930 15406
rect 7230 15404 7236 15468
rect 7300 15466 7306 15468
rect 7373 15466 7439 15469
rect 7300 15464 7439 15466
rect 7300 15408 7378 15464
rect 7434 15408 7439 15464
rect 7300 15406 7439 15408
rect 7300 15404 7306 15406
rect 7373 15403 7439 15406
rect 7598 15404 7604 15468
rect 7668 15466 7674 15468
rect 7833 15466 7899 15469
rect 7668 15464 7899 15466
rect 7668 15408 7838 15464
rect 7894 15408 7899 15464
rect 7668 15406 7899 15408
rect 7668 15404 7674 15406
rect 7833 15403 7899 15406
rect 9724 15330 9844 15360
rect 6870 15270 9844 15330
rect 3006 15264 3322 15265
rect 3006 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3322 15264
rect 9724 15240 9844 15270
rect 3006 15199 3322 15200
rect 0 15058 120 15088
rect 749 15058 815 15061
rect 0 15056 815 15058
rect 0 15000 754 15056
rect 810 15000 815 15056
rect 0 14998 815 15000
rect 0 14968 120 14998
rect 749 14995 815 14998
rect 9029 15058 9095 15061
rect 9724 15058 9844 15088
rect 9029 15056 9844 15058
rect 9029 15000 9034 15056
rect 9090 15000 9844 15056
rect 9029 14998 9844 15000
rect 9029 14995 9095 14998
rect 9724 14968 9844 14998
rect 6913 14922 6979 14925
rect 7557 14922 7623 14925
rect 6913 14920 7623 14922
rect 6913 14864 6918 14920
rect 6974 14864 7562 14920
rect 7618 14864 7623 14920
rect 6913 14862 7623 14864
rect 6913 14859 6979 14862
rect 7557 14859 7623 14862
rect 8845 14786 8911 14789
rect 9724 14786 9844 14816
rect 8845 14784 9844 14786
rect 8845 14728 8850 14784
rect 8906 14728 9844 14784
rect 8845 14726 9844 14728
rect 8845 14723 8911 14726
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 7946 14720 8262 14721
rect 7946 14656 7952 14720
rect 8016 14656 8032 14720
rect 8096 14656 8112 14720
rect 8176 14656 8192 14720
rect 8256 14656 8262 14720
rect 9724 14696 9844 14726
rect 7946 14655 8262 14656
rect 7649 14514 7715 14517
rect 9724 14514 9844 14544
rect 7649 14512 9844 14514
rect 7649 14456 7654 14512
rect 7710 14456 9844 14512
rect 7649 14454 9844 14456
rect 7649 14451 7715 14454
rect 9724 14424 9844 14454
rect 7557 14242 7623 14245
rect 9724 14242 9844 14272
rect 7557 14240 9844 14242
rect 7557 14184 7562 14240
rect 7618 14184 9844 14240
rect 7557 14182 9844 14184
rect 7557 14179 7623 14182
rect 3006 14176 3322 14177
rect 3006 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3322 14176
rect 9724 14152 9844 14182
rect 3006 14111 3322 14112
rect 9397 13970 9463 13973
rect 9724 13970 9844 14000
rect 9397 13968 9844 13970
rect 9397 13912 9402 13968
rect 9458 13912 9844 13968
rect 9397 13910 9844 13912
rect 9397 13907 9463 13910
rect 9724 13880 9844 13910
rect 1853 13834 1919 13837
rect 6177 13836 6243 13837
rect 4654 13834 4660 13836
rect 1853 13832 4660 13834
rect 1853 13776 1858 13832
rect 1914 13776 4660 13832
rect 1853 13774 4660 13776
rect 1853 13771 1919 13774
rect 4654 13772 4660 13774
rect 4724 13772 4730 13836
rect 6126 13834 6132 13836
rect 6086 13774 6132 13834
rect 6196 13832 6243 13836
rect 6238 13776 6243 13832
rect 6126 13772 6132 13774
rect 6196 13772 6243 13776
rect 6177 13771 6243 13772
rect 0 13698 120 13728
rect 1025 13698 1091 13701
rect 0 13696 1091 13698
rect 0 13640 1030 13696
rect 1086 13640 1091 13696
rect 0 13638 1091 13640
rect 0 13608 120 13638
rect 1025 13635 1091 13638
rect 8569 13698 8635 13701
rect 9724 13698 9844 13728
rect 8569 13696 9844 13698
rect 8569 13640 8574 13696
rect 8630 13640 9844 13696
rect 8569 13638 9844 13640
rect 8569 13635 8635 13638
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 7946 13632 8262 13633
rect 7946 13568 7952 13632
rect 8016 13568 8032 13632
rect 8096 13568 8112 13632
rect 8176 13568 8192 13632
rect 8256 13568 8262 13632
rect 9724 13608 9844 13638
rect 7946 13567 8262 13568
rect 8753 13426 8819 13429
rect 9724 13426 9844 13456
rect 8753 13424 9844 13426
rect 8753 13368 8758 13424
rect 8814 13368 9844 13424
rect 8753 13366 9844 13368
rect 8753 13363 8819 13366
rect 9724 13336 9844 13366
rect 8477 13154 8543 13157
rect 9724 13154 9844 13184
rect 8477 13152 9844 13154
rect 8477 13096 8482 13152
rect 8538 13096 9844 13152
rect 8477 13094 9844 13096
rect 8477 13091 8543 13094
rect 3006 13088 3322 13089
rect 3006 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3322 13088
rect 9724 13064 9844 13094
rect 3006 13023 3322 13024
rect 8293 12882 8359 12885
rect 9724 12882 9844 12912
rect 8293 12880 9844 12882
rect 8293 12824 8298 12880
rect 8354 12824 9844 12880
rect 8293 12822 9844 12824
rect 8293 12819 8359 12822
rect 9724 12792 9844 12822
rect 9489 12610 9555 12613
rect 9724 12610 9844 12640
rect 9489 12608 9844 12610
rect 9489 12552 9494 12608
rect 9550 12552 9844 12608
rect 9489 12550 9844 12552
rect 9489 12547 9555 12550
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 7946 12544 8262 12545
rect 7946 12480 7952 12544
rect 8016 12480 8032 12544
rect 8096 12480 8112 12544
rect 8176 12480 8192 12544
rect 8256 12480 8262 12544
rect 9724 12520 9844 12550
rect 7946 12479 8262 12480
rect 0 12338 120 12368
rect 749 12338 815 12341
rect 0 12336 815 12338
rect 0 12280 754 12336
rect 810 12280 815 12336
rect 0 12278 815 12280
rect 0 12248 120 12278
rect 749 12275 815 12278
rect 8753 12338 8819 12341
rect 9724 12338 9844 12368
rect 8753 12336 9844 12338
rect 8753 12280 8758 12336
rect 8814 12280 9844 12336
rect 8753 12278 9844 12280
rect 8753 12275 8819 12278
rect 9724 12248 9844 12278
rect 9581 12066 9647 12069
rect 9724 12066 9844 12096
rect 9581 12064 9844 12066
rect 9581 12008 9586 12064
rect 9642 12008 9844 12064
rect 9581 12006 9844 12008
rect 9581 12003 9647 12006
rect 3006 12000 3322 12001
rect 3006 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3322 12000
rect 9724 11976 9844 12006
rect 3006 11935 3322 11936
rect 9438 11732 9444 11796
rect 9508 11794 9514 11796
rect 9724 11794 9844 11824
rect 9508 11734 9844 11794
rect 9508 11732 9514 11734
rect 9724 11704 9844 11734
rect 1710 11596 1716 11660
rect 1780 11658 1786 11660
rect 1853 11658 1919 11661
rect 1780 11656 1919 11658
rect 1780 11600 1858 11656
rect 1914 11600 1919 11656
rect 1780 11598 1919 11600
rect 1780 11596 1786 11598
rect 1853 11595 1919 11598
rect 5993 11658 6059 11661
rect 6310 11658 6316 11660
rect 5993 11656 6316 11658
rect 5993 11600 5998 11656
rect 6054 11600 6316 11656
rect 5993 11598 6316 11600
rect 5993 11595 6059 11598
rect 6310 11596 6316 11598
rect 6380 11596 6386 11660
rect 8661 11522 8727 11525
rect 9724 11522 9844 11552
rect 8661 11520 9844 11522
rect 8661 11464 8666 11520
rect 8722 11464 9844 11520
rect 8661 11462 9844 11464
rect 8661 11459 8727 11462
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 7946 11456 8262 11457
rect 7946 11392 7952 11456
rect 8016 11392 8032 11456
rect 8096 11392 8112 11456
rect 8176 11392 8192 11456
rect 8256 11392 8262 11456
rect 9724 11432 9844 11462
rect 7946 11391 8262 11392
rect 9254 11188 9260 11252
rect 9324 11250 9330 11252
rect 9724 11250 9844 11280
rect 9324 11190 9844 11250
rect 9324 11188 9330 11190
rect 9724 11160 9844 11190
rect 2865 11114 2931 11117
rect 2865 11112 3618 11114
rect 2865 11056 2870 11112
rect 2926 11056 3618 11112
rect 2865 11054 3618 11056
rect 2865 11051 2931 11054
rect 0 10978 120 11008
rect 933 10978 999 10981
rect 0 10976 999 10978
rect 0 10920 938 10976
rect 994 10920 999 10976
rect 0 10918 999 10920
rect 3558 10978 3618 11054
rect 9724 10978 9844 11008
rect 3558 10918 9844 10978
rect 0 10888 120 10918
rect 933 10915 999 10918
rect 3006 10912 3322 10913
rect 3006 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3322 10912
rect 9724 10888 9844 10918
rect 3006 10847 3322 10848
rect 6494 10644 6500 10708
rect 6564 10706 6570 10708
rect 9724 10706 9844 10736
rect 6564 10646 9844 10706
rect 6564 10644 6570 10646
rect 9724 10616 9844 10646
rect 8937 10434 9003 10437
rect 9724 10434 9844 10464
rect 8937 10432 9844 10434
rect 8937 10376 8942 10432
rect 8998 10376 9844 10432
rect 8937 10374 9844 10376
rect 8937 10371 9003 10374
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 7946 10368 8262 10369
rect 7946 10304 7952 10368
rect 8016 10304 8032 10368
rect 8096 10304 8112 10368
rect 8176 10304 8192 10368
rect 8256 10304 8262 10368
rect 9724 10344 9844 10374
rect 7946 10303 8262 10304
rect 8753 10162 8819 10165
rect 9724 10162 9844 10192
rect 8753 10160 9844 10162
rect 8753 10104 8758 10160
rect 8814 10104 9844 10160
rect 8753 10102 9844 10104
rect 8753 10099 8819 10102
rect 9724 10072 9844 10102
rect 8477 9890 8543 9893
rect 9724 9890 9844 9920
rect 8477 9888 9844 9890
rect 8477 9832 8482 9888
rect 8538 9832 9844 9888
rect 8477 9830 9844 9832
rect 8477 9827 8543 9830
rect 3006 9824 3322 9825
rect 3006 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3322 9824
rect 9724 9800 9844 9830
rect 3006 9759 3322 9760
rect 0 9618 120 9648
rect 565 9618 631 9621
rect 0 9616 631 9618
rect 0 9560 570 9616
rect 626 9560 631 9616
rect 0 9558 631 9560
rect 0 9528 120 9558
rect 565 9555 631 9558
rect 8293 9618 8359 9621
rect 9724 9618 9844 9648
rect 8293 9616 9844 9618
rect 8293 9560 8298 9616
rect 8354 9560 9844 9616
rect 8293 9558 9844 9560
rect 8293 9555 8359 9558
rect 9724 9528 9844 9558
rect 7649 9482 7715 9485
rect 8702 9482 8708 9484
rect 7649 9480 8708 9482
rect 7649 9424 7654 9480
rect 7710 9424 8708 9480
rect 7649 9422 8708 9424
rect 7649 9419 7715 9422
rect 8702 9420 8708 9422
rect 8772 9420 8778 9484
rect 8385 9346 8451 9349
rect 9724 9346 9844 9376
rect 8385 9344 9844 9346
rect 8385 9288 8390 9344
rect 8446 9288 9844 9344
rect 8385 9286 9844 9288
rect 8385 9283 8451 9286
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 7946 9280 8262 9281
rect 7946 9216 7952 9280
rect 8016 9216 8032 9280
rect 8096 9216 8112 9280
rect 8176 9216 8192 9280
rect 8256 9216 8262 9280
rect 9724 9256 9844 9286
rect 7946 9215 8262 9216
rect 6913 9074 6979 9077
rect 9724 9074 9844 9104
rect 6913 9072 9844 9074
rect 6913 9016 6918 9072
rect 6974 9016 9844 9072
rect 6913 9014 9844 9016
rect 6913 9011 6979 9014
rect 9724 8984 9844 9014
rect 7097 8802 7163 8805
rect 9724 8802 9844 8832
rect 7097 8800 9844 8802
rect 7097 8744 7102 8800
rect 7158 8744 9844 8800
rect 7097 8742 9844 8744
rect 7097 8739 7163 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 9724 8712 9844 8742
rect 3006 8671 3322 8672
rect 9438 8468 9444 8532
rect 9508 8530 9514 8532
rect 9724 8530 9844 8560
rect 9508 8470 9844 8530
rect 9508 8468 9514 8470
rect 9724 8440 9844 8470
rect 0 8258 120 8288
rect 473 8258 539 8261
rect 0 8256 539 8258
rect 0 8200 478 8256
rect 534 8200 539 8256
rect 0 8198 539 8200
rect 0 8168 120 8198
rect 473 8195 539 8198
rect 4613 8258 4679 8261
rect 5717 8258 5783 8261
rect 4613 8256 5783 8258
rect 4613 8200 4618 8256
rect 4674 8200 5722 8256
rect 5778 8200 5783 8256
rect 4613 8198 5783 8200
rect 4613 8195 4679 8198
rect 5717 8195 5783 8198
rect 8385 8258 8451 8261
rect 9724 8258 9844 8288
rect 8385 8256 9844 8258
rect 8385 8200 8390 8256
rect 8446 8200 9844 8256
rect 8385 8198 9844 8200
rect 8385 8195 8451 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 9724 8168 9844 8198
rect 7946 8127 8262 8128
rect 7005 7986 7071 7989
rect 9724 7986 9844 8016
rect 7005 7984 9844 7986
rect 7005 7928 7010 7984
rect 7066 7928 9844 7984
rect 7005 7926 9844 7928
rect 7005 7923 7071 7926
rect 9724 7896 9844 7926
rect 7833 7714 7899 7717
rect 9724 7714 9844 7744
rect 7833 7712 9844 7714
rect 7833 7656 7838 7712
rect 7894 7656 9844 7712
rect 7833 7654 9844 7656
rect 7833 7651 7899 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 9724 7624 9844 7654
rect 3006 7583 3322 7584
rect 7189 7442 7255 7445
rect 9724 7442 9844 7472
rect 7189 7440 9844 7442
rect 7189 7384 7194 7440
rect 7250 7384 9844 7440
rect 7189 7382 9844 7384
rect 7189 7379 7255 7382
rect 9724 7352 9844 7382
rect 5809 7306 5875 7309
rect 5809 7304 9368 7306
rect 5809 7248 5814 7304
rect 5870 7248 9368 7304
rect 5809 7246 9368 7248
rect 5809 7243 5875 7246
rect 9308 7170 9368 7246
rect 9724 7170 9844 7200
rect 9308 7110 9844 7170
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 9724 7080 9844 7110
rect 7946 7039 8262 7040
rect 0 6898 120 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 120 6838
rect 2773 6835 2839 6838
rect 6729 6898 6795 6901
rect 9724 6898 9844 6928
rect 6729 6896 9844 6898
rect 6729 6840 6734 6896
rect 6790 6840 9844 6896
rect 6729 6838 9844 6840
rect 6729 6835 6795 6838
rect 9724 6808 9844 6838
rect 7281 6626 7347 6629
rect 9724 6626 9844 6656
rect 7281 6624 9844 6626
rect 7281 6568 7286 6624
rect 7342 6568 9844 6624
rect 7281 6566 9844 6568
rect 7281 6563 7347 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 9724 6536 9844 6566
rect 3006 6495 3322 6496
rect 9724 6357 9844 6384
rect 9673 6352 9844 6357
rect 9673 6296 9678 6352
rect 9734 6296 9844 6352
rect 9673 6291 9844 6296
rect 9724 6264 9844 6291
rect 5901 6218 5967 6221
rect 5901 6216 8402 6218
rect 5901 6160 5906 6216
rect 5962 6160 8402 6216
rect 5901 6158 8402 6160
rect 5901 6155 5967 6158
rect 8342 6082 8402 6158
rect 9724 6082 9844 6112
rect 8342 6022 9844 6082
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 9724 5992 9844 6022
rect 7946 5951 8262 5952
rect 6361 5810 6427 5813
rect 9724 5810 9844 5840
rect 6361 5808 9844 5810
rect 6361 5752 6366 5808
rect 6422 5752 9844 5808
rect 6361 5750 9844 5752
rect 6361 5747 6427 5750
rect 9724 5720 9844 5750
rect 0 5538 120 5568
rect 197 5538 263 5541
rect 0 5536 263 5538
rect 0 5480 202 5536
rect 258 5480 263 5536
rect 0 5478 263 5480
rect 0 5448 120 5478
rect 197 5475 263 5478
rect 7833 5538 7899 5541
rect 9724 5538 9844 5568
rect 7833 5536 9844 5538
rect 7833 5480 7838 5536
rect 7894 5480 9844 5536
rect 7833 5478 9844 5480
rect 7833 5475 7899 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 9724 5448 9844 5478
rect 3006 5407 3322 5408
rect 7741 5266 7807 5269
rect 9724 5266 9844 5296
rect 7741 5264 9844 5266
rect 7741 5208 7746 5264
rect 7802 5208 9844 5264
rect 7741 5206 9844 5208
rect 7741 5203 7807 5206
rect 9724 5176 9844 5206
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 0 4178 120 4208
rect 381 4178 447 4181
rect 0 4176 447 4178
rect 0 4120 386 4176
rect 442 4120 447 4176
rect 0 4118 447 4120
rect 0 4088 120 4118
rect 381 4115 447 4118
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 0 2821 120 2848
rect 0 2816 171 2821
rect 0 2760 110 2816
rect 166 2760 171 2816
rect 0 2755 171 2760
rect 0 2728 120 2755
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 0 1458 120 1488
rect 657 1458 723 1461
rect 0 1456 723 1458
rect 0 1400 662 1456
rect 718 1400 723 1456
rect 0 1398 723 1400
rect 0 1368 120 1398
rect 657 1395 723 1398
rect 3049 1322 3115 1325
rect 3734 1322 3740 1324
rect 3049 1320 3740 1322
rect 3049 1264 3054 1320
rect 3110 1264 3740 1320
rect 3049 1262 3740 1264
rect 3049 1259 3115 1262
rect 3734 1260 3740 1262
rect 3804 1260 3810 1324
rect 6678 1260 6684 1324
rect 6748 1322 6754 1324
rect 9489 1322 9555 1325
rect 6748 1320 9555 1322
rect 6748 1264 9494 1320
rect 9550 1264 9555 1320
rect 6748 1262 9555 1264
rect 6748 1260 6754 1262
rect 9489 1259 9555 1262
rect 3550 1124 3556 1188
rect 3620 1186 3626 1188
rect 7189 1186 7255 1189
rect 3620 1184 7255 1186
rect 3620 1128 7194 1184
rect 7250 1128 7255 1184
rect 3620 1126 7255 1128
rect 3620 1124 3626 1126
rect 7189 1123 7255 1126
rect 5390 988 5396 1052
rect 5460 1050 5466 1052
rect 9029 1050 9095 1053
rect 5460 1048 9095 1050
rect 5460 992 9034 1048
rect 9090 992 9095 1048
rect 5460 990 9095 992
rect 5460 988 5466 990
rect 9029 987 9095 990
rect 5206 36 5212 100
rect 5276 98 5282 100
rect 7649 98 7715 101
rect 5276 96 7715 98
rect 5276 40 7654 96
rect 7710 40 7715 96
rect 5276 38 7715 40
rect 5276 36 5282 38
rect 7649 35 7715 38
<< via3 >>
rect 3012 42460 3076 42464
rect 3012 42404 3016 42460
rect 3016 42404 3072 42460
rect 3072 42404 3076 42460
rect 3012 42400 3076 42404
rect 3092 42460 3156 42464
rect 3092 42404 3096 42460
rect 3096 42404 3152 42460
rect 3152 42404 3156 42460
rect 3092 42400 3156 42404
rect 3172 42460 3236 42464
rect 3172 42404 3176 42460
rect 3176 42404 3232 42460
rect 3232 42404 3236 42460
rect 3172 42400 3236 42404
rect 3252 42460 3316 42464
rect 3252 42404 3256 42460
rect 3256 42404 3312 42460
rect 3312 42404 3316 42460
rect 3252 42400 3316 42404
rect 1952 41916 2016 41920
rect 1952 41860 1956 41916
rect 1956 41860 2012 41916
rect 2012 41860 2016 41916
rect 1952 41856 2016 41860
rect 2032 41916 2096 41920
rect 2032 41860 2036 41916
rect 2036 41860 2092 41916
rect 2092 41860 2096 41916
rect 2032 41856 2096 41860
rect 2112 41916 2176 41920
rect 2112 41860 2116 41916
rect 2116 41860 2172 41916
rect 2172 41860 2176 41916
rect 2112 41856 2176 41860
rect 2192 41916 2256 41920
rect 2192 41860 2196 41916
rect 2196 41860 2252 41916
rect 2252 41860 2256 41916
rect 2192 41856 2256 41860
rect 7952 41916 8016 41920
rect 7952 41860 7956 41916
rect 7956 41860 8012 41916
rect 8012 41860 8016 41916
rect 7952 41856 8016 41860
rect 8032 41916 8096 41920
rect 8032 41860 8036 41916
rect 8036 41860 8092 41916
rect 8092 41860 8096 41916
rect 8032 41856 8096 41860
rect 8112 41916 8176 41920
rect 8112 41860 8116 41916
rect 8116 41860 8172 41916
rect 8172 41860 8176 41916
rect 8112 41856 8176 41860
rect 8192 41916 8256 41920
rect 8192 41860 8196 41916
rect 8196 41860 8252 41916
rect 8252 41860 8256 41916
rect 8192 41856 8256 41860
rect 1532 41652 1596 41716
rect 1716 41440 1780 41444
rect 1716 41384 1730 41440
rect 1730 41384 1780 41440
rect 1716 41380 1780 41384
rect 5028 41440 5092 41444
rect 5028 41384 5042 41440
rect 5042 41384 5092 41440
rect 5028 41380 5092 41384
rect 3012 41372 3076 41376
rect 3012 41316 3016 41372
rect 3016 41316 3072 41372
rect 3072 41316 3076 41372
rect 3012 41312 3076 41316
rect 3092 41372 3156 41376
rect 3092 41316 3096 41372
rect 3096 41316 3152 41372
rect 3152 41316 3156 41372
rect 3092 41312 3156 41316
rect 3172 41372 3236 41376
rect 3172 41316 3176 41372
rect 3176 41316 3232 41372
rect 3232 41316 3236 41372
rect 3172 41312 3236 41316
rect 3252 41372 3316 41376
rect 3252 41316 3256 41372
rect 3256 41316 3312 41372
rect 3312 41316 3316 41372
rect 3252 41312 3316 41316
rect 1952 40828 2016 40832
rect 1952 40772 1956 40828
rect 1956 40772 2012 40828
rect 2012 40772 2016 40828
rect 1952 40768 2016 40772
rect 2032 40828 2096 40832
rect 2032 40772 2036 40828
rect 2036 40772 2092 40828
rect 2092 40772 2096 40828
rect 2032 40768 2096 40772
rect 2112 40828 2176 40832
rect 2112 40772 2116 40828
rect 2116 40772 2172 40828
rect 2172 40772 2176 40828
rect 2112 40768 2176 40772
rect 2192 40828 2256 40832
rect 2192 40772 2196 40828
rect 2196 40772 2252 40828
rect 2252 40772 2256 40828
rect 2192 40768 2256 40772
rect 7952 40828 8016 40832
rect 7952 40772 7956 40828
rect 7956 40772 8012 40828
rect 8012 40772 8016 40828
rect 7952 40768 8016 40772
rect 8032 40828 8096 40832
rect 8032 40772 8036 40828
rect 8036 40772 8092 40828
rect 8092 40772 8096 40828
rect 8032 40768 8096 40772
rect 8112 40828 8176 40832
rect 8112 40772 8116 40828
rect 8116 40772 8172 40828
rect 8172 40772 8176 40828
rect 8112 40768 8176 40772
rect 8192 40828 8256 40832
rect 8192 40772 8196 40828
rect 8196 40772 8252 40828
rect 8252 40772 8256 40828
rect 8192 40768 8256 40772
rect 3012 40284 3076 40288
rect 3012 40228 3016 40284
rect 3016 40228 3072 40284
rect 3072 40228 3076 40284
rect 3012 40224 3076 40228
rect 3092 40284 3156 40288
rect 3092 40228 3096 40284
rect 3096 40228 3152 40284
rect 3152 40228 3156 40284
rect 3092 40224 3156 40228
rect 3172 40284 3236 40288
rect 3172 40228 3176 40284
rect 3176 40228 3232 40284
rect 3232 40228 3236 40284
rect 3172 40224 3236 40228
rect 3252 40284 3316 40288
rect 3252 40228 3256 40284
rect 3256 40228 3312 40284
rect 3312 40228 3316 40284
rect 3252 40224 3316 40228
rect 1952 39740 2016 39744
rect 1952 39684 1956 39740
rect 1956 39684 2012 39740
rect 2012 39684 2016 39740
rect 1952 39680 2016 39684
rect 2032 39740 2096 39744
rect 2032 39684 2036 39740
rect 2036 39684 2092 39740
rect 2092 39684 2096 39740
rect 2032 39680 2096 39684
rect 2112 39740 2176 39744
rect 2112 39684 2116 39740
rect 2116 39684 2172 39740
rect 2172 39684 2176 39740
rect 2112 39680 2176 39684
rect 2192 39740 2256 39744
rect 2192 39684 2196 39740
rect 2196 39684 2252 39740
rect 2252 39684 2256 39740
rect 2192 39680 2256 39684
rect 7952 39740 8016 39744
rect 7952 39684 7956 39740
rect 7956 39684 8012 39740
rect 8012 39684 8016 39740
rect 7952 39680 8016 39684
rect 8032 39740 8096 39744
rect 8032 39684 8036 39740
rect 8036 39684 8092 39740
rect 8092 39684 8096 39740
rect 8032 39680 8096 39684
rect 8112 39740 8176 39744
rect 8112 39684 8116 39740
rect 8116 39684 8172 39740
rect 8172 39684 8176 39740
rect 8112 39680 8176 39684
rect 8192 39740 8256 39744
rect 8192 39684 8196 39740
rect 8196 39684 8252 39740
rect 8252 39684 8256 39740
rect 8192 39680 8256 39684
rect 3012 39196 3076 39200
rect 3012 39140 3016 39196
rect 3016 39140 3072 39196
rect 3072 39140 3076 39196
rect 3012 39136 3076 39140
rect 3092 39196 3156 39200
rect 3092 39140 3096 39196
rect 3096 39140 3152 39196
rect 3152 39140 3156 39196
rect 3092 39136 3156 39140
rect 3172 39196 3236 39200
rect 3172 39140 3176 39196
rect 3176 39140 3232 39196
rect 3232 39140 3236 39196
rect 3172 39136 3236 39140
rect 3252 39196 3316 39200
rect 3252 39140 3256 39196
rect 3256 39140 3312 39196
rect 3312 39140 3316 39196
rect 3252 39136 3316 39140
rect 1952 38652 2016 38656
rect 1952 38596 1956 38652
rect 1956 38596 2012 38652
rect 2012 38596 2016 38652
rect 1952 38592 2016 38596
rect 2032 38652 2096 38656
rect 2032 38596 2036 38652
rect 2036 38596 2092 38652
rect 2092 38596 2096 38652
rect 2032 38592 2096 38596
rect 2112 38652 2176 38656
rect 2112 38596 2116 38652
rect 2116 38596 2172 38652
rect 2172 38596 2176 38652
rect 2112 38592 2176 38596
rect 2192 38652 2256 38656
rect 2192 38596 2196 38652
rect 2196 38596 2252 38652
rect 2252 38596 2256 38652
rect 2192 38592 2256 38596
rect 7952 38652 8016 38656
rect 7952 38596 7956 38652
rect 7956 38596 8012 38652
rect 8012 38596 8016 38652
rect 7952 38592 8016 38596
rect 8032 38652 8096 38656
rect 8032 38596 8036 38652
rect 8036 38596 8092 38652
rect 8092 38596 8096 38652
rect 8032 38592 8096 38596
rect 8112 38652 8176 38656
rect 8112 38596 8116 38652
rect 8116 38596 8172 38652
rect 8172 38596 8176 38652
rect 8112 38592 8176 38596
rect 8192 38652 8256 38656
rect 8192 38596 8196 38652
rect 8196 38596 8252 38652
rect 8252 38596 8256 38652
rect 8192 38592 8256 38596
rect 3012 38108 3076 38112
rect 3012 38052 3016 38108
rect 3016 38052 3072 38108
rect 3072 38052 3076 38108
rect 3012 38048 3076 38052
rect 3092 38108 3156 38112
rect 3092 38052 3096 38108
rect 3096 38052 3152 38108
rect 3152 38052 3156 38108
rect 3092 38048 3156 38052
rect 3172 38108 3236 38112
rect 3172 38052 3176 38108
rect 3176 38052 3232 38108
rect 3232 38052 3236 38108
rect 3172 38048 3236 38052
rect 3252 38108 3316 38112
rect 3252 38052 3256 38108
rect 3256 38052 3312 38108
rect 3312 38052 3316 38108
rect 3252 38048 3316 38052
rect 1952 37564 2016 37568
rect 1952 37508 1956 37564
rect 1956 37508 2012 37564
rect 2012 37508 2016 37564
rect 1952 37504 2016 37508
rect 2032 37564 2096 37568
rect 2032 37508 2036 37564
rect 2036 37508 2092 37564
rect 2092 37508 2096 37564
rect 2032 37504 2096 37508
rect 2112 37564 2176 37568
rect 2112 37508 2116 37564
rect 2116 37508 2172 37564
rect 2172 37508 2176 37564
rect 2112 37504 2176 37508
rect 2192 37564 2256 37568
rect 2192 37508 2196 37564
rect 2196 37508 2252 37564
rect 2252 37508 2256 37564
rect 2192 37504 2256 37508
rect 7952 37564 8016 37568
rect 7952 37508 7956 37564
rect 7956 37508 8012 37564
rect 8012 37508 8016 37564
rect 7952 37504 8016 37508
rect 8032 37564 8096 37568
rect 8032 37508 8036 37564
rect 8036 37508 8092 37564
rect 8092 37508 8096 37564
rect 8032 37504 8096 37508
rect 8112 37564 8176 37568
rect 8112 37508 8116 37564
rect 8116 37508 8172 37564
rect 8172 37508 8176 37564
rect 8112 37504 8176 37508
rect 8192 37564 8256 37568
rect 8192 37508 8196 37564
rect 8196 37508 8252 37564
rect 8252 37508 8256 37564
rect 8192 37504 8256 37508
rect 3012 37020 3076 37024
rect 3012 36964 3016 37020
rect 3016 36964 3072 37020
rect 3072 36964 3076 37020
rect 3012 36960 3076 36964
rect 3092 37020 3156 37024
rect 3092 36964 3096 37020
rect 3096 36964 3152 37020
rect 3152 36964 3156 37020
rect 3092 36960 3156 36964
rect 3172 37020 3236 37024
rect 3172 36964 3176 37020
rect 3176 36964 3232 37020
rect 3232 36964 3236 37020
rect 3172 36960 3236 36964
rect 3252 37020 3316 37024
rect 3252 36964 3256 37020
rect 3256 36964 3312 37020
rect 3312 36964 3316 37020
rect 3252 36960 3316 36964
rect 1952 36476 2016 36480
rect 1952 36420 1956 36476
rect 1956 36420 2012 36476
rect 2012 36420 2016 36476
rect 1952 36416 2016 36420
rect 2032 36476 2096 36480
rect 2032 36420 2036 36476
rect 2036 36420 2092 36476
rect 2092 36420 2096 36476
rect 2032 36416 2096 36420
rect 2112 36476 2176 36480
rect 2112 36420 2116 36476
rect 2116 36420 2172 36476
rect 2172 36420 2176 36476
rect 2112 36416 2176 36420
rect 2192 36476 2256 36480
rect 2192 36420 2196 36476
rect 2196 36420 2252 36476
rect 2252 36420 2256 36476
rect 2192 36416 2256 36420
rect 7952 36476 8016 36480
rect 7952 36420 7956 36476
rect 7956 36420 8012 36476
rect 8012 36420 8016 36476
rect 7952 36416 8016 36420
rect 8032 36476 8096 36480
rect 8032 36420 8036 36476
rect 8036 36420 8092 36476
rect 8092 36420 8096 36476
rect 8032 36416 8096 36420
rect 8112 36476 8176 36480
rect 8112 36420 8116 36476
rect 8116 36420 8172 36476
rect 8172 36420 8176 36476
rect 8112 36416 8176 36420
rect 8192 36476 8256 36480
rect 8192 36420 8196 36476
rect 8196 36420 8252 36476
rect 8252 36420 8256 36476
rect 8192 36416 8256 36420
rect 3012 35932 3076 35936
rect 3012 35876 3016 35932
rect 3016 35876 3072 35932
rect 3072 35876 3076 35932
rect 3012 35872 3076 35876
rect 3092 35932 3156 35936
rect 3092 35876 3096 35932
rect 3096 35876 3152 35932
rect 3152 35876 3156 35932
rect 3092 35872 3156 35876
rect 3172 35932 3236 35936
rect 3172 35876 3176 35932
rect 3176 35876 3232 35932
rect 3232 35876 3236 35932
rect 3172 35872 3236 35876
rect 3252 35932 3316 35936
rect 3252 35876 3256 35932
rect 3256 35876 3312 35932
rect 3312 35876 3316 35932
rect 3252 35872 3316 35876
rect 1952 35388 2016 35392
rect 1952 35332 1956 35388
rect 1956 35332 2012 35388
rect 2012 35332 2016 35388
rect 1952 35328 2016 35332
rect 2032 35388 2096 35392
rect 2032 35332 2036 35388
rect 2036 35332 2092 35388
rect 2092 35332 2096 35388
rect 2032 35328 2096 35332
rect 2112 35388 2176 35392
rect 2112 35332 2116 35388
rect 2116 35332 2172 35388
rect 2172 35332 2176 35388
rect 2112 35328 2176 35332
rect 2192 35388 2256 35392
rect 2192 35332 2196 35388
rect 2196 35332 2252 35388
rect 2252 35332 2256 35388
rect 2192 35328 2256 35332
rect 7952 35388 8016 35392
rect 7952 35332 7956 35388
rect 7956 35332 8012 35388
rect 8012 35332 8016 35388
rect 7952 35328 8016 35332
rect 8032 35388 8096 35392
rect 8032 35332 8036 35388
rect 8036 35332 8092 35388
rect 8092 35332 8096 35388
rect 8032 35328 8096 35332
rect 8112 35388 8176 35392
rect 8112 35332 8116 35388
rect 8116 35332 8172 35388
rect 8172 35332 8176 35388
rect 8112 35328 8176 35332
rect 8192 35388 8256 35392
rect 8192 35332 8196 35388
rect 8196 35332 8252 35388
rect 8252 35332 8256 35388
rect 8192 35328 8256 35332
rect 3012 34844 3076 34848
rect 3012 34788 3016 34844
rect 3016 34788 3072 34844
rect 3072 34788 3076 34844
rect 3012 34784 3076 34788
rect 3092 34844 3156 34848
rect 3092 34788 3096 34844
rect 3096 34788 3152 34844
rect 3152 34788 3156 34844
rect 3092 34784 3156 34788
rect 3172 34844 3236 34848
rect 3172 34788 3176 34844
rect 3176 34788 3232 34844
rect 3232 34788 3236 34844
rect 3172 34784 3236 34788
rect 3252 34844 3316 34848
rect 3252 34788 3256 34844
rect 3256 34788 3312 34844
rect 3312 34788 3316 34844
rect 3252 34784 3316 34788
rect 1952 34300 2016 34304
rect 1952 34244 1956 34300
rect 1956 34244 2012 34300
rect 2012 34244 2016 34300
rect 1952 34240 2016 34244
rect 2032 34300 2096 34304
rect 2032 34244 2036 34300
rect 2036 34244 2092 34300
rect 2092 34244 2096 34300
rect 2032 34240 2096 34244
rect 2112 34300 2176 34304
rect 2112 34244 2116 34300
rect 2116 34244 2172 34300
rect 2172 34244 2176 34300
rect 2112 34240 2176 34244
rect 2192 34300 2256 34304
rect 2192 34244 2196 34300
rect 2196 34244 2252 34300
rect 2252 34244 2256 34300
rect 2192 34240 2256 34244
rect 7952 34300 8016 34304
rect 7952 34244 7956 34300
rect 7956 34244 8012 34300
rect 8012 34244 8016 34300
rect 7952 34240 8016 34244
rect 8032 34300 8096 34304
rect 8032 34244 8036 34300
rect 8036 34244 8092 34300
rect 8092 34244 8096 34300
rect 8032 34240 8096 34244
rect 8112 34300 8176 34304
rect 8112 34244 8116 34300
rect 8116 34244 8172 34300
rect 8172 34244 8176 34300
rect 8112 34240 8176 34244
rect 8192 34300 8256 34304
rect 8192 34244 8196 34300
rect 8196 34244 8252 34300
rect 8252 34244 8256 34300
rect 8192 34240 8256 34244
rect 3012 33756 3076 33760
rect 3012 33700 3016 33756
rect 3016 33700 3072 33756
rect 3072 33700 3076 33756
rect 3012 33696 3076 33700
rect 3092 33756 3156 33760
rect 3092 33700 3096 33756
rect 3096 33700 3152 33756
rect 3152 33700 3156 33756
rect 3092 33696 3156 33700
rect 3172 33756 3236 33760
rect 3172 33700 3176 33756
rect 3176 33700 3232 33756
rect 3232 33700 3236 33756
rect 3172 33696 3236 33700
rect 3252 33756 3316 33760
rect 3252 33700 3256 33756
rect 3256 33700 3312 33756
rect 3312 33700 3316 33756
rect 3252 33696 3316 33700
rect 4660 33492 4724 33556
rect 1952 33212 2016 33216
rect 1952 33156 1956 33212
rect 1956 33156 2012 33212
rect 2012 33156 2016 33212
rect 1952 33152 2016 33156
rect 2032 33212 2096 33216
rect 2032 33156 2036 33212
rect 2036 33156 2092 33212
rect 2092 33156 2096 33212
rect 2032 33152 2096 33156
rect 2112 33212 2176 33216
rect 2112 33156 2116 33212
rect 2116 33156 2172 33212
rect 2172 33156 2176 33212
rect 2112 33152 2176 33156
rect 2192 33212 2256 33216
rect 2192 33156 2196 33212
rect 2196 33156 2252 33212
rect 2252 33156 2256 33212
rect 2192 33152 2256 33156
rect 7952 33212 8016 33216
rect 7952 33156 7956 33212
rect 7956 33156 8012 33212
rect 8012 33156 8016 33212
rect 7952 33152 8016 33156
rect 8032 33212 8096 33216
rect 8032 33156 8036 33212
rect 8036 33156 8092 33212
rect 8092 33156 8096 33212
rect 8032 33152 8096 33156
rect 8112 33212 8176 33216
rect 8112 33156 8116 33212
rect 8116 33156 8172 33212
rect 8172 33156 8176 33212
rect 8112 33152 8176 33156
rect 8192 33212 8256 33216
rect 8192 33156 8196 33212
rect 8196 33156 8252 33212
rect 8252 33156 8256 33212
rect 8192 33152 8256 33156
rect 3012 32668 3076 32672
rect 3012 32612 3016 32668
rect 3016 32612 3072 32668
rect 3072 32612 3076 32668
rect 3012 32608 3076 32612
rect 3092 32668 3156 32672
rect 3092 32612 3096 32668
rect 3096 32612 3152 32668
rect 3152 32612 3156 32668
rect 3092 32608 3156 32612
rect 3172 32668 3236 32672
rect 3172 32612 3176 32668
rect 3176 32612 3232 32668
rect 3232 32612 3236 32668
rect 3172 32608 3236 32612
rect 3252 32668 3316 32672
rect 3252 32612 3256 32668
rect 3256 32612 3312 32668
rect 3312 32612 3316 32668
rect 3252 32608 3316 32612
rect 1952 32124 2016 32128
rect 1952 32068 1956 32124
rect 1956 32068 2012 32124
rect 2012 32068 2016 32124
rect 1952 32064 2016 32068
rect 2032 32124 2096 32128
rect 2032 32068 2036 32124
rect 2036 32068 2092 32124
rect 2092 32068 2096 32124
rect 2032 32064 2096 32068
rect 2112 32124 2176 32128
rect 2112 32068 2116 32124
rect 2116 32068 2172 32124
rect 2172 32068 2176 32124
rect 2112 32064 2176 32068
rect 2192 32124 2256 32128
rect 2192 32068 2196 32124
rect 2196 32068 2252 32124
rect 2252 32068 2256 32124
rect 2192 32064 2256 32068
rect 7952 32124 8016 32128
rect 7952 32068 7956 32124
rect 7956 32068 8012 32124
rect 8012 32068 8016 32124
rect 7952 32064 8016 32068
rect 8032 32124 8096 32128
rect 8032 32068 8036 32124
rect 8036 32068 8092 32124
rect 8092 32068 8096 32124
rect 8032 32064 8096 32068
rect 8112 32124 8176 32128
rect 8112 32068 8116 32124
rect 8116 32068 8172 32124
rect 8172 32068 8176 32124
rect 8112 32064 8176 32068
rect 8192 32124 8256 32128
rect 8192 32068 8196 32124
rect 8196 32068 8252 32124
rect 8252 32068 8256 32124
rect 8192 32064 8256 32068
rect 3012 31580 3076 31584
rect 3012 31524 3016 31580
rect 3016 31524 3072 31580
rect 3072 31524 3076 31580
rect 3012 31520 3076 31524
rect 3092 31580 3156 31584
rect 3092 31524 3096 31580
rect 3096 31524 3152 31580
rect 3152 31524 3156 31580
rect 3092 31520 3156 31524
rect 3172 31580 3236 31584
rect 3172 31524 3176 31580
rect 3176 31524 3232 31580
rect 3232 31524 3236 31580
rect 3172 31520 3236 31524
rect 3252 31580 3316 31584
rect 3252 31524 3256 31580
rect 3256 31524 3312 31580
rect 3312 31524 3316 31580
rect 3252 31520 3316 31524
rect 1952 31036 2016 31040
rect 1952 30980 1956 31036
rect 1956 30980 2012 31036
rect 2012 30980 2016 31036
rect 1952 30976 2016 30980
rect 2032 31036 2096 31040
rect 2032 30980 2036 31036
rect 2036 30980 2092 31036
rect 2092 30980 2096 31036
rect 2032 30976 2096 30980
rect 2112 31036 2176 31040
rect 2112 30980 2116 31036
rect 2116 30980 2172 31036
rect 2172 30980 2176 31036
rect 2112 30976 2176 30980
rect 2192 31036 2256 31040
rect 2192 30980 2196 31036
rect 2196 30980 2252 31036
rect 2252 30980 2256 31036
rect 2192 30976 2256 30980
rect 7952 31036 8016 31040
rect 7952 30980 7956 31036
rect 7956 30980 8012 31036
rect 8012 30980 8016 31036
rect 7952 30976 8016 30980
rect 8032 31036 8096 31040
rect 8032 30980 8036 31036
rect 8036 30980 8092 31036
rect 8092 30980 8096 31036
rect 8032 30976 8096 30980
rect 8112 31036 8176 31040
rect 8112 30980 8116 31036
rect 8116 30980 8172 31036
rect 8172 30980 8176 31036
rect 8112 30976 8176 30980
rect 8192 31036 8256 31040
rect 8192 30980 8196 31036
rect 8196 30980 8252 31036
rect 8252 30980 8256 31036
rect 8192 30976 8256 30980
rect 3012 30492 3076 30496
rect 3012 30436 3016 30492
rect 3016 30436 3072 30492
rect 3072 30436 3076 30492
rect 3012 30432 3076 30436
rect 3092 30492 3156 30496
rect 3092 30436 3096 30492
rect 3096 30436 3152 30492
rect 3152 30436 3156 30492
rect 3092 30432 3156 30436
rect 3172 30492 3236 30496
rect 3172 30436 3176 30492
rect 3176 30436 3232 30492
rect 3232 30436 3236 30492
rect 3172 30432 3236 30436
rect 3252 30492 3316 30496
rect 3252 30436 3256 30492
rect 3256 30436 3312 30492
rect 3312 30436 3316 30492
rect 3252 30432 3316 30436
rect 1952 29948 2016 29952
rect 1952 29892 1956 29948
rect 1956 29892 2012 29948
rect 2012 29892 2016 29948
rect 1952 29888 2016 29892
rect 2032 29948 2096 29952
rect 2032 29892 2036 29948
rect 2036 29892 2092 29948
rect 2092 29892 2096 29948
rect 2032 29888 2096 29892
rect 2112 29948 2176 29952
rect 2112 29892 2116 29948
rect 2116 29892 2172 29948
rect 2172 29892 2176 29948
rect 2112 29888 2176 29892
rect 2192 29948 2256 29952
rect 2192 29892 2196 29948
rect 2196 29892 2252 29948
rect 2252 29892 2256 29948
rect 2192 29888 2256 29892
rect 7952 29948 8016 29952
rect 7952 29892 7956 29948
rect 7956 29892 8012 29948
rect 8012 29892 8016 29948
rect 7952 29888 8016 29892
rect 8032 29948 8096 29952
rect 8032 29892 8036 29948
rect 8036 29892 8092 29948
rect 8092 29892 8096 29948
rect 8032 29888 8096 29892
rect 8112 29948 8176 29952
rect 8112 29892 8116 29948
rect 8116 29892 8172 29948
rect 8172 29892 8176 29948
rect 8112 29888 8176 29892
rect 8192 29948 8256 29952
rect 8192 29892 8196 29948
rect 8196 29892 8252 29948
rect 8252 29892 8256 29948
rect 8192 29888 8256 29892
rect 3012 29404 3076 29408
rect 3012 29348 3016 29404
rect 3016 29348 3072 29404
rect 3072 29348 3076 29404
rect 3012 29344 3076 29348
rect 3092 29404 3156 29408
rect 3092 29348 3096 29404
rect 3096 29348 3152 29404
rect 3152 29348 3156 29404
rect 3092 29344 3156 29348
rect 3172 29404 3236 29408
rect 3172 29348 3176 29404
rect 3176 29348 3232 29404
rect 3232 29348 3236 29404
rect 3172 29344 3236 29348
rect 3252 29404 3316 29408
rect 3252 29348 3256 29404
rect 3256 29348 3312 29404
rect 3312 29348 3316 29404
rect 3252 29344 3316 29348
rect 3924 29004 3988 29068
rect 1952 28860 2016 28864
rect 1952 28804 1956 28860
rect 1956 28804 2012 28860
rect 2012 28804 2016 28860
rect 1952 28800 2016 28804
rect 2032 28860 2096 28864
rect 2032 28804 2036 28860
rect 2036 28804 2092 28860
rect 2092 28804 2096 28860
rect 2032 28800 2096 28804
rect 2112 28860 2176 28864
rect 2112 28804 2116 28860
rect 2116 28804 2172 28860
rect 2172 28804 2176 28860
rect 2112 28800 2176 28804
rect 2192 28860 2256 28864
rect 2192 28804 2196 28860
rect 2196 28804 2252 28860
rect 2252 28804 2256 28860
rect 2192 28800 2256 28804
rect 7952 28860 8016 28864
rect 7952 28804 7956 28860
rect 7956 28804 8012 28860
rect 8012 28804 8016 28860
rect 7952 28800 8016 28804
rect 8032 28860 8096 28864
rect 8032 28804 8036 28860
rect 8036 28804 8092 28860
rect 8092 28804 8096 28860
rect 8032 28800 8096 28804
rect 8112 28860 8176 28864
rect 8112 28804 8116 28860
rect 8116 28804 8172 28860
rect 8172 28804 8176 28860
rect 8112 28800 8176 28804
rect 8192 28860 8256 28864
rect 8192 28804 8196 28860
rect 8196 28804 8252 28860
rect 8252 28804 8256 28860
rect 8192 28800 8256 28804
rect 3012 28316 3076 28320
rect 3012 28260 3016 28316
rect 3016 28260 3072 28316
rect 3072 28260 3076 28316
rect 3012 28256 3076 28260
rect 3092 28316 3156 28320
rect 3092 28260 3096 28316
rect 3096 28260 3152 28316
rect 3152 28260 3156 28316
rect 3092 28256 3156 28260
rect 3172 28316 3236 28320
rect 3172 28260 3176 28316
rect 3176 28260 3232 28316
rect 3232 28260 3236 28316
rect 3172 28256 3236 28260
rect 3252 28316 3316 28320
rect 3252 28260 3256 28316
rect 3256 28260 3312 28316
rect 3312 28260 3316 28316
rect 3252 28256 3316 28260
rect 1952 27772 2016 27776
rect 1952 27716 1956 27772
rect 1956 27716 2012 27772
rect 2012 27716 2016 27772
rect 1952 27712 2016 27716
rect 2032 27772 2096 27776
rect 2032 27716 2036 27772
rect 2036 27716 2092 27772
rect 2092 27716 2096 27772
rect 2032 27712 2096 27716
rect 2112 27772 2176 27776
rect 2112 27716 2116 27772
rect 2116 27716 2172 27772
rect 2172 27716 2176 27772
rect 2112 27712 2176 27716
rect 2192 27772 2256 27776
rect 2192 27716 2196 27772
rect 2196 27716 2252 27772
rect 2252 27716 2256 27772
rect 2192 27712 2256 27716
rect 7952 27772 8016 27776
rect 7952 27716 7956 27772
rect 7956 27716 8012 27772
rect 8012 27716 8016 27772
rect 7952 27712 8016 27716
rect 8032 27772 8096 27776
rect 8032 27716 8036 27772
rect 8036 27716 8092 27772
rect 8092 27716 8096 27772
rect 8032 27712 8096 27716
rect 8112 27772 8176 27776
rect 8112 27716 8116 27772
rect 8116 27716 8172 27772
rect 8172 27716 8176 27772
rect 8112 27712 8176 27716
rect 8192 27772 8256 27776
rect 8192 27716 8196 27772
rect 8196 27716 8252 27772
rect 8252 27716 8256 27772
rect 8192 27712 8256 27716
rect 3012 27228 3076 27232
rect 3012 27172 3016 27228
rect 3016 27172 3072 27228
rect 3072 27172 3076 27228
rect 3012 27168 3076 27172
rect 3092 27228 3156 27232
rect 3092 27172 3096 27228
rect 3096 27172 3152 27228
rect 3152 27172 3156 27228
rect 3092 27168 3156 27172
rect 3172 27228 3236 27232
rect 3172 27172 3176 27228
rect 3176 27172 3232 27228
rect 3232 27172 3236 27228
rect 3172 27168 3236 27172
rect 3252 27228 3316 27232
rect 3252 27172 3256 27228
rect 3256 27172 3312 27228
rect 3312 27172 3316 27228
rect 3252 27168 3316 27172
rect 1952 26684 2016 26688
rect 1952 26628 1956 26684
rect 1956 26628 2012 26684
rect 2012 26628 2016 26684
rect 1952 26624 2016 26628
rect 2032 26684 2096 26688
rect 2032 26628 2036 26684
rect 2036 26628 2092 26684
rect 2092 26628 2096 26684
rect 2032 26624 2096 26628
rect 2112 26684 2176 26688
rect 2112 26628 2116 26684
rect 2116 26628 2172 26684
rect 2172 26628 2176 26684
rect 2112 26624 2176 26628
rect 2192 26684 2256 26688
rect 2192 26628 2196 26684
rect 2196 26628 2252 26684
rect 2252 26628 2256 26684
rect 2192 26624 2256 26628
rect 7952 26684 8016 26688
rect 7952 26628 7956 26684
rect 7956 26628 8012 26684
rect 8012 26628 8016 26684
rect 7952 26624 8016 26628
rect 8032 26684 8096 26688
rect 8032 26628 8036 26684
rect 8036 26628 8092 26684
rect 8092 26628 8096 26684
rect 8032 26624 8096 26628
rect 8112 26684 8176 26688
rect 8112 26628 8116 26684
rect 8116 26628 8172 26684
rect 8172 26628 8176 26684
rect 8112 26624 8176 26628
rect 8192 26684 8256 26688
rect 8192 26628 8196 26684
rect 8196 26628 8252 26684
rect 8252 26628 8256 26684
rect 8192 26624 8256 26628
rect 7604 26284 7668 26348
rect 3012 26140 3076 26144
rect 3012 26084 3016 26140
rect 3016 26084 3072 26140
rect 3072 26084 3076 26140
rect 3012 26080 3076 26084
rect 3092 26140 3156 26144
rect 3092 26084 3096 26140
rect 3096 26084 3152 26140
rect 3152 26084 3156 26140
rect 3092 26080 3156 26084
rect 3172 26140 3236 26144
rect 3172 26084 3176 26140
rect 3176 26084 3232 26140
rect 3232 26084 3236 26140
rect 3172 26080 3236 26084
rect 3252 26140 3316 26144
rect 3252 26084 3256 26140
rect 3256 26084 3312 26140
rect 3312 26084 3316 26140
rect 3252 26080 3316 26084
rect 1952 25596 2016 25600
rect 1952 25540 1956 25596
rect 1956 25540 2012 25596
rect 2012 25540 2016 25596
rect 1952 25536 2016 25540
rect 2032 25596 2096 25600
rect 2032 25540 2036 25596
rect 2036 25540 2092 25596
rect 2092 25540 2096 25596
rect 2032 25536 2096 25540
rect 2112 25596 2176 25600
rect 2112 25540 2116 25596
rect 2116 25540 2172 25596
rect 2172 25540 2176 25596
rect 2112 25536 2176 25540
rect 2192 25596 2256 25600
rect 2192 25540 2196 25596
rect 2196 25540 2252 25596
rect 2252 25540 2256 25596
rect 2192 25536 2256 25540
rect 7952 25596 8016 25600
rect 7952 25540 7956 25596
rect 7956 25540 8012 25596
rect 8012 25540 8016 25596
rect 7952 25536 8016 25540
rect 8032 25596 8096 25600
rect 8032 25540 8036 25596
rect 8036 25540 8092 25596
rect 8092 25540 8096 25596
rect 8032 25536 8096 25540
rect 8112 25596 8176 25600
rect 8112 25540 8116 25596
rect 8116 25540 8172 25596
rect 8172 25540 8176 25596
rect 8112 25536 8176 25540
rect 8192 25596 8256 25600
rect 8192 25540 8196 25596
rect 8196 25540 8252 25596
rect 8252 25540 8256 25596
rect 8192 25536 8256 25540
rect 3556 25196 3620 25260
rect 3012 25052 3076 25056
rect 3012 24996 3016 25052
rect 3016 24996 3072 25052
rect 3072 24996 3076 25052
rect 3012 24992 3076 24996
rect 3092 25052 3156 25056
rect 3092 24996 3096 25052
rect 3096 24996 3152 25052
rect 3152 24996 3156 25052
rect 3092 24992 3156 24996
rect 3172 25052 3236 25056
rect 3172 24996 3176 25052
rect 3176 24996 3232 25052
rect 3232 24996 3236 25052
rect 3172 24992 3236 24996
rect 3252 25052 3316 25056
rect 3252 24996 3256 25052
rect 3256 24996 3312 25052
rect 3312 24996 3316 25052
rect 3252 24992 3316 24996
rect 7236 24788 7300 24852
rect 1952 24508 2016 24512
rect 1952 24452 1956 24508
rect 1956 24452 2012 24508
rect 2012 24452 2016 24508
rect 1952 24448 2016 24452
rect 2032 24508 2096 24512
rect 2032 24452 2036 24508
rect 2036 24452 2092 24508
rect 2092 24452 2096 24508
rect 2032 24448 2096 24452
rect 2112 24508 2176 24512
rect 2112 24452 2116 24508
rect 2116 24452 2172 24508
rect 2172 24452 2176 24508
rect 2112 24448 2176 24452
rect 2192 24508 2256 24512
rect 2192 24452 2196 24508
rect 2196 24452 2252 24508
rect 2252 24452 2256 24508
rect 2192 24448 2256 24452
rect 7952 24508 8016 24512
rect 7952 24452 7956 24508
rect 7956 24452 8012 24508
rect 8012 24452 8016 24508
rect 7952 24448 8016 24452
rect 8032 24508 8096 24512
rect 8032 24452 8036 24508
rect 8036 24452 8092 24508
rect 8092 24452 8096 24508
rect 8032 24448 8096 24452
rect 8112 24508 8176 24512
rect 8112 24452 8116 24508
rect 8116 24452 8172 24508
rect 8172 24452 8176 24508
rect 8112 24448 8176 24452
rect 8192 24508 8256 24512
rect 8192 24452 8196 24508
rect 8196 24452 8252 24508
rect 8252 24452 8256 24508
rect 8192 24448 8256 24452
rect 5396 23972 5460 24036
rect 3012 23964 3076 23968
rect 3012 23908 3016 23964
rect 3016 23908 3072 23964
rect 3072 23908 3076 23964
rect 3012 23904 3076 23908
rect 3092 23964 3156 23968
rect 3092 23908 3096 23964
rect 3096 23908 3152 23964
rect 3152 23908 3156 23964
rect 3092 23904 3156 23908
rect 3172 23964 3236 23968
rect 3172 23908 3176 23964
rect 3176 23908 3232 23964
rect 3232 23908 3236 23964
rect 3172 23904 3236 23908
rect 3252 23964 3316 23968
rect 3252 23908 3256 23964
rect 3256 23908 3312 23964
rect 3312 23908 3316 23964
rect 3252 23904 3316 23908
rect 3740 23488 3804 23492
rect 3740 23432 3754 23488
rect 3754 23432 3804 23488
rect 3740 23428 3804 23432
rect 5212 23428 5276 23492
rect 6500 23428 6564 23492
rect 1952 23420 2016 23424
rect 1952 23364 1956 23420
rect 1956 23364 2012 23420
rect 2012 23364 2016 23420
rect 1952 23360 2016 23364
rect 2032 23420 2096 23424
rect 2032 23364 2036 23420
rect 2036 23364 2092 23420
rect 2092 23364 2096 23420
rect 2032 23360 2096 23364
rect 2112 23420 2176 23424
rect 2112 23364 2116 23420
rect 2116 23364 2172 23420
rect 2172 23364 2176 23420
rect 2112 23360 2176 23364
rect 2192 23420 2256 23424
rect 2192 23364 2196 23420
rect 2196 23364 2252 23420
rect 2252 23364 2256 23420
rect 2192 23360 2256 23364
rect 7952 23420 8016 23424
rect 7952 23364 7956 23420
rect 7956 23364 8012 23420
rect 8012 23364 8016 23420
rect 7952 23360 8016 23364
rect 8032 23420 8096 23424
rect 8032 23364 8036 23420
rect 8036 23364 8092 23420
rect 8092 23364 8096 23420
rect 8032 23360 8096 23364
rect 8112 23420 8176 23424
rect 8112 23364 8116 23420
rect 8116 23364 8172 23420
rect 8172 23364 8176 23420
rect 8112 23360 8176 23364
rect 8192 23420 8256 23424
rect 8192 23364 8196 23420
rect 8196 23364 8252 23420
rect 8252 23364 8256 23420
rect 8192 23360 8256 23364
rect 3012 22876 3076 22880
rect 3012 22820 3016 22876
rect 3016 22820 3072 22876
rect 3072 22820 3076 22876
rect 3012 22816 3076 22820
rect 3092 22876 3156 22880
rect 3092 22820 3096 22876
rect 3096 22820 3152 22876
rect 3152 22820 3156 22876
rect 3092 22816 3156 22820
rect 3172 22876 3236 22880
rect 3172 22820 3176 22876
rect 3176 22820 3232 22876
rect 3232 22820 3236 22876
rect 3172 22816 3236 22820
rect 3252 22876 3316 22880
rect 3252 22820 3256 22876
rect 3256 22820 3312 22876
rect 3312 22820 3316 22876
rect 3252 22816 3316 22820
rect 9444 22748 9508 22812
rect 7420 22476 7484 22540
rect 9444 22476 9508 22540
rect 1952 22332 2016 22336
rect 1952 22276 1956 22332
rect 1956 22276 2012 22332
rect 2012 22276 2016 22332
rect 1952 22272 2016 22276
rect 2032 22332 2096 22336
rect 2032 22276 2036 22332
rect 2036 22276 2092 22332
rect 2092 22276 2096 22332
rect 2032 22272 2096 22276
rect 2112 22332 2176 22336
rect 2112 22276 2116 22332
rect 2116 22276 2172 22332
rect 2172 22276 2176 22332
rect 2112 22272 2176 22276
rect 2192 22332 2256 22336
rect 2192 22276 2196 22332
rect 2196 22276 2252 22332
rect 2252 22276 2256 22332
rect 2192 22272 2256 22276
rect 7952 22332 8016 22336
rect 7952 22276 7956 22332
rect 7956 22276 8012 22332
rect 8012 22276 8016 22332
rect 7952 22272 8016 22276
rect 8032 22332 8096 22336
rect 8032 22276 8036 22332
rect 8036 22276 8092 22332
rect 8092 22276 8096 22332
rect 8032 22272 8096 22276
rect 8112 22332 8176 22336
rect 8112 22276 8116 22332
rect 8116 22276 8172 22332
rect 8172 22276 8176 22332
rect 8112 22272 8176 22276
rect 8192 22332 8256 22336
rect 8192 22276 8196 22332
rect 8196 22276 8252 22332
rect 8252 22276 8256 22332
rect 8192 22272 8256 22276
rect 7236 22128 7300 22132
rect 7236 22072 7286 22128
rect 7286 22072 7300 22128
rect 7236 22068 7300 22072
rect 3012 21788 3076 21792
rect 3012 21732 3016 21788
rect 3016 21732 3072 21788
rect 3072 21732 3076 21788
rect 3012 21728 3076 21732
rect 3092 21788 3156 21792
rect 3092 21732 3096 21788
rect 3096 21732 3152 21788
rect 3152 21732 3156 21788
rect 3092 21728 3156 21732
rect 3172 21788 3236 21792
rect 3172 21732 3176 21788
rect 3176 21732 3232 21788
rect 3232 21732 3236 21788
rect 3172 21728 3236 21732
rect 3252 21788 3316 21792
rect 3252 21732 3256 21788
rect 3256 21732 3312 21788
rect 3312 21732 3316 21788
rect 3252 21728 3316 21732
rect 8340 21388 8404 21452
rect 1952 21244 2016 21248
rect 1952 21188 1956 21244
rect 1956 21188 2012 21244
rect 2012 21188 2016 21244
rect 1952 21184 2016 21188
rect 2032 21244 2096 21248
rect 2032 21188 2036 21244
rect 2036 21188 2092 21244
rect 2092 21188 2096 21244
rect 2032 21184 2096 21188
rect 2112 21244 2176 21248
rect 2112 21188 2116 21244
rect 2116 21188 2172 21244
rect 2172 21188 2176 21244
rect 2112 21184 2176 21188
rect 2192 21244 2256 21248
rect 2192 21188 2196 21244
rect 2196 21188 2252 21244
rect 2252 21188 2256 21244
rect 2192 21184 2256 21188
rect 7952 21244 8016 21248
rect 7952 21188 7956 21244
rect 7956 21188 8012 21244
rect 8012 21188 8016 21244
rect 7952 21184 8016 21188
rect 8032 21244 8096 21248
rect 8032 21188 8036 21244
rect 8036 21188 8092 21244
rect 8092 21188 8096 21244
rect 8032 21184 8096 21188
rect 8112 21244 8176 21248
rect 8112 21188 8116 21244
rect 8116 21188 8172 21244
rect 8172 21188 8176 21244
rect 8112 21184 8176 21188
rect 8192 21244 8256 21248
rect 8192 21188 8196 21244
rect 8196 21188 8252 21244
rect 8252 21188 8256 21244
rect 8192 21184 8256 21188
rect 6684 21040 6748 21044
rect 6684 20984 6734 21040
rect 6734 20984 6748 21040
rect 6684 20980 6748 20984
rect 6132 20844 6196 20908
rect 6316 20708 6380 20772
rect 3012 20700 3076 20704
rect 3012 20644 3016 20700
rect 3016 20644 3072 20700
rect 3072 20644 3076 20700
rect 3012 20640 3076 20644
rect 3092 20700 3156 20704
rect 3092 20644 3096 20700
rect 3096 20644 3152 20700
rect 3152 20644 3156 20700
rect 3092 20640 3156 20644
rect 3172 20700 3236 20704
rect 3172 20644 3176 20700
rect 3176 20644 3232 20700
rect 3232 20644 3236 20700
rect 3172 20640 3236 20644
rect 3252 20700 3316 20704
rect 3252 20644 3256 20700
rect 3256 20644 3312 20700
rect 3312 20644 3316 20700
rect 3252 20640 3316 20644
rect 9260 20572 9324 20636
rect 8708 20436 8772 20500
rect 7236 20300 7300 20364
rect 1952 20156 2016 20160
rect 1952 20100 1956 20156
rect 1956 20100 2012 20156
rect 2012 20100 2016 20156
rect 1952 20096 2016 20100
rect 2032 20156 2096 20160
rect 2032 20100 2036 20156
rect 2036 20100 2092 20156
rect 2092 20100 2096 20156
rect 2032 20096 2096 20100
rect 2112 20156 2176 20160
rect 2112 20100 2116 20156
rect 2116 20100 2172 20156
rect 2172 20100 2176 20156
rect 2112 20096 2176 20100
rect 2192 20156 2256 20160
rect 2192 20100 2196 20156
rect 2196 20100 2252 20156
rect 2252 20100 2256 20156
rect 2192 20096 2256 20100
rect 7952 20156 8016 20160
rect 7952 20100 7956 20156
rect 7956 20100 8012 20156
rect 8012 20100 8016 20156
rect 7952 20096 8016 20100
rect 8032 20156 8096 20160
rect 8032 20100 8036 20156
rect 8036 20100 8092 20156
rect 8092 20100 8096 20156
rect 8032 20096 8096 20100
rect 8112 20156 8176 20160
rect 8112 20100 8116 20156
rect 8116 20100 8172 20156
rect 8172 20100 8176 20156
rect 8112 20096 8176 20100
rect 8192 20156 8256 20160
rect 8192 20100 8196 20156
rect 8196 20100 8252 20156
rect 8252 20100 8256 20156
rect 8192 20096 8256 20100
rect 3012 19612 3076 19616
rect 3012 19556 3016 19612
rect 3016 19556 3072 19612
rect 3072 19556 3076 19612
rect 3012 19552 3076 19556
rect 3092 19612 3156 19616
rect 3092 19556 3096 19612
rect 3096 19556 3152 19612
rect 3152 19556 3156 19612
rect 3092 19552 3156 19556
rect 3172 19612 3236 19616
rect 3172 19556 3176 19612
rect 3176 19556 3232 19612
rect 3232 19556 3236 19612
rect 3172 19552 3236 19556
rect 3252 19612 3316 19616
rect 3252 19556 3256 19612
rect 3256 19556 3312 19612
rect 3312 19556 3316 19612
rect 3252 19552 3316 19556
rect 3924 19484 3988 19548
rect 1952 19068 2016 19072
rect 1952 19012 1956 19068
rect 1956 19012 2012 19068
rect 2012 19012 2016 19068
rect 1952 19008 2016 19012
rect 2032 19068 2096 19072
rect 2032 19012 2036 19068
rect 2036 19012 2092 19068
rect 2092 19012 2096 19068
rect 2032 19008 2096 19012
rect 2112 19068 2176 19072
rect 2112 19012 2116 19068
rect 2116 19012 2172 19068
rect 2172 19012 2176 19068
rect 2112 19008 2176 19012
rect 2192 19068 2256 19072
rect 2192 19012 2196 19068
rect 2196 19012 2252 19068
rect 2252 19012 2256 19068
rect 2192 19008 2256 19012
rect 7952 19068 8016 19072
rect 7952 19012 7956 19068
rect 7956 19012 8012 19068
rect 8012 19012 8016 19068
rect 7952 19008 8016 19012
rect 8032 19068 8096 19072
rect 8032 19012 8036 19068
rect 8036 19012 8092 19068
rect 8092 19012 8096 19068
rect 8032 19008 8096 19012
rect 8112 19068 8176 19072
rect 8112 19012 8116 19068
rect 8116 19012 8172 19068
rect 8172 19012 8176 19068
rect 8112 19008 8176 19012
rect 8192 19068 8256 19072
rect 8192 19012 8196 19068
rect 8196 19012 8252 19068
rect 8252 19012 8256 19068
rect 8192 19008 8256 19012
rect 3012 18524 3076 18528
rect 3012 18468 3016 18524
rect 3016 18468 3072 18524
rect 3072 18468 3076 18524
rect 3012 18464 3076 18468
rect 3092 18524 3156 18528
rect 3092 18468 3096 18524
rect 3096 18468 3152 18524
rect 3152 18468 3156 18524
rect 3092 18464 3156 18468
rect 3172 18524 3236 18528
rect 3172 18468 3176 18524
rect 3176 18468 3232 18524
rect 3232 18468 3236 18524
rect 3172 18464 3236 18468
rect 3252 18524 3316 18528
rect 3252 18468 3256 18524
rect 3256 18468 3312 18524
rect 3312 18468 3316 18524
rect 3252 18464 3316 18468
rect 1952 17980 2016 17984
rect 1952 17924 1956 17980
rect 1956 17924 2012 17980
rect 2012 17924 2016 17980
rect 1952 17920 2016 17924
rect 2032 17980 2096 17984
rect 2032 17924 2036 17980
rect 2036 17924 2092 17980
rect 2092 17924 2096 17980
rect 2032 17920 2096 17924
rect 2112 17980 2176 17984
rect 2112 17924 2116 17980
rect 2116 17924 2172 17980
rect 2172 17924 2176 17980
rect 2112 17920 2176 17924
rect 2192 17980 2256 17984
rect 2192 17924 2196 17980
rect 2196 17924 2252 17980
rect 2252 17924 2256 17980
rect 2192 17920 2256 17924
rect 7952 17980 8016 17984
rect 7952 17924 7956 17980
rect 7956 17924 8012 17980
rect 8012 17924 8016 17980
rect 7952 17920 8016 17924
rect 8032 17980 8096 17984
rect 8032 17924 8036 17980
rect 8036 17924 8092 17980
rect 8092 17924 8096 17980
rect 8032 17920 8096 17924
rect 8112 17980 8176 17984
rect 8112 17924 8116 17980
rect 8116 17924 8172 17980
rect 8172 17924 8176 17980
rect 8112 17920 8176 17924
rect 8192 17980 8256 17984
rect 8192 17924 8196 17980
rect 8196 17924 8252 17980
rect 8252 17924 8256 17980
rect 8192 17920 8256 17924
rect 7420 17852 7484 17916
rect 8340 17640 8404 17644
rect 8340 17584 8390 17640
rect 8390 17584 8404 17640
rect 8340 17580 8404 17584
rect 3012 17436 3076 17440
rect 3012 17380 3016 17436
rect 3016 17380 3072 17436
rect 3072 17380 3076 17436
rect 3012 17376 3076 17380
rect 3092 17436 3156 17440
rect 3092 17380 3096 17436
rect 3096 17380 3152 17436
rect 3152 17380 3156 17436
rect 3092 17376 3156 17380
rect 3172 17436 3236 17440
rect 3172 17380 3176 17436
rect 3176 17380 3232 17436
rect 3232 17380 3236 17436
rect 3172 17376 3236 17380
rect 3252 17436 3316 17440
rect 3252 17380 3256 17436
rect 3256 17380 3312 17436
rect 3312 17380 3316 17436
rect 3252 17376 3316 17380
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 7952 16892 8016 16896
rect 7952 16836 7956 16892
rect 7956 16836 8012 16892
rect 8012 16836 8016 16892
rect 7952 16832 8016 16836
rect 8032 16892 8096 16896
rect 8032 16836 8036 16892
rect 8036 16836 8092 16892
rect 8092 16836 8096 16892
rect 8032 16832 8096 16836
rect 8112 16892 8176 16896
rect 8112 16836 8116 16892
rect 8116 16836 8172 16892
rect 8172 16836 8176 16892
rect 8112 16832 8176 16836
rect 8192 16892 8256 16896
rect 8192 16836 8196 16892
rect 8196 16836 8252 16892
rect 8252 16836 8256 16892
rect 8192 16832 8256 16836
rect 3012 16348 3076 16352
rect 3012 16292 3016 16348
rect 3016 16292 3072 16348
rect 3072 16292 3076 16348
rect 3012 16288 3076 16292
rect 3092 16348 3156 16352
rect 3092 16292 3096 16348
rect 3096 16292 3152 16348
rect 3152 16292 3156 16348
rect 3092 16288 3156 16292
rect 3172 16348 3236 16352
rect 3172 16292 3176 16348
rect 3176 16292 3232 16348
rect 3232 16292 3236 16348
rect 3172 16288 3236 16292
rect 3252 16348 3316 16352
rect 3252 16292 3256 16348
rect 3256 16292 3312 16348
rect 3312 16292 3316 16348
rect 3252 16288 3316 16292
rect 1532 16220 1596 16284
rect 5028 16220 5092 16284
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 7952 15804 8016 15808
rect 7952 15748 7956 15804
rect 7956 15748 8012 15804
rect 8012 15748 8016 15804
rect 7952 15744 8016 15748
rect 8032 15804 8096 15808
rect 8032 15748 8036 15804
rect 8036 15748 8092 15804
rect 8092 15748 8096 15804
rect 8032 15744 8096 15748
rect 8112 15804 8176 15808
rect 8112 15748 8116 15804
rect 8116 15748 8172 15804
rect 8172 15748 8176 15804
rect 8112 15744 8176 15748
rect 8192 15804 8256 15808
rect 8192 15748 8196 15804
rect 8196 15748 8252 15804
rect 8252 15748 8256 15804
rect 8192 15744 8256 15748
rect 7236 15404 7300 15468
rect 7604 15404 7668 15468
rect 3012 15260 3076 15264
rect 3012 15204 3016 15260
rect 3016 15204 3072 15260
rect 3072 15204 3076 15260
rect 3012 15200 3076 15204
rect 3092 15260 3156 15264
rect 3092 15204 3096 15260
rect 3096 15204 3152 15260
rect 3152 15204 3156 15260
rect 3092 15200 3156 15204
rect 3172 15260 3236 15264
rect 3172 15204 3176 15260
rect 3176 15204 3232 15260
rect 3232 15204 3236 15260
rect 3172 15200 3236 15204
rect 3252 15260 3316 15264
rect 3252 15204 3256 15260
rect 3256 15204 3312 15260
rect 3312 15204 3316 15260
rect 3252 15200 3316 15204
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 7952 14716 8016 14720
rect 7952 14660 7956 14716
rect 7956 14660 8012 14716
rect 8012 14660 8016 14716
rect 7952 14656 8016 14660
rect 8032 14716 8096 14720
rect 8032 14660 8036 14716
rect 8036 14660 8092 14716
rect 8092 14660 8096 14716
rect 8032 14656 8096 14660
rect 8112 14716 8176 14720
rect 8112 14660 8116 14716
rect 8116 14660 8172 14716
rect 8172 14660 8176 14716
rect 8112 14656 8176 14660
rect 8192 14716 8256 14720
rect 8192 14660 8196 14716
rect 8196 14660 8252 14716
rect 8252 14660 8256 14716
rect 8192 14656 8256 14660
rect 3012 14172 3076 14176
rect 3012 14116 3016 14172
rect 3016 14116 3072 14172
rect 3072 14116 3076 14172
rect 3012 14112 3076 14116
rect 3092 14172 3156 14176
rect 3092 14116 3096 14172
rect 3096 14116 3152 14172
rect 3152 14116 3156 14172
rect 3092 14112 3156 14116
rect 3172 14172 3236 14176
rect 3172 14116 3176 14172
rect 3176 14116 3232 14172
rect 3232 14116 3236 14172
rect 3172 14112 3236 14116
rect 3252 14172 3316 14176
rect 3252 14116 3256 14172
rect 3256 14116 3312 14172
rect 3312 14116 3316 14172
rect 3252 14112 3316 14116
rect 4660 13772 4724 13836
rect 6132 13832 6196 13836
rect 6132 13776 6182 13832
rect 6182 13776 6196 13832
rect 6132 13772 6196 13776
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 7952 13628 8016 13632
rect 7952 13572 7956 13628
rect 7956 13572 8012 13628
rect 8012 13572 8016 13628
rect 7952 13568 8016 13572
rect 8032 13628 8096 13632
rect 8032 13572 8036 13628
rect 8036 13572 8092 13628
rect 8092 13572 8096 13628
rect 8032 13568 8096 13572
rect 8112 13628 8176 13632
rect 8112 13572 8116 13628
rect 8116 13572 8172 13628
rect 8172 13572 8176 13628
rect 8112 13568 8176 13572
rect 8192 13628 8256 13632
rect 8192 13572 8196 13628
rect 8196 13572 8252 13628
rect 8252 13572 8256 13628
rect 8192 13568 8256 13572
rect 3012 13084 3076 13088
rect 3012 13028 3016 13084
rect 3016 13028 3072 13084
rect 3072 13028 3076 13084
rect 3012 13024 3076 13028
rect 3092 13084 3156 13088
rect 3092 13028 3096 13084
rect 3096 13028 3152 13084
rect 3152 13028 3156 13084
rect 3092 13024 3156 13028
rect 3172 13084 3236 13088
rect 3172 13028 3176 13084
rect 3176 13028 3232 13084
rect 3232 13028 3236 13084
rect 3172 13024 3236 13028
rect 3252 13084 3316 13088
rect 3252 13028 3256 13084
rect 3256 13028 3312 13084
rect 3312 13028 3316 13084
rect 3252 13024 3316 13028
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 7952 12540 8016 12544
rect 7952 12484 7956 12540
rect 7956 12484 8012 12540
rect 8012 12484 8016 12540
rect 7952 12480 8016 12484
rect 8032 12540 8096 12544
rect 8032 12484 8036 12540
rect 8036 12484 8092 12540
rect 8092 12484 8096 12540
rect 8032 12480 8096 12484
rect 8112 12540 8176 12544
rect 8112 12484 8116 12540
rect 8116 12484 8172 12540
rect 8172 12484 8176 12540
rect 8112 12480 8176 12484
rect 8192 12540 8256 12544
rect 8192 12484 8196 12540
rect 8196 12484 8252 12540
rect 8252 12484 8256 12540
rect 8192 12480 8256 12484
rect 3012 11996 3076 12000
rect 3012 11940 3016 11996
rect 3016 11940 3072 11996
rect 3072 11940 3076 11996
rect 3012 11936 3076 11940
rect 3092 11996 3156 12000
rect 3092 11940 3096 11996
rect 3096 11940 3152 11996
rect 3152 11940 3156 11996
rect 3092 11936 3156 11940
rect 3172 11996 3236 12000
rect 3172 11940 3176 11996
rect 3176 11940 3232 11996
rect 3232 11940 3236 11996
rect 3172 11936 3236 11940
rect 3252 11996 3316 12000
rect 3252 11940 3256 11996
rect 3256 11940 3312 11996
rect 3312 11940 3316 11996
rect 3252 11936 3316 11940
rect 9444 11732 9508 11796
rect 1716 11596 1780 11660
rect 6316 11596 6380 11660
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 7952 11452 8016 11456
rect 7952 11396 7956 11452
rect 7956 11396 8012 11452
rect 8012 11396 8016 11452
rect 7952 11392 8016 11396
rect 8032 11452 8096 11456
rect 8032 11396 8036 11452
rect 8036 11396 8092 11452
rect 8092 11396 8096 11452
rect 8032 11392 8096 11396
rect 8112 11452 8176 11456
rect 8112 11396 8116 11452
rect 8116 11396 8172 11452
rect 8172 11396 8176 11452
rect 8112 11392 8176 11396
rect 8192 11452 8256 11456
rect 8192 11396 8196 11452
rect 8196 11396 8252 11452
rect 8252 11396 8256 11452
rect 8192 11392 8256 11396
rect 9260 11188 9324 11252
rect 3012 10908 3076 10912
rect 3012 10852 3016 10908
rect 3016 10852 3072 10908
rect 3072 10852 3076 10908
rect 3012 10848 3076 10852
rect 3092 10908 3156 10912
rect 3092 10852 3096 10908
rect 3096 10852 3152 10908
rect 3152 10852 3156 10908
rect 3092 10848 3156 10852
rect 3172 10908 3236 10912
rect 3172 10852 3176 10908
rect 3176 10852 3232 10908
rect 3232 10852 3236 10908
rect 3172 10848 3236 10852
rect 3252 10908 3316 10912
rect 3252 10852 3256 10908
rect 3256 10852 3312 10908
rect 3312 10852 3316 10908
rect 3252 10848 3316 10852
rect 6500 10644 6564 10708
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 7952 10364 8016 10368
rect 7952 10308 7956 10364
rect 7956 10308 8012 10364
rect 8012 10308 8016 10364
rect 7952 10304 8016 10308
rect 8032 10364 8096 10368
rect 8032 10308 8036 10364
rect 8036 10308 8092 10364
rect 8092 10308 8096 10364
rect 8032 10304 8096 10308
rect 8112 10364 8176 10368
rect 8112 10308 8116 10364
rect 8116 10308 8172 10364
rect 8172 10308 8176 10364
rect 8112 10304 8176 10308
rect 8192 10364 8256 10368
rect 8192 10308 8196 10364
rect 8196 10308 8252 10364
rect 8252 10308 8256 10364
rect 8192 10304 8256 10308
rect 3012 9820 3076 9824
rect 3012 9764 3016 9820
rect 3016 9764 3072 9820
rect 3072 9764 3076 9820
rect 3012 9760 3076 9764
rect 3092 9820 3156 9824
rect 3092 9764 3096 9820
rect 3096 9764 3152 9820
rect 3152 9764 3156 9820
rect 3092 9760 3156 9764
rect 3172 9820 3236 9824
rect 3172 9764 3176 9820
rect 3176 9764 3232 9820
rect 3232 9764 3236 9820
rect 3172 9760 3236 9764
rect 3252 9820 3316 9824
rect 3252 9764 3256 9820
rect 3256 9764 3312 9820
rect 3312 9764 3316 9820
rect 3252 9760 3316 9764
rect 8708 9420 8772 9484
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 7952 9276 8016 9280
rect 7952 9220 7956 9276
rect 7956 9220 8012 9276
rect 8012 9220 8016 9276
rect 7952 9216 8016 9220
rect 8032 9276 8096 9280
rect 8032 9220 8036 9276
rect 8036 9220 8092 9276
rect 8092 9220 8096 9276
rect 8032 9216 8096 9220
rect 8112 9276 8176 9280
rect 8112 9220 8116 9276
rect 8116 9220 8172 9276
rect 8172 9220 8176 9276
rect 8112 9216 8176 9220
rect 8192 9276 8256 9280
rect 8192 9220 8196 9276
rect 8196 9220 8252 9276
rect 8252 9220 8256 9276
rect 8192 9216 8256 9220
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9444 8468 9508 8532
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 3740 1260 3804 1324
rect 6684 1260 6748 1324
rect 3556 1124 3620 1188
rect 5396 988 5460 1052
rect 5212 36 5276 100
<< metal4 >>
rect 1944 41920 2264 45016
rect 1944 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2264 41920
rect 1531 41716 1597 41717
rect 1531 41652 1532 41716
rect 1596 41652 1597 41716
rect 1531 41651 1597 41652
rect 1534 16285 1594 41651
rect 1715 41444 1781 41445
rect 1715 41380 1716 41444
rect 1780 41380 1781 41444
rect 1715 41379 1781 41380
rect 1531 16284 1597 16285
rect 1531 16220 1532 16284
rect 1596 16220 1597 16284
rect 1531 16219 1597 16220
rect 1718 11661 1778 41379
rect 1944 40832 2264 41856
rect 1944 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2264 40832
rect 1944 39744 2264 40768
rect 1944 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2264 39744
rect 1944 38656 2264 39680
rect 1944 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2264 38656
rect 1944 37568 2264 38592
rect 1944 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2264 37568
rect 1944 36480 2264 37504
rect 1944 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2264 36480
rect 1944 35392 2264 36416
rect 1944 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2264 35392
rect 1944 34304 2264 35328
rect 1944 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2264 34304
rect 1944 33216 2264 34240
rect 1944 33152 1952 33216
rect 2016 33152 2032 33216
rect 2096 33152 2112 33216
rect 2176 33152 2192 33216
rect 2256 33152 2264 33216
rect 1944 32128 2264 33152
rect 1944 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2264 32128
rect 1944 31040 2264 32064
rect 1944 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2264 31040
rect 1944 29952 2264 30976
rect 1944 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2264 29952
rect 1944 28864 2264 29888
rect 1944 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2264 28864
rect 1944 27776 2264 28800
rect 1944 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2264 27776
rect 1944 26688 2264 27712
rect 1944 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2264 26688
rect 1944 25600 2264 26624
rect 1944 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2264 25600
rect 1944 24512 2264 25536
rect 1944 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2264 24512
rect 1944 23424 2264 24448
rect 1944 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2264 23424
rect 1944 22336 2264 23360
rect 1944 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2264 22336
rect 1944 21248 2264 22272
rect 1944 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2264 21248
rect 1944 20160 2264 21184
rect 1944 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2264 20160
rect 1944 19072 2264 20096
rect 1944 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2264 19072
rect 1944 17984 2264 19008
rect 1944 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2264 17984
rect 1944 16896 2264 17920
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 12544 2264 13568
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1715 11660 1781 11661
rect 1715 11596 1716 11660
rect 1780 11596 1781 11660
rect 1715 11595 1781 11596
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 42464 3324 45016
rect 3004 42400 3012 42464
rect 3076 42400 3092 42464
rect 3156 42400 3172 42464
rect 3236 42400 3252 42464
rect 3316 42400 3324 42464
rect 3004 41376 3324 42400
rect 7944 41920 8264 45016
rect 7944 41856 7952 41920
rect 8016 41856 8032 41920
rect 8096 41856 8112 41920
rect 8176 41856 8192 41920
rect 8256 41856 8264 41920
rect 5027 41444 5093 41445
rect 5027 41380 5028 41444
rect 5092 41380 5093 41444
rect 5027 41379 5093 41380
rect 3004 41312 3012 41376
rect 3076 41312 3092 41376
rect 3156 41312 3172 41376
rect 3236 41312 3252 41376
rect 3316 41312 3324 41376
rect 3004 40288 3324 41312
rect 3004 40224 3012 40288
rect 3076 40224 3092 40288
rect 3156 40224 3172 40288
rect 3236 40224 3252 40288
rect 3316 40224 3324 40288
rect 3004 39200 3324 40224
rect 3004 39136 3012 39200
rect 3076 39136 3092 39200
rect 3156 39136 3172 39200
rect 3236 39136 3252 39200
rect 3316 39136 3324 39200
rect 3004 38112 3324 39136
rect 3004 38048 3012 38112
rect 3076 38048 3092 38112
rect 3156 38048 3172 38112
rect 3236 38048 3252 38112
rect 3316 38048 3324 38112
rect 3004 37024 3324 38048
rect 3004 36960 3012 37024
rect 3076 36960 3092 37024
rect 3156 36960 3172 37024
rect 3236 36960 3252 37024
rect 3316 36960 3324 37024
rect 3004 35936 3324 36960
rect 3004 35872 3012 35936
rect 3076 35872 3092 35936
rect 3156 35872 3172 35936
rect 3236 35872 3252 35936
rect 3316 35872 3324 35936
rect 3004 34848 3324 35872
rect 3004 34784 3012 34848
rect 3076 34784 3092 34848
rect 3156 34784 3172 34848
rect 3236 34784 3252 34848
rect 3316 34784 3324 34848
rect 3004 33760 3324 34784
rect 3004 33696 3012 33760
rect 3076 33696 3092 33760
rect 3156 33696 3172 33760
rect 3236 33696 3252 33760
rect 3316 33696 3324 33760
rect 3004 32672 3324 33696
rect 4659 33556 4725 33557
rect 4659 33492 4660 33556
rect 4724 33492 4725 33556
rect 4659 33491 4725 33492
rect 3004 32608 3012 32672
rect 3076 32608 3092 32672
rect 3156 32608 3172 32672
rect 3236 32608 3252 32672
rect 3316 32608 3324 32672
rect 3004 31584 3324 32608
rect 3004 31520 3012 31584
rect 3076 31520 3092 31584
rect 3156 31520 3172 31584
rect 3236 31520 3252 31584
rect 3316 31520 3324 31584
rect 3004 30496 3324 31520
rect 3004 30432 3012 30496
rect 3076 30432 3092 30496
rect 3156 30432 3172 30496
rect 3236 30432 3252 30496
rect 3316 30432 3324 30496
rect 3004 29408 3324 30432
rect 3004 29344 3012 29408
rect 3076 29344 3092 29408
rect 3156 29344 3172 29408
rect 3236 29344 3252 29408
rect 3316 29344 3324 29408
rect 3004 28320 3324 29344
rect 3923 29068 3989 29069
rect 3923 29004 3924 29068
rect 3988 29004 3989 29068
rect 3923 29003 3989 29004
rect 3004 28256 3012 28320
rect 3076 28256 3092 28320
rect 3156 28256 3172 28320
rect 3236 28256 3252 28320
rect 3316 28256 3324 28320
rect 3004 27232 3324 28256
rect 3004 27168 3012 27232
rect 3076 27168 3092 27232
rect 3156 27168 3172 27232
rect 3236 27168 3252 27232
rect 3316 27168 3324 27232
rect 3004 26144 3324 27168
rect 3004 26080 3012 26144
rect 3076 26080 3092 26144
rect 3156 26080 3172 26144
rect 3236 26080 3252 26144
rect 3316 26080 3324 26144
rect 3004 25056 3324 26080
rect 3555 25260 3621 25261
rect 3555 25196 3556 25260
rect 3620 25196 3621 25260
rect 3555 25195 3621 25196
rect 3004 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3172 25056
rect 3236 24992 3252 25056
rect 3316 24992 3324 25056
rect 3004 23968 3324 24992
rect 3004 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3172 23968
rect 3236 23904 3252 23968
rect 3316 23904 3324 23968
rect 3004 22880 3324 23904
rect 3004 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3172 22880
rect 3236 22816 3252 22880
rect 3316 22816 3324 22880
rect 3004 21792 3324 22816
rect 3004 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3172 21792
rect 3236 21728 3252 21792
rect 3316 21728 3324 21792
rect 3004 20704 3324 21728
rect 3004 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3172 20704
rect 3236 20640 3252 20704
rect 3316 20640 3324 20704
rect 3004 19616 3324 20640
rect 3004 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3324 19616
rect 3004 18528 3324 19552
rect 3004 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3324 18528
rect 3004 17440 3324 18464
rect 3004 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3324 17440
rect 3004 16352 3324 17376
rect 3004 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3324 16352
rect 3004 15264 3324 16288
rect 3004 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3324 15264
rect 3004 14176 3324 15200
rect 3004 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3324 14176
rect 3004 13088 3324 14112
rect 3004 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3324 13088
rect 3004 12000 3324 13024
rect 3004 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3324 12000
rect 3004 10912 3324 11936
rect 3004 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3324 10912
rect 3004 9824 3324 10848
rect 3004 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3324 9824
rect 3004 8736 3324 9760
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 3558 1189 3618 25195
rect 3739 23492 3805 23493
rect 3739 23428 3740 23492
rect 3804 23428 3805 23492
rect 3739 23427 3805 23428
rect 3742 1325 3802 23427
rect 3926 19549 3986 29003
rect 3923 19548 3989 19549
rect 3923 19484 3924 19548
rect 3988 19484 3989 19548
rect 3923 19483 3989 19484
rect 4662 13837 4722 33491
rect 5030 16285 5090 41379
rect 7944 40832 8264 41856
rect 7944 40768 7952 40832
rect 8016 40768 8032 40832
rect 8096 40768 8112 40832
rect 8176 40768 8192 40832
rect 8256 40768 8264 40832
rect 7944 39744 8264 40768
rect 7944 39680 7952 39744
rect 8016 39680 8032 39744
rect 8096 39680 8112 39744
rect 8176 39680 8192 39744
rect 8256 39680 8264 39744
rect 7944 38656 8264 39680
rect 7944 38592 7952 38656
rect 8016 38592 8032 38656
rect 8096 38592 8112 38656
rect 8176 38592 8192 38656
rect 8256 38592 8264 38656
rect 7944 37568 8264 38592
rect 7944 37504 7952 37568
rect 8016 37504 8032 37568
rect 8096 37504 8112 37568
rect 8176 37504 8192 37568
rect 8256 37504 8264 37568
rect 7944 36480 8264 37504
rect 7944 36416 7952 36480
rect 8016 36416 8032 36480
rect 8096 36416 8112 36480
rect 8176 36416 8192 36480
rect 8256 36416 8264 36480
rect 7944 35392 8264 36416
rect 7944 35328 7952 35392
rect 8016 35328 8032 35392
rect 8096 35328 8112 35392
rect 8176 35328 8192 35392
rect 8256 35328 8264 35392
rect 7944 34304 8264 35328
rect 7944 34240 7952 34304
rect 8016 34240 8032 34304
rect 8096 34240 8112 34304
rect 8176 34240 8192 34304
rect 8256 34240 8264 34304
rect 7944 33216 8264 34240
rect 7944 33152 7952 33216
rect 8016 33152 8032 33216
rect 8096 33152 8112 33216
rect 8176 33152 8192 33216
rect 8256 33152 8264 33216
rect 7944 32128 8264 33152
rect 7944 32064 7952 32128
rect 8016 32064 8032 32128
rect 8096 32064 8112 32128
rect 8176 32064 8192 32128
rect 8256 32064 8264 32128
rect 7944 31040 8264 32064
rect 7944 30976 7952 31040
rect 8016 30976 8032 31040
rect 8096 30976 8112 31040
rect 8176 30976 8192 31040
rect 8256 30976 8264 31040
rect 7944 29952 8264 30976
rect 7944 29888 7952 29952
rect 8016 29888 8032 29952
rect 8096 29888 8112 29952
rect 8176 29888 8192 29952
rect 8256 29888 8264 29952
rect 7944 28864 8264 29888
rect 7944 28800 7952 28864
rect 8016 28800 8032 28864
rect 8096 28800 8112 28864
rect 8176 28800 8192 28864
rect 8256 28800 8264 28864
rect 7944 27776 8264 28800
rect 7944 27712 7952 27776
rect 8016 27712 8032 27776
rect 8096 27712 8112 27776
rect 8176 27712 8192 27776
rect 8256 27712 8264 27776
rect 7944 26688 8264 27712
rect 7944 26624 7952 26688
rect 8016 26624 8032 26688
rect 8096 26624 8112 26688
rect 8176 26624 8192 26688
rect 8256 26624 8264 26688
rect 7603 26348 7669 26349
rect 7603 26284 7604 26348
rect 7668 26284 7669 26348
rect 7603 26283 7669 26284
rect 7235 24852 7301 24853
rect 7235 24788 7236 24852
rect 7300 24788 7301 24852
rect 7235 24787 7301 24788
rect 5395 24036 5461 24037
rect 5395 23972 5396 24036
rect 5460 23972 5461 24036
rect 5395 23971 5461 23972
rect 5211 23492 5277 23493
rect 5211 23428 5212 23492
rect 5276 23428 5277 23492
rect 5211 23427 5277 23428
rect 5027 16284 5093 16285
rect 5027 16220 5028 16284
rect 5092 16220 5093 16284
rect 5027 16219 5093 16220
rect 4659 13836 4725 13837
rect 4659 13772 4660 13836
rect 4724 13772 4725 13836
rect 4659 13771 4725 13772
rect 3739 1324 3805 1325
rect 3739 1260 3740 1324
rect 3804 1260 3805 1324
rect 3739 1259 3805 1260
rect 3555 1188 3621 1189
rect 3555 1124 3556 1188
rect 3620 1124 3621 1188
rect 3555 1123 3621 1124
rect 5214 101 5274 23427
rect 5398 1053 5458 23971
rect 6499 23492 6565 23493
rect 6499 23428 6500 23492
rect 6564 23428 6565 23492
rect 6499 23427 6565 23428
rect 6131 20908 6197 20909
rect 6131 20844 6132 20908
rect 6196 20844 6197 20908
rect 6131 20843 6197 20844
rect 6134 13837 6194 20843
rect 6315 20772 6381 20773
rect 6315 20708 6316 20772
rect 6380 20708 6381 20772
rect 6315 20707 6381 20708
rect 6131 13836 6197 13837
rect 6131 13772 6132 13836
rect 6196 13772 6197 13836
rect 6131 13771 6197 13772
rect 6318 11661 6378 20707
rect 6315 11660 6381 11661
rect 6315 11596 6316 11660
rect 6380 11596 6381 11660
rect 6315 11595 6381 11596
rect 6502 10709 6562 23427
rect 7238 22133 7298 24787
rect 7419 22540 7485 22541
rect 7419 22476 7420 22540
rect 7484 22476 7485 22540
rect 7419 22475 7485 22476
rect 7235 22132 7301 22133
rect 7235 22068 7236 22132
rect 7300 22068 7301 22132
rect 7235 22067 7301 22068
rect 6683 21044 6749 21045
rect 6683 20980 6684 21044
rect 6748 20980 6749 21044
rect 6683 20979 6749 20980
rect 6499 10708 6565 10709
rect 6499 10644 6500 10708
rect 6564 10644 6565 10708
rect 6499 10643 6565 10644
rect 6686 1325 6746 20979
rect 7235 20364 7301 20365
rect 7235 20300 7236 20364
rect 7300 20300 7301 20364
rect 7235 20299 7301 20300
rect 7238 15469 7298 20299
rect 7422 17917 7482 22475
rect 7419 17916 7485 17917
rect 7419 17852 7420 17916
rect 7484 17852 7485 17916
rect 7419 17851 7485 17852
rect 7606 15469 7666 26283
rect 7944 25600 8264 26624
rect 7944 25536 7952 25600
rect 8016 25536 8032 25600
rect 8096 25536 8112 25600
rect 8176 25536 8192 25600
rect 8256 25536 8264 25600
rect 7944 24512 8264 25536
rect 7944 24448 7952 24512
rect 8016 24448 8032 24512
rect 8096 24448 8112 24512
rect 8176 24448 8192 24512
rect 8256 24448 8264 24512
rect 7944 23424 8264 24448
rect 7944 23360 7952 23424
rect 8016 23360 8032 23424
rect 8096 23360 8112 23424
rect 8176 23360 8192 23424
rect 8256 23360 8264 23424
rect 7944 22336 8264 23360
rect 9443 22812 9509 22813
rect 9443 22748 9444 22812
rect 9508 22810 9509 22812
rect 9508 22750 9690 22810
rect 9508 22748 9509 22750
rect 9443 22747 9509 22748
rect 9443 22540 9509 22541
rect 9443 22476 9444 22540
rect 9508 22476 9509 22540
rect 9443 22475 9509 22476
rect 7944 22272 7952 22336
rect 8016 22272 8032 22336
rect 8096 22272 8112 22336
rect 8176 22272 8192 22336
rect 8256 22272 8264 22336
rect 7944 21248 8264 22272
rect 8339 21452 8405 21453
rect 8339 21388 8340 21452
rect 8404 21388 8405 21452
rect 8339 21387 8405 21388
rect 7944 21184 7952 21248
rect 8016 21184 8032 21248
rect 8096 21184 8112 21248
rect 8176 21184 8192 21248
rect 8256 21184 8264 21248
rect 7944 20160 8264 21184
rect 7944 20096 7952 20160
rect 8016 20096 8032 20160
rect 8096 20096 8112 20160
rect 8176 20096 8192 20160
rect 8256 20096 8264 20160
rect 7944 19072 8264 20096
rect 7944 19008 7952 19072
rect 8016 19008 8032 19072
rect 8096 19008 8112 19072
rect 8176 19008 8192 19072
rect 8256 19008 8264 19072
rect 7944 17984 8264 19008
rect 7944 17920 7952 17984
rect 8016 17920 8032 17984
rect 8096 17920 8112 17984
rect 8176 17920 8192 17984
rect 8256 17920 8264 17984
rect 7944 16896 8264 17920
rect 8342 17645 8402 21387
rect 9259 20636 9325 20637
rect 9259 20572 9260 20636
rect 9324 20572 9325 20636
rect 9259 20571 9325 20572
rect 8707 20500 8773 20501
rect 8707 20436 8708 20500
rect 8772 20436 8773 20500
rect 8707 20435 8773 20436
rect 8339 17644 8405 17645
rect 8339 17580 8340 17644
rect 8404 17580 8405 17644
rect 8339 17579 8405 17580
rect 7944 16832 7952 16896
rect 8016 16832 8032 16896
rect 8096 16832 8112 16896
rect 8176 16832 8192 16896
rect 8256 16832 8264 16896
rect 7944 15808 8264 16832
rect 7944 15744 7952 15808
rect 8016 15744 8032 15808
rect 8096 15744 8112 15808
rect 8176 15744 8192 15808
rect 8256 15744 8264 15808
rect 7235 15468 7301 15469
rect 7235 15404 7236 15468
rect 7300 15404 7301 15468
rect 7235 15403 7301 15404
rect 7603 15468 7669 15469
rect 7603 15404 7604 15468
rect 7668 15404 7669 15468
rect 7603 15403 7669 15404
rect 7944 14720 8264 15744
rect 7944 14656 7952 14720
rect 8016 14656 8032 14720
rect 8096 14656 8112 14720
rect 8176 14656 8192 14720
rect 8256 14656 8264 14720
rect 7944 13632 8264 14656
rect 7944 13568 7952 13632
rect 8016 13568 8032 13632
rect 8096 13568 8112 13632
rect 8176 13568 8192 13632
rect 8256 13568 8264 13632
rect 7944 12544 8264 13568
rect 7944 12480 7952 12544
rect 8016 12480 8032 12544
rect 8096 12480 8112 12544
rect 8176 12480 8192 12544
rect 8256 12480 8264 12544
rect 7944 11456 8264 12480
rect 7944 11392 7952 11456
rect 8016 11392 8032 11456
rect 8096 11392 8112 11456
rect 8176 11392 8192 11456
rect 8256 11392 8264 11456
rect 7944 10368 8264 11392
rect 7944 10304 7952 10368
rect 8016 10304 8032 10368
rect 8096 10304 8112 10368
rect 8176 10304 8192 10368
rect 8256 10304 8264 10368
rect 7944 9280 8264 10304
rect 8710 9485 8770 20435
rect 9262 11253 9322 20571
rect 9446 11797 9506 22475
rect 9443 11796 9509 11797
rect 9443 11732 9444 11796
rect 9508 11732 9509 11796
rect 9443 11731 9509 11732
rect 9259 11252 9325 11253
rect 9259 11188 9260 11252
rect 9324 11188 9325 11252
rect 9259 11187 9325 11188
rect 8707 9484 8773 9485
rect 8707 9420 8708 9484
rect 8772 9420 8773 9484
rect 8707 9419 8773 9420
rect 7944 9216 7952 9280
rect 8016 9216 8032 9280
rect 8096 9216 8112 9280
rect 8176 9216 8192 9280
rect 8256 9216 8264 9280
rect 7944 8192 8264 9216
rect 9443 8532 9509 8533
rect 9443 8468 9444 8532
rect 9508 8530 9509 8532
rect 9630 8530 9690 22750
rect 9508 8470 9690 8530
rect 9508 8468 9509 8470
rect 9443 8467 9509 8468
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 6683 1324 6749 1325
rect 6683 1260 6684 1324
rect 6748 1260 6749 1324
rect 6683 1259 6749 1260
rect 5395 1052 5461 1053
rect 5395 988 5396 1052
rect 5460 988 5461 1052
rect 5395 987 5461 988
rect 5211 100 5277 101
rect 5211 36 5212 100
rect 5276 36 5277 100
rect 5211 35 5277 36
rect 7944 0 8264 2688
use sky130_fd_sc_hd__buf_1  _000_
timestamp -3599
transform 1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform -1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _004_
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _005_
timestamp -3599
transform 1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform -1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _009_
timestamp -3599
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _011_
timestamp -3599
transform -1 0 7728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _012_
timestamp -3599
transform 1 0 7820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _013_
timestamp -3599
transform -1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _014_
timestamp -3599
transform -1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _015_
timestamp -3599
transform 1 0 5612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 6716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _018_
timestamp -3599
transform 1 0 7084 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _019_
timestamp -3599
transform -1 0 7728 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _020_
timestamp -3599
transform -1 0 7728 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _021_
timestamp -3599
transform -1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _022_
timestamp -3599
transform -1 0 7728 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _023_
timestamp -3599
transform -1 0 7360 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _024_
timestamp -3599
transform -1 0 7544 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _025_
timestamp -3599
transform -1 0 7360 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _026_
timestamp -3599
transform -1 0 7268 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _027_
timestamp -3599
transform -1 0 7452 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _028_
timestamp -3599
transform -1 0 6992 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _029_
timestamp -3599
transform 1 0 5060 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 6440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_
timestamp -3599
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp -3599
transform -1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp -3599
transform -1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp -3599
transform -1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp -3599
transform -1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp -3599
transform -1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp -3599
transform -1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp -3599
transform -1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _039_
timestamp -3599
transform 1 0 6716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform -1 0 8188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _041_
timestamp -3599
transform 1 0 7820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp -3599
transform -1 0 7544 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform -1 0 7452 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp -3599
transform -1 0 7268 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform -1 0 7268 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform -1 0 7544 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform -1 0 7728 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform -1 0 7728 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform -1 0 1840 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 2852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform -1 0 2300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp -3599
transform -1 0 3036 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp -3599
transform -1 0 2852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp -3599
transform -1 0 2668 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp -3599
transform -1 0 2300 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp -3599
transform 1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp -3599
transform -1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp -3599
transform 1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp -3599
transform 1 0 1564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp -3599
transform 1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp -3599
transform 1 0 1564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp -3599
transform 1 0 1840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp -3599
transform -1 0 1932 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp -3599
transform -1 0 1840 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp -3599
transform -1 0 2300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp -3599
transform 1 0 2392 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp -3599
transform -1 0 2668 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp -3599
transform 1 0 2484 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp -3599
transform -1 0 2944 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp -3599
transform -1 0 3036 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp -3599
transform -1 0 7728 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp -3599
transform -1 0 2300 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp -3599
transform -1 0 7728 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp -3599
transform -1 0 7728 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform -1 0 7728 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp -3599
transform -1 0 7728 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform -1 0 7912 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp -3599
transform -1 0 7728 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp -3599
transform 1 0 7728 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _080_
timestamp -3599
transform -1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _081_
timestamp -3599
transform -1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _082_
timestamp -3599
transform -1 0 2024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _083_
timestamp -3599
transform 1 0 1932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _084_
timestamp -3599
transform 1 0 2392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _085_
timestamp -3599
transform -1 0 3680 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _086_
timestamp -3599
transform -1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp -3599
transform 1 0 3588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _088_
timestamp -3599
transform 1 0 4692 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform -1 0 4968 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _090_
timestamp -3599
transform 1 0 5336 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _091_
timestamp -3599
transform 1 0 4600 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _092_
timestamp -3599
transform 1 0 4508 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp -3599
transform -1 0 3588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _094_
timestamp -3599
transform 1 0 2944 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _095_
timestamp -3599
transform 1 0 4876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp -3599
transform 1 0 6992 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp -3599
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _098_
timestamp -3599
transform 1 0 6992 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _099_
timestamp -3599
transform 1 0 6716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp -3599
transform 1 0 1656 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 2760 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 2944 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform 1 0 4876 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 6992 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform 1 0 6992 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform 1 0 3588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 7636 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 7452 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 7268 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6
timestamp -3599
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp -3599
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12
timestamp -3599
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18
timestamp -3599
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21
timestamp -3599
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp -3599
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35
timestamp -3599
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp -3599
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp -3599
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47
timestamp -3599
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50
timestamp -3599
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60
timestamp -3599
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp -3599
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp -3599
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp -3599
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78
timestamp -3599
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6
timestamp -3599
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_9
timestamp -3599
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_12
timestamp -3599
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_15
timestamp -3599
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_18
timestamp -3599
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_21
timestamp -3599
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_24
timestamp -3599
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp -3599
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_30
timestamp -3599
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_33
timestamp -3599
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_36
timestamp -3599
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_39
timestamp -3599
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_42
timestamp -3599
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_45
timestamp -3599
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_48
timestamp -3599
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_60
timestamp -3599
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_63
timestamp -3599
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_66
timestamp -3599
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp -3599
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_72
timestamp -3599
transform 1 0 7728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_76
timestamp -3599
transform 1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_79
timestamp -3599
transform 1 0 8372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_6
timestamp -3599
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_9
timestamp -3599
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_12
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_18
timestamp -3599
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_21
timestamp -3599
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_24
timestamp -3599
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp -3599
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_35
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_38
timestamp -3599
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp -3599
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_44
timestamp -3599
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_47
timestamp -3599
transform 1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp -3599
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp -3599
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp -3599
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_59
timestamp -3599
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_62
timestamp -3599
transform 1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_65
timestamp -3599
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp -3599
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_71
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_6
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_9
timestamp -3599
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_12
timestamp -3599
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_18
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_21
timestamp -3599
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_24
timestamp -3599
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp -3599
transform 1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_30
timestamp -3599
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_33
timestamp -3599
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_36
timestamp -3599
transform 1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_39
timestamp -3599
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_42
timestamp -3599
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_45
timestamp -3599
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_48
timestamp -3599
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp -3599
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_60
timestamp -3599
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_63
timestamp -3599
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_66
timestamp -3599
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_70
timestamp -3599
transform 1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_73
timestamp -3599
transform 1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_76
timestamp -3599
transform 1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_79
timestamp -3599
transform 1 0 8372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_6
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp -3599
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_12
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_18
timestamp -3599
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_21
timestamp -3599
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_24
timestamp -3599
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp -3599
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_35
timestamp -3599
transform 1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp -3599
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_44
timestamp -3599
transform 1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_47
timestamp -3599
transform 1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_50
timestamp -3599
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_56
timestamp -3599
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_59
timestamp -3599
transform 1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_62
timestamp -3599
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp -3599
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_68
timestamp -3599
transform 1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_71
timestamp -3599
transform 1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_74
timestamp -3599
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_6
timestamp -3599
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_9
timestamp -3599
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp -3599
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_18
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_21
timestamp -3599
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp -3599
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_33
timestamp -3599
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_36
timestamp -3599
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_42
timestamp -3599
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_45
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_48
timestamp -3599
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_60
timestamp -3599
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_63
timestamp -3599
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_66
timestamp -3599
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_72
timestamp -3599
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp -3599
transform 1 0 8280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_6
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_9
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_12
timestamp -3599
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_15
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_18
timestamp -3599
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_21
timestamp -3599
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_24
timestamp -3599
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_38
timestamp -3599
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_44
timestamp -3599
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_47
timestamp -3599
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_50
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_54
timestamp -3599
transform 1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_57
timestamp -3599
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_60
timestamp -3599
transform 1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_63
timestamp -3599
transform 1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_66
timestamp -3599
transform 1 0 7176 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_69
timestamp -3599
transform 1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_72
timestamp -3599
transform 1 0 7728 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_75
timestamp -3599
transform 1 0 8004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_78
timestamp -3599
transform 1 0 8280 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_6
timestamp -3599
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_9
timestamp -3599
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_12
timestamp -3599
transform 1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_18
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_21
timestamp -3599
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_30
timestamp -3599
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_33
timestamp -3599
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_36
timestamp -3599
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_39
timestamp -3599
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_42
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_45
timestamp -3599
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_48
timestamp -3599
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp -3599
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_60
timestamp -3599
transform 1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_63
timestamp -3599
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp -3599
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_75
timestamp -3599
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp -3599
transform 1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_6
timestamp -3599
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_9
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_12
timestamp -3599
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp -3599
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_18
timestamp -3599
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_21
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp -3599
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_35
timestamp -3599
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp -3599
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp -3599
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_47
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_50
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp -3599
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_56
timestamp -3599
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_59
timestamp -3599
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_68
timestamp -3599
transform 1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_71
timestamp -3599
transform 1 0 7636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_75
timestamp -3599
transform 1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp -3599
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6
timestamp -3599
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_9
timestamp -3599
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_12
timestamp -3599
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp -3599
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_18
timestamp -3599
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_21
timestamp -3599
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_24
timestamp -3599
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp -3599
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_30
timestamp -3599
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_33
timestamp -3599
transform 1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_36
timestamp -3599
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_39
timestamp -3599
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_42
timestamp -3599
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_45
timestamp -3599
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_48
timestamp -3599
transform 1 0 5520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_51
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp -3599
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_60
timestamp -3599
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_63
timestamp -3599
transform 1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_66
timestamp -3599
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_72
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_75
timestamp -3599
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp -3599
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_6
timestamp -3599
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_9
timestamp -3599
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_12
timestamp -3599
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_18
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_24
timestamp -3599
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp -3599
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_35
timestamp -3599
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_38
timestamp -3599
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_44
timestamp -3599
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_47
timestamp -3599
transform 1 0 5428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_50
timestamp -3599
transform 1 0 5704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_53
timestamp -3599
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_56
timestamp -3599
transform 1 0 6256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_59
timestamp -3599
transform 1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_62
timestamp -3599
transform 1 0 6808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_67
timestamp -3599
transform 1 0 7268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_70
timestamp -3599
transform 1 0 7544 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_73
timestamp -3599
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_76
timestamp -3599
transform 1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_79
timestamp -3599
transform 1 0 8372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_6
timestamp -3599
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_9
timestamp -3599
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_12
timestamp -3599
transform 1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_15
timestamp -3599
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_18
timestamp -3599
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_21
timestamp -3599
transform 1 0 3036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_24
timestamp -3599
transform 1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_27
timestamp -3599
transform 1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_30
timestamp -3599
transform 1 0 3864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_33
timestamp -3599
transform 1 0 4140 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_36
timestamp -3599
transform 1 0 4416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_39
timestamp -3599
transform 1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_42
timestamp -3599
transform 1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_45
timestamp -3599
transform 1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_48
timestamp -3599
transform 1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_51
timestamp -3599
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp -3599
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_60
timestamp -3599
transform 1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_63
timestamp -3599
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_66
timestamp -3599
transform 1 0 7176 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_69
timestamp -3599
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_72
timestamp -3599
transform 1 0 7728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_75
timestamp -3599
transform 1 0 8004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp -3599
transform 1 0 8280 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp -3599
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_6
timestamp -3599
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_9
timestamp -3599
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_12
timestamp -3599
transform 1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_15
timestamp -3599
transform 1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_18
timestamp -3599
transform 1 0 2760 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_21
timestamp -3599
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_24
timestamp -3599
transform 1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp -3599
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp -3599
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp -3599
transform 1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_35
timestamp -3599
transform 1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_38
timestamp -3599
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_41
timestamp -3599
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_44
timestamp -3599
transform 1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_47
timestamp -3599
transform 1 0 5428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_50
timestamp -3599
transform 1 0 5704 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_53
timestamp -3599
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_56
timestamp -3599
transform 1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_59
timestamp -3599
transform 1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_62
timestamp -3599
transform 1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_68
timestamp -3599
transform 1 0 7360 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_71
timestamp -3599
transform 1 0 7636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_74
timestamp -3599
transform 1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_77
timestamp -3599
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp -3599
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_6
timestamp -3599
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_9
timestamp -3599
transform 1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_12
timestamp -3599
transform 1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_15
timestamp -3599
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_18
timestamp -3599
transform 1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_21
timestamp -3599
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_24
timestamp -3599
transform 1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_27
timestamp -3599
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_30
timestamp -3599
transform 1 0 3864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_33
timestamp -3599
transform 1 0 4140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_36
timestamp -3599
transform 1 0 4416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_39
timestamp -3599
transform 1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_42
timestamp -3599
transform 1 0 4968 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_45
timestamp -3599
transform 1 0 5244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_48
timestamp -3599
transform 1 0 5520 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_51
timestamp -3599
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp -3599
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp -3599
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_60
timestamp -3599
transform 1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_66
timestamp -3599
transform 1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_69
timestamp -3599
transform 1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_72
timestamp -3599
transform 1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_75
timestamp -3599
transform 1 0 8004 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_78
timestamp -3599
transform 1 0 8280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp -3599
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_6
timestamp -3599
transform 1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_9
timestamp -3599
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_12
timestamp -3599
transform 1 0 2208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_15
timestamp -3599
transform 1 0 2484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_18
timestamp -3599
transform 1 0 2760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_21
timestamp -3599
transform 1 0 3036 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_24
timestamp -3599
transform 1 0 3312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp -3599
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_29
timestamp -3599
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_32
timestamp -3599
transform 1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_35
timestamp -3599
transform 1 0 4324 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_38
timestamp -3599
transform 1 0 4600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_41
timestamp -3599
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_44
timestamp -3599
transform 1 0 5152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_47
timestamp -3599
transform 1 0 5428 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_50
timestamp -3599
transform 1 0 5704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_53
timestamp -3599
transform 1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_56
timestamp -3599
transform 1 0 6256 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_59
timestamp -3599
transform 1 0 6532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_62
timestamp -3599
transform 1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_65
timestamp -3599
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_68
timestamp -3599
transform 1 0 7360 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_71
timestamp -3599
transform 1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_74
timestamp -3599
transform 1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_77
timestamp -3599
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp -3599
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_6
timestamp -3599
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_9
timestamp -3599
transform 1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_12
timestamp -3599
transform 1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_15
timestamp -3599
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_18
timestamp -3599
transform 1 0 2760 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_21
timestamp -3599
transform 1 0 3036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_24
timestamp -3599
transform 1 0 3312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp -3599
transform 1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_30
timestamp -3599
transform 1 0 3864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_33
timestamp -3599
transform 1 0 4140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_36
timestamp -3599
transform 1 0 4416 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_39
timestamp -3599
transform 1 0 4692 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_42
timestamp -3599
transform 1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_45
timestamp -3599
transform 1 0 5244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_48
timestamp -3599
transform 1 0 5520 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_51
timestamp -3599
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp -3599
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp -3599
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp -3599
transform 1 0 6624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_64
timestamp -3599
transform 1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_67
timestamp -3599
transform 1 0 7268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_70
timestamp -3599
transform 1 0 7544 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_73
timestamp -3599
transform 1 0 7820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_76
timestamp -3599
transform 1 0 8096 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_79
timestamp -3599
transform 1 0 8372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp -3599
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp -3599
transform 1 0 1656 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_11
timestamp -3599
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_14
timestamp -3599
transform 1 0 2392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_17
timestamp -3599
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_20
timestamp -3599
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_23
timestamp -3599
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp -3599
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_29
timestamp -3599
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp -3599
transform 1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_35
timestamp -3599
transform 1 0 4324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_38
timestamp -3599
transform 1 0 4600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp -3599
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_44
timestamp -3599
transform 1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_47
timestamp -3599
transform 1 0 5428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_52
timestamp -3599
transform 1 0 5888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_55
timestamp -3599
transform 1 0 6164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_58
timestamp -3599
transform 1 0 6440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_61
timestamp -3599
transform 1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_64
timestamp -3599
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_67
timestamp -3599
transform 1 0 7268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_70
timestamp -3599
transform 1 0 7544 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_73
timestamp -3599
transform 1 0 7820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_76
timestamp -3599
transform 1 0 8096 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_79
timestamp -3599
transform 1 0 8372 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp -3599
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_6
timestamp -3599
transform 1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_9
timestamp -3599
transform 1 0 1932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_12
timestamp -3599
transform 1 0 2208 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_15
timestamp -3599
transform 1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_18
timestamp -3599
transform 1 0 2760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_21
timestamp -3599
transform 1 0 3036 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_24
timestamp -3599
transform 1 0 3312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_27
timestamp -3599
transform 1 0 3588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_30
timestamp -3599
transform 1 0 3864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_33
timestamp -3599
transform 1 0 4140 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_36
timestamp -3599
transform 1 0 4416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_39
timestamp -3599
transform 1 0 4692 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_42
timestamp -3599
transform 1 0 4968 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_45
timestamp -3599
transform 1 0 5244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_48
timestamp -3599
transform 1 0 5520 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_51
timestamp -3599
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp -3599
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_57
timestamp -3599
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_60
timestamp -3599
transform 1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_63
timestamp -3599
transform 1 0 6900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_66
timestamp -3599
transform 1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_69
timestamp -3599
transform 1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_72
timestamp -3599
transform 1 0 7728 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_76
timestamp -3599
transform 1 0 8096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_79
timestamp -3599
transform 1 0 8372 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp -3599
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_6
timestamp -3599
transform 1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_9
timestamp -3599
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_12
timestamp -3599
transform 1 0 2208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_15
timestamp -3599
transform 1 0 2484 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_18
timestamp -3599
transform 1 0 2760 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_21
timestamp -3599
transform 1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_24
timestamp -3599
transform 1 0 3312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -3599
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp -3599
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp -3599
transform 1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_35
timestamp -3599
transform 1 0 4324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_38
timestamp -3599
transform 1 0 4600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_41
timestamp -3599
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_44
timestamp -3599
transform 1 0 5152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_47
timestamp -3599
transform 1 0 5428 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_53
timestamp -3599
transform 1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_56
timestamp -3599
transform 1 0 6256 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_59
timestamp -3599
transform 1 0 6532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_62
timestamp -3599
transform 1 0 6808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_65
timestamp -3599
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_68
timestamp -3599
transform 1 0 7360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_72
timestamp -3599
transform 1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_75
timestamp -3599
transform 1 0 8004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_78
timestamp -3599
transform 1 0 8280 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp -3599
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_6
timestamp -3599
transform 1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_9
timestamp -3599
transform 1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_12
timestamp -3599
transform 1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_15
timestamp -3599
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_18
timestamp -3599
transform 1 0 2760 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_21
timestamp -3599
transform 1 0 3036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_24
timestamp -3599
transform 1 0 3312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_27
timestamp -3599
transform 1 0 3588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_30
timestamp -3599
transform 1 0 3864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_33
timestamp -3599
transform 1 0 4140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_36
timestamp -3599
transform 1 0 4416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_39
timestamp -3599
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_42
timestamp -3599
transform 1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_45
timestamp -3599
transform 1 0 5244 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_48
timestamp -3599
transform 1 0 5520 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_51
timestamp -3599
transform 1 0 5796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp -3599
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp -3599
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_60
timestamp -3599
transform 1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_63
timestamp -3599
transform 1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_66
timestamp -3599
transform 1 0 7176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_69
timestamp -3599
transform 1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_72
timestamp -3599
transform 1 0 7728 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_75
timestamp -3599
transform 1 0 8004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp -3599
transform 1 0 8280 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp -3599
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_9
timestamp -3599
transform 1 0 1932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_12
timestamp -3599
transform 1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_15
timestamp -3599
transform 1 0 2484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_18
timestamp -3599
transform 1 0 2760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_21
timestamp -3599
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_24
timestamp -3599
transform 1 0 3312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp -3599
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_29
timestamp -3599
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp -3599
transform 1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_35
timestamp -3599
transform 1 0 4324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_38
timestamp -3599
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_41
timestamp -3599
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_44
timestamp -3599
transform 1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_47
timestamp -3599
transform 1 0 5428 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_50
timestamp -3599
transform 1 0 5704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_53
timestamp -3599
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_56
timestamp -3599
transform 1 0 6256 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_59
timestamp -3599
transform 1 0 6532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_62
timestamp -3599
transform 1 0 6808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_65
timestamp -3599
transform 1 0 7084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_68
timestamp -3599
transform 1 0 7360 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp -3599
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_76
timestamp -3599
transform 1 0 8096 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_79
timestamp -3599
transform 1 0 8372 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp -3599
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_6
timestamp -3599
transform 1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_9
timestamp -3599
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_12
timestamp -3599
transform 1 0 2208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_15
timestamp -3599
transform 1 0 2484 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_18
timestamp -3599
transform 1 0 2760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_21
timestamp -3599
transform 1 0 3036 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_24
timestamp -3599
transform 1 0 3312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_27
timestamp -3599
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_30
timestamp -3599
transform 1 0 3864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_33
timestamp -3599
transform 1 0 4140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_36
timestamp -3599
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_39
timestamp -3599
transform 1 0 4692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_42
timestamp -3599
transform 1 0 4968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_45
timestamp -3599
transform 1 0 5244 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_48
timestamp -3599
transform 1 0 5520 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_51
timestamp -3599
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp -3599
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp -3599
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_60
timestamp -3599
transform 1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_63
timestamp -3599
transform 1 0 6900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_66
timestamp -3599
transform 1 0 7176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp -3599
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_72
timestamp -3599
transform 1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_75
timestamp -3599
transform 1 0 8004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_78
timestamp -3599
transform 1 0 8280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp -3599
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_6
timestamp -3599
transform 1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_12
timestamp -3599
transform 1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_15
timestamp -3599
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_18
timestamp -3599
transform 1 0 2760 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_21
timestamp -3599
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_24
timestamp -3599
transform 1 0 3312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp -3599
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_29
timestamp -3599
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp -3599
transform 1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_35
timestamp -3599
transform 1 0 4324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_38
timestamp -3599
transform 1 0 4600 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_41
timestamp -3599
transform 1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_44
timestamp -3599
transform 1 0 5152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_47
timestamp -3599
transform 1 0 5428 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_50
timestamp -3599
transform 1 0 5704 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_53
timestamp -3599
transform 1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_56
timestamp -3599
transform 1 0 6256 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp -3599
transform 1 0 6532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_64
timestamp -3599
transform 1 0 6992 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_67
timestamp -3599
transform 1 0 7268 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_70
timestamp -3599
transform 1 0 7544 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_73
timestamp -3599
transform 1 0 7820 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_77
timestamp -3599
transform 1 0 8188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp -3599
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_6
timestamp -3599
transform 1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_9
timestamp -3599
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_12
timestamp -3599
transform 1 0 2208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_15
timestamp -3599
transform 1 0 2484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_18
timestamp -3599
transform 1 0 2760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_21
timestamp -3599
transform 1 0 3036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_24
timestamp -3599
transform 1 0 3312 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_27
timestamp -3599
transform 1 0 3588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_30
timestamp -3599
transform 1 0 3864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_33
timestamp -3599
transform 1 0 4140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_36
timestamp -3599
transform 1 0 4416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_39
timestamp -3599
transform 1 0 4692 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_42
timestamp -3599
transform 1 0 4968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_45
timestamp -3599
transform 1 0 5244 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_48
timestamp -3599
transform 1 0 5520 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_51
timestamp -3599
transform 1 0 5796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp -3599
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_60
timestamp -3599
transform 1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_63
timestamp -3599
transform 1 0 6900 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_66
timestamp -3599
transform 1 0 7176 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_69
timestamp -3599
transform 1 0 7452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_72
timestamp -3599
transform 1 0 7728 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_75
timestamp -3599
transform 1 0 8004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp -3599
transform 1 0 8280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp -3599
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_6
timestamp -3599
transform 1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_9
timestamp -3599
transform 1 0 1932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_13
timestamp -3599
transform 1 0 2300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_16
timestamp -3599
transform 1 0 2576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_19
timestamp -3599
transform 1 0 2852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_22
timestamp -3599
transform 1 0 3128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp -3599
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_29
timestamp -3599
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp -3599
transform 1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_35
timestamp -3599
transform 1 0 4324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_38
timestamp -3599
transform 1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_41
timestamp -3599
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_44
timestamp -3599
transform 1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_47
timestamp -3599
transform 1 0 5428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_50
timestamp -3599
transform 1 0 5704 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_53
timestamp -3599
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_56
timestamp -3599
transform 1 0 6256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_59
timestamp -3599
transform 1 0 6532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_62
timestamp -3599
transform 1 0 6808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_65
timestamp -3599
transform 1 0 7084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_68
timestamp -3599
transform 1 0 7360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_71
timestamp -3599
transform 1 0 7636 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_74
timestamp -3599
transform 1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_77
timestamp -3599
transform 1 0 8188 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp -3599
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_6
timestamp -3599
transform 1 0 1656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_11
timestamp -3599
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_14
timestamp -3599
transform 1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_17
timestamp -3599
transform 1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_20
timestamp -3599
transform 1 0 2944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_23
timestamp -3599
transform 1 0 3220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_26
timestamp -3599
transform 1 0 3496 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_29
timestamp -3599
transform 1 0 3772 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_32
timestamp -3599
transform 1 0 4048 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_35
timestamp -3599
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_38
timestamp -3599
transform 1 0 4600 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_42
timestamp -3599
transform 1 0 4968 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_45
timestamp -3599
transform 1 0 5244 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_48
timestamp -3599
transform 1 0 5520 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_51
timestamp -3599
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp -3599
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_60
timestamp -3599
transform 1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_63
timestamp -3599
transform 1 0 6900 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_66
timestamp -3599
transform 1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_71
timestamp -3599
transform 1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_74
timestamp -3599
transform 1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_77
timestamp -3599
transform 1 0 8188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp -3599
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_6
timestamp -3599
transform 1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_9
timestamp -3599
transform 1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_12
timestamp -3599
transform 1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_15
timestamp -3599
transform 1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_18
timestamp -3599
transform 1 0 2760 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_21
timestamp -3599
transform 1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_24
timestamp -3599
transform 1 0 3312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp -3599
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp -3599
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_32
timestamp -3599
transform 1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_35
timestamp -3599
transform 1 0 4324 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_38
timestamp -3599
transform 1 0 4600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_41
timestamp -3599
transform 1 0 4876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_44
timestamp -3599
transform 1 0 5152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_47
timestamp -3599
transform 1 0 5428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_50
timestamp -3599
transform 1 0 5704 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_53
timestamp -3599
transform 1 0 5980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_56
timestamp -3599
transform 1 0 6256 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_59
timestamp -3599
transform 1 0 6532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_62
timestamp -3599
transform 1 0 6808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_65
timestamp -3599
transform 1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_68
timestamp -3599
transform 1 0 7360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_71
timestamp -3599
transform 1 0 7636 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_74
timestamp -3599
transform 1 0 7912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_77
timestamp -3599
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp -3599
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_6
timestamp -3599
transform 1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_9
timestamp -3599
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_12
timestamp -3599
transform 1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_15
timestamp -3599
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_18
timestamp -3599
transform 1 0 2760 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_21
timestamp -3599
transform 1 0 3036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_24
timestamp -3599
transform 1 0 3312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_27
timestamp -3599
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_30
timestamp -3599
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_33
timestamp -3599
transform 1 0 4140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_36
timestamp -3599
transform 1 0 4416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_39
timestamp -3599
transform 1 0 4692 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_42
timestamp -3599
transform 1 0 4968 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_45
timestamp -3599
transform 1 0 5244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_48
timestamp -3599
transform 1 0 5520 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_51
timestamp -3599
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp -3599
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp -3599
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_60
timestamp -3599
transform 1 0 6624 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_66
timestamp -3599
transform 1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_69
timestamp -3599
transform 1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_72
timestamp -3599
transform 1 0 7728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_75
timestamp -3599
transform 1 0 8004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_78
timestamp -3599
transform 1 0 8280 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp -3599
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_8
timestamp -3599
transform 1 0 1840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_11
timestamp -3599
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_14
timestamp -3599
transform 1 0 2392 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_17
timestamp -3599
transform 1 0 2668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_20
timestamp -3599
transform 1 0 2944 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_23
timestamp -3599
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp -3599
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp -3599
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp -3599
transform 1 0 4048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_35
timestamp -3599
transform 1 0 4324 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_38
timestamp -3599
transform 1 0 4600 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_41
timestamp -3599
transform 1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_44
timestamp -3599
transform 1 0 5152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_47
timestamp -3599
transform 1 0 5428 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_50
timestamp -3599
transform 1 0 5704 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_53
timestamp -3599
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_56
timestamp -3599
transform 1 0 6256 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_59
timestamp -3599
transform 1 0 6532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_63
timestamp -3599
transform 1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_66
timestamp -3599
transform 1 0 7176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_69
timestamp -3599
transform 1 0 7452 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_72
timestamp -3599
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_75
timestamp -3599
transform 1 0 8004 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_78
timestamp -3599
transform 1 0 8280 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp -3599
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_6
timestamp -3599
transform 1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_9
timestamp -3599
transform 1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_12
timestamp -3599
transform 1 0 2208 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_15
timestamp -3599
transform 1 0 2484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_18
timestamp -3599
transform 1 0 2760 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_21
timestamp -3599
transform 1 0 3036 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_24
timestamp -3599
transform 1 0 3312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_27
timestamp -3599
transform 1 0 3588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_30
timestamp -3599
transform 1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_33
timestamp -3599
transform 1 0 4140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp -3599
transform 1 0 4416 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_41
timestamp -3599
transform 1 0 4876 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_44
timestamp -3599
transform 1 0 5152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_47
timestamp -3599
transform 1 0 5428 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_50
timestamp -3599
transform 1 0 5704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp -3599
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp -3599
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_60
timestamp -3599
transform 1 0 6624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_63
timestamp -3599
transform 1 0 6900 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp -3599
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_72
timestamp -3599
transform 1 0 7728 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_75
timestamp -3599
transform 1 0 8004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp -3599
transform 1 0 8280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp -3599
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_6
timestamp -3599
transform 1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_9
timestamp -3599
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_12
timestamp -3599
transform 1 0 2208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_15
timestamp -3599
transform 1 0 2484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_18
timestamp -3599
transform 1 0 2760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_21
timestamp -3599
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_24
timestamp -3599
transform 1 0 3312 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp -3599
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp -3599
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_32
timestamp -3599
transform 1 0 4048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_35
timestamp -3599
transform 1 0 4324 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_38
timestamp -3599
transform 1 0 4600 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_41
timestamp -3599
transform 1 0 4876 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_44
timestamp -3599
transform 1 0 5152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_47
timestamp -3599
transform 1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_50
timestamp -3599
transform 1 0 5704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_53
timestamp -3599
transform 1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_56
timestamp -3599
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_59
timestamp -3599
transform 1 0 6532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_62
timestamp -3599
transform 1 0 6808 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_68
timestamp -3599
transform 1 0 7360 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp -3599
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_9
timestamp -3599
transform 1 0 1932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_12
timestamp -3599
transform 1 0 2208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_15
timestamp -3599
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_18
timestamp -3599
transform 1 0 2760 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_21
timestamp -3599
transform 1 0 3036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_30
timestamp -3599
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_33
timestamp -3599
transform 1 0 4140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_36
timestamp -3599
transform 1 0 4416 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_39
timestamp -3599
transform 1 0 4692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_42
timestamp -3599
transform 1 0 4968 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_45
timestamp -3599
transform 1 0 5244 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_48
timestamp -3599
transform 1 0 5520 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_51
timestamp -3599
transform 1 0 5796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp -3599
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp -3599
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_61
timestamp -3599
transform 1 0 6716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_64
timestamp -3599
transform 1 0 6992 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_67
timestamp -3599
transform 1 0 7268 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp -3599
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_6
timestamp -3599
transform 1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_9
timestamp -3599
transform 1 0 1932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp -3599
transform 1 0 2208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_17
timestamp -3599
transform 1 0 2668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_20
timestamp -3599
transform 1 0 2944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_23
timestamp -3599
transform 1 0 3220 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp -3599
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_29
timestamp -3599
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_32
timestamp -3599
transform 1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_35
timestamp -3599
transform 1 0 4324 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_38
timestamp -3599
transform 1 0 4600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_42
timestamp -3599
transform 1 0 4968 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_45
timestamp -3599
transform 1 0 5244 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_48
timestamp -3599
transform 1 0 5520 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_51
timestamp -3599
transform 1 0 5796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_54
timestamp -3599
transform 1 0 6072 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_57
timestamp -3599
transform 1 0 6348 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_60
timestamp -3599
transform 1 0 6624 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_63
timestamp -3599
transform 1 0 6900 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_66
timestamp -3599
transform 1 0 7176 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_69
timestamp -3599
transform 1 0 7452 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp -3599
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_6
timestamp -3599
transform 1 0 1656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_9
timestamp -3599
transform 1 0 1932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_12
timestamp -3599
transform 1 0 2208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_15
timestamp -3599
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_18
timestamp -3599
transform 1 0 2760 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_21
timestamp -3599
transform 1 0 3036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_24
timestamp -3599
transform 1 0 3312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_27
timestamp -3599
transform 1 0 3588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_30
timestamp -3599
transform 1 0 3864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_33
timestamp -3599
transform 1 0 4140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_36
timestamp -3599
transform 1 0 4416 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_39
timestamp -3599
transform 1 0 4692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_42
timestamp -3599
transform 1 0 4968 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_49
timestamp -3599
transform 1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_52
timestamp -3599
transform 1 0 5888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp -3599
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_57
timestamp -3599
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_60
timestamp -3599
transform 1 0 6624 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_63
timestamp -3599
transform 1 0 6900 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_66
timestamp -3599
transform 1 0 7176 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_69
timestamp -3599
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp -3599
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_6
timestamp -3599
transform 1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_9
timestamp -3599
transform 1 0 1932 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_12
timestamp -3599
transform 1 0 2208 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_15
timestamp -3599
transform 1 0 2484 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_18
timestamp -3599
transform 1 0 2760 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_21
timestamp -3599
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_24
timestamp -3599
transform 1 0 3312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp -3599
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_29
timestamp -3599
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_32
timestamp -3599
transform 1 0 4048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_35
timestamp -3599
transform 1 0 4324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_38
timestamp -3599
transform 1 0 4600 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_41
timestamp -3599
transform 1 0 4876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_44
timestamp -3599
transform 1 0 5152 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_47
timestamp -3599
transform 1 0 5428 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_50
timestamp -3599
transform 1 0 5704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_53
timestamp -3599
transform 1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_56
timestamp -3599
transform 1 0 6256 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_59
timestamp -3599
transform 1 0 6532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_64
timestamp -3599
transform 1 0 6992 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_67
timestamp -3599
transform 1 0 7268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_70
timestamp -3599
transform 1 0 7544 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp -3599
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_8
timestamp -3599
transform 1 0 1840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_11
timestamp -3599
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_14
timestamp -3599
transform 1 0 2392 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_17
timestamp -3599
transform 1 0 2668 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_20
timestamp -3599
transform 1 0 2944 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_23
timestamp -3599
transform 1 0 3220 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_26
timestamp -3599
transform 1 0 3496 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_29
timestamp -3599
transform 1 0 3772 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_32
timestamp -3599
transform 1 0 4048 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_35
timestamp -3599
transform 1 0 4324 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_38
timestamp -3599
transform 1 0 4600 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_41
timestamp -3599
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_44
timestamp -3599
transform 1 0 5152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_47
timestamp -3599
transform 1 0 5428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_50
timestamp -3599
transform 1 0 5704 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp -3599
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_57
timestamp -3599
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_60
timestamp -3599
transform 1 0 6624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_63
timestamp -3599
transform 1 0 6900 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_66
timestamp -3599
transform 1 0 7176 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_69
timestamp -3599
transform 1 0 7452 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp -3599
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_6
timestamp -3599
transform 1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_9
timestamp -3599
transform 1 0 1932 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_12
timestamp -3599
transform 1 0 2208 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_15
timestamp -3599
transform 1 0 2484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_18
timestamp -3599
transform 1 0 2760 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_21
timestamp -3599
transform 1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_24
timestamp -3599
transform 1 0 3312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp -3599
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_29
timestamp -3599
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_32
timestamp -3599
transform 1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_35
timestamp -3599
transform 1 0 4324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_40
timestamp -3599
transform 1 0 4784 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_43
timestamp -3599
transform 1 0 5060 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_46
timestamp -3599
transform 1 0 5336 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_49
timestamp -3599
transform 1 0 5612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_52
timestamp -3599
transform 1 0 5888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_55
timestamp -3599
transform 1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_58
timestamp -3599
transform 1 0 6440 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_66
timestamp -3599
transform 1 0 7176 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_70
timestamp -3599
transform 1 0 7544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp -3599
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_6
timestamp -3599
transform 1 0 1656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_11
timestamp -3599
transform 1 0 2116 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_14
timestamp -3599
transform 1 0 2392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_17
timestamp -3599
transform 1 0 2668 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_20
timestamp -3599
transform 1 0 2944 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_23
timestamp -3599
transform 1 0 3220 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_26
timestamp -3599
transform 1 0 3496 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_30
timestamp -3599
transform 1 0 3864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_33
timestamp -3599
transform 1 0 4140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_36
timestamp -3599
transform 1 0 4416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_39
timestamp -3599
transform 1 0 4692 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_42
timestamp -3599
transform 1 0 4968 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_45
timestamp -3599
transform 1 0 5244 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_48
timestamp -3599
transform 1 0 5520 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_51
timestamp -3599
transform 1 0 5796 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp -3599
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp -3599
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_60
timestamp -3599
transform 1 0 6624 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_63
timestamp -3599
transform 1 0 6900 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_67
timestamp -3599
transform 1 0 7268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_71
timestamp -3599
transform 1 0 7636 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp -3599
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_6
timestamp -3599
transform 1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_9
timestamp -3599
transform 1 0 1932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_12
timestamp -3599
transform 1 0 2208 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_15
timestamp -3599
transform 1 0 2484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_18
timestamp -3599
transform 1 0 2760 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_21
timestamp -3599
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_24
timestamp -3599
transform 1 0 3312 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp -3599
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp -3599
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_32
timestamp -3599
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_35
timestamp -3599
transform 1 0 4324 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_38
timestamp -3599
transform 1 0 4600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_41
timestamp -3599
transform 1 0 4876 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_44
timestamp -3599
transform 1 0 5152 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_47
timestamp -3599
transform 1 0 5428 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_50
timestamp -3599
transform 1 0 5704 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_53
timestamp -3599
transform 1 0 5980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_56
timestamp -3599
transform 1 0 6256 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_59
timestamp -3599
transform 1 0 6532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_62
timestamp -3599
transform 1 0 6808 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_65
timestamp -3599
transform 1 0 7084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_68
timestamp -3599
transform 1 0 7360 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp -3599
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_6
timestamp -3599
transform 1 0 1656 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_10
timestamp -3599
transform 1 0 2024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_13
timestamp -3599
transform 1 0 2300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_16
timestamp -3599
transform 1 0 2576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_19
timestamp -3599
transform 1 0 2852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_22
timestamp -3599
transform 1 0 3128 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_25
timestamp -3599
transform 1 0 3404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_28
timestamp -3599
transform 1 0 3680 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_31
timestamp -3599
transform 1 0 3956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_34
timestamp -3599
transform 1 0 4232 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_37
timestamp -3599
transform 1 0 4508 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_40
timestamp -3599
transform 1 0 4784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_43
timestamp -3599
transform 1 0 5060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_46
timestamp -3599
transform 1 0 5336 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_49
timestamp -3599
transform 1 0 5612 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_52
timestamp -3599
transform 1 0 5888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp -3599
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp -3599
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_60
timestamp -3599
transform 1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_63
timestamp -3599
transform 1 0 6900 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_66
timestamp -3599
transform 1 0 7176 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_69
timestamp -3599
transform 1 0 7452 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp -3599
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_6
timestamp -3599
transform 1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_9
timestamp -3599
transform 1 0 1932 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_12
timestamp -3599
transform 1 0 2208 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_15
timestamp -3599
transform 1 0 2484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_18
timestamp -3599
transform 1 0 2760 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_21
timestamp -3599
transform 1 0 3036 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_24
timestamp -3599
transform 1 0 3312 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_29
timestamp -3599
transform 1 0 3772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_32
timestamp -3599
transform 1 0 4048 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_35
timestamp -3599
transform 1 0 4324 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_38
timestamp -3599
transform 1 0 4600 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_44
timestamp -3599
transform 1 0 5152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_47
timestamp -3599
transform 1 0 5428 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_50
timestamp -3599
transform 1 0 5704 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_53
timestamp -3599
transform 1 0 5980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_56
timestamp -3599
transform 1 0 6256 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_59
timestamp -3599
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_62
timestamp -3599
transform 1 0 6808 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_66
timestamp -3599
transform 1 0 7176 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp -3599
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_6
timestamp -3599
transform 1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_9
timestamp -3599
transform 1 0 1932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_12
timestamp -3599
transform 1 0 2208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_15
timestamp -3599
transform 1 0 2484 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_18
timestamp -3599
transform 1 0 2760 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_21
timestamp -3599
transform 1 0 3036 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_24
timestamp -3599
transform 1 0 3312 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_27
timestamp -3599
transform 1 0 3588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_30
timestamp -3599
transform 1 0 3864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_33
timestamp -3599
transform 1 0 4140 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_36
timestamp -3599
transform 1 0 4416 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_39
timestamp -3599
transform 1 0 4692 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_42
timestamp -3599
transform 1 0 4968 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_45
timestamp -3599
transform 1 0 5244 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_48
timestamp -3599
transform 1 0 5520 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_51
timestamp -3599
transform 1 0 5796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp -3599
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_57
timestamp -3599
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_60
timestamp -3599
transform 1 0 6624 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_63
timestamp -3599
transform 1 0 6900 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_70
timestamp -3599
transform 1 0 7544 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_3
timestamp -3599
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_10
timestamp -3599
transform 1 0 2024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_13
timestamp -3599
transform 1 0 2300 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_16
timestamp -3599
transform 1 0 2576 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_19
timestamp -3599
transform 1 0 2852 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_22
timestamp -3599
transform 1 0 3128 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp -3599
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_29
timestamp -3599
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_32
timestamp -3599
transform 1 0 4048 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_35
timestamp -3599
transform 1 0 4324 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_38
timestamp -3599
transform 1 0 4600 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_41
timestamp -3599
transform 1 0 4876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_44
timestamp -3599
transform 1 0 5152 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_47
timestamp -3599
transform 1 0 5428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_50
timestamp -3599
transform 1 0 5704 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_53
timestamp -3599
transform 1 0 5980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_56
timestamp -3599
transform 1 0 6256 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_59
timestamp -3599
transform 1 0 6532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_62
timestamp -3599
transform 1 0 6808 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_65
timestamp -3599
transform 1 0 7084 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_69
timestamp -3599
transform 1 0 7452 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_3
timestamp -3599
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_6
timestamp -3599
transform 1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_12
timestamp -3599
transform 1 0 2208 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_15
timestamp -3599
transform 1 0 2484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_18
timestamp -3599
transform 1 0 2760 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_23
timestamp -3599
transform 1 0 3220 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_26
timestamp -3599
transform 1 0 3496 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_29
timestamp -3599
transform 1 0 3772 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_32
timestamp -3599
transform 1 0 4048 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_35
timestamp -3599
transform 1 0 4324 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_38
timestamp -3599
transform 1 0 4600 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_41
timestamp -3599
transform 1 0 4876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_44
timestamp -3599
transform 1 0 5152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_47
timestamp -3599
transform 1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_50
timestamp -3599
transform 1 0 5704 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp -3599
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_57
timestamp -3599
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_60
timestamp -3599
transform 1 0 6624 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_63
timestamp -3599
transform 1 0 6900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_67
timestamp -3599
transform 1 0 7268 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_70
timestamp -3599
transform 1 0 7544 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_3
timestamp -3599
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_6
timestamp -3599
transform 1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_9
timestamp -3599
transform 1 0 1932 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_12
timestamp -3599
transform 1 0 2208 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_15
timestamp -3599
transform 1 0 2484 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_18
timestamp -3599
transform 1 0 2760 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_21
timestamp -3599
transform 1 0 3036 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_24
timestamp -3599
transform 1 0 3312 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp -3599
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_29
timestamp -3599
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_32
timestamp -3599
transform 1 0 4048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_35
timestamp -3599
transform 1 0 4324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_38
timestamp -3599
transform 1 0 4600 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_41
timestamp -3599
transform 1 0 4876 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_44
timestamp -3599
transform 1 0 5152 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_47
timestamp -3599
transform 1 0 5428 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_50
timestamp -3599
transform 1 0 5704 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_53
timestamp -3599
transform 1 0 5980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_56
timestamp -3599
transform 1 0 6256 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_59
timestamp -3599
transform 1 0 6532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_62
timestamp -3599
transform 1 0 6808 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_69
timestamp -3599
transform 1 0 7452 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_3
timestamp -3599
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_6
timestamp -3599
transform 1 0 1656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_9
timestamp -3599
transform 1 0 1932 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_12
timestamp -3599
transform 1 0 2208 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_15
timestamp -3599
transform 1 0 2484 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_18
timestamp -3599
transform 1 0 2760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_21
timestamp -3599
transform 1 0 3036 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_24
timestamp -3599
transform 1 0 3312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_27
timestamp -3599
transform 1 0 3588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_30
timestamp -3599
transform 1 0 3864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_33
timestamp -3599
transform 1 0 4140 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_36
timestamp -3599
transform 1 0 4416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_39
timestamp -3599
transform 1 0 4692 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_42
timestamp -3599
transform 1 0 4968 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_45
timestamp -3599
transform 1 0 5244 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_48
timestamp -3599
transform 1 0 5520 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_51
timestamp -3599
transform 1 0 5796 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp -3599
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_57
timestamp -3599
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_60
timestamp -3599
transform 1 0 6624 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_63
timestamp -3599
transform 1 0 6900 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_66
timestamp -3599
transform 1 0 7176 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_70
timestamp -3599
transform 1 0 7544 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_3
timestamp -3599
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_6
timestamp -3599
transform 1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_9
timestamp -3599
transform 1 0 1932 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_12
timestamp -3599
transform 1 0 2208 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_17
timestamp -3599
transform 1 0 2668 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_20
timestamp -3599
transform 1 0 2944 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_23
timestamp -3599
transform 1 0 3220 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp -3599
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_29
timestamp -3599
transform 1 0 3772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_32
timestamp -3599
transform 1 0 4048 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_35
timestamp -3599
transform 1 0 4324 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_38
timestamp -3599
transform 1 0 4600 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_41
timestamp -3599
transform 1 0 4876 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_44
timestamp -3599
transform 1 0 5152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_47
timestamp -3599
transform 1 0 5428 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_50
timestamp -3599
transform 1 0 5704 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp -3599
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_56
timestamp -3599
transform 1 0 6256 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_59
timestamp -3599
transform 1 0 6532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_62
timestamp -3599
transform 1 0 6808 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_65
timestamp -3599
transform 1 0 7084 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_68
timestamp -3599
transform 1 0 7360 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_3
timestamp -3599
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_6
timestamp -3599
transform 1 0 1656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_9
timestamp -3599
transform 1 0 1932 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_12
timestamp -3599
transform 1 0 2208 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_15
timestamp -3599
transform 1 0 2484 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_18
timestamp -3599
transform 1 0 2760 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_21
timestamp -3599
transform 1 0 3036 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_24
timestamp -3599
transform 1 0 3312 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_27
timestamp -3599
transform 1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_30
timestamp -3599
transform 1 0 3864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_33
timestamp -3599
transform 1 0 4140 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_36
timestamp -3599
transform 1 0 4416 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_39
timestamp -3599
transform 1 0 4692 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_42
timestamp -3599
transform 1 0 4968 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_45
timestamp -3599
transform 1 0 5244 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_48
timestamp -3599
transform 1 0 5520 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_51
timestamp -3599
transform 1 0 5796 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp -3599
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_57
timestamp -3599
transform 1 0 6348 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_60
timestamp -3599
transform 1 0 6624 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_63
timestamp -3599
transform 1 0 6900 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_66
timestamp -3599
transform 1 0 7176 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_3
timestamp -3599
transform 1 0 1380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_6
timestamp -3599
transform 1 0 1656 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_9
timestamp -3599
transform 1 0 1932 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_12
timestamp -3599
transform 1 0 2208 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_15
timestamp -3599
transform 1 0 2484 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_18
timestamp -3599
transform 1 0 2760 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_21
timestamp -3599
transform 1 0 3036 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_24
timestamp -3599
transform 1 0 3312 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp -3599
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_29
timestamp -3599
transform 1 0 3772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_32
timestamp -3599
transform 1 0 4048 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_35
timestamp -3599
transform 1 0 4324 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_38
timestamp -3599
transform 1 0 4600 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_41
timestamp -3599
transform 1 0 4876 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_44
timestamp -3599
transform 1 0 5152 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_47
timestamp -3599
transform 1 0 5428 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_50
timestamp -3599
transform 1 0 5704 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_53
timestamp -3599
transform 1 0 5980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_56
timestamp -3599
transform 1 0 6256 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_59
timestamp -3599
transform 1 0 6532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_62
timestamp -3599
transform 1 0 6808 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_65
timestamp -3599
transform 1 0 7084 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_68
timestamp -3599
transform 1 0 7360 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_3
timestamp -3599
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_6
timestamp -3599
transform 1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_9
timestamp -3599
transform 1 0 1932 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_12
timestamp -3599
transform 1 0 2208 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_18
timestamp -3599
transform 1 0 2760 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_21
timestamp -3599
transform 1 0 3036 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_24
timestamp -3599
transform 1 0 3312 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_27
timestamp -3599
transform 1 0 3588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_30
timestamp -3599
transform 1 0 3864 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_33
timestamp -3599
transform 1 0 4140 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_36
timestamp -3599
transform 1 0 4416 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_39
timestamp -3599
transform 1 0 4692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_42
timestamp -3599
transform 1 0 4968 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_45
timestamp -3599
transform 1 0 5244 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_48
timestamp -3599
transform 1 0 5520 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_51
timestamp -3599
transform 1 0 5796 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp -3599
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_57
timestamp -3599
transform 1 0 6348 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_60
timestamp -3599
transform 1 0 6624 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_63
timestamp -3599
transform 1 0 6900 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_68
timestamp -3599
transform 1 0 7360 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_71
timestamp -3599
transform 1 0 7636 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_3
timestamp -3599
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_6
timestamp -3599
transform 1 0 1656 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_9
timestamp -3599
transform 1 0 1932 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_12
timestamp -3599
transform 1 0 2208 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_15
timestamp -3599
transform 1 0 2484 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_18
timestamp -3599
transform 1 0 2760 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_21
timestamp -3599
transform 1 0 3036 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_24
timestamp -3599
transform 1 0 3312 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp -3599
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_29
timestamp -3599
transform 1 0 3772 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_32
timestamp -3599
transform 1 0 4048 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_35
timestamp -3599
transform 1 0 4324 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_38
timestamp -3599
transform 1 0 4600 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_41
timestamp -3599
transform 1 0 4876 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_44
timestamp -3599
transform 1 0 5152 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_47
timestamp -3599
transform 1 0 5428 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_50
timestamp -3599
transform 1 0 5704 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_53
timestamp -3599
transform 1 0 5980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_56
timestamp -3599
transform 1 0 6256 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_59
timestamp -3599
transform 1 0 6532 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_62
timestamp -3599
transform 1 0 6808 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_65
timestamp -3599
transform 1 0 7084 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_70
timestamp -3599
transform 1 0 7544 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp -3599
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_8
timestamp -3599
transform 1 0 1840 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_11
timestamp -3599
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_14
timestamp -3599
transform 1 0 2392 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_19
timestamp -3599
transform 1 0 2852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_22
timestamp -3599
transform 1 0 3128 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_25
timestamp -3599
transform 1 0 3404 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_28
timestamp -3599
transform 1 0 3680 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_31
timestamp -3599
transform 1 0 3956 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_34
timestamp -3599
transform 1 0 4232 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_37
timestamp -3599
transform 1 0 4508 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_40
timestamp -3599
transform 1 0 4784 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_43
timestamp -3599
transform 1 0 5060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_46
timestamp -3599
transform 1 0 5336 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_49
timestamp -3599
transform 1 0 5612 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_52
timestamp -3599
transform 1 0 5888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp -3599
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_57
timestamp -3599
transform 1 0 6348 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_60
timestamp -3599
transform 1 0 6624 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_63
timestamp -3599
transform 1 0 6900 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_68
timestamp -3599
transform 1 0 7360 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_71
timestamp -3599
transform 1 0 7636 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_3
timestamp -3599
transform 1 0 1380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_6
timestamp -3599
transform 1 0 1656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_9
timestamp -3599
transform 1 0 1932 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_12
timestamp -3599
transform 1 0 2208 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_15
timestamp -3599
transform 1 0 2484 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_18
timestamp -3599
transform 1 0 2760 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_21
timestamp -3599
transform 1 0 3036 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_24
timestamp -3599
transform 1 0 3312 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp -3599
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_29
timestamp -3599
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_32
timestamp -3599
transform 1 0 4048 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_35
timestamp -3599
transform 1 0 4324 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_38
timestamp -3599
transform 1 0 4600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_41
timestamp -3599
transform 1 0 4876 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_44
timestamp -3599
transform 1 0 5152 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_47
timestamp -3599
transform 1 0 5428 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_50
timestamp -3599
transform 1 0 5704 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_53
timestamp -3599
transform 1 0 5980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_56
timestamp -3599
transform 1 0 6256 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_59
timestamp -3599
transform 1 0 6532 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_62
timestamp -3599
transform 1 0 6808 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_67
timestamp -3599
transform 1 0 7268 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_70
timestamp -3599
transform 1 0 7544 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_3
timestamp -3599
transform 1 0 1380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_6
timestamp -3599
transform 1 0 1656 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_9
timestamp -3599
transform 1 0 1932 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_13
timestamp -3599
transform 1 0 2300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_16
timestamp -3599
transform 1 0 2576 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_20
timestamp -3599
transform 1 0 2944 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_23
timestamp -3599
transform 1 0 3220 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_26
timestamp -3599
transform 1 0 3496 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_29
timestamp -3599
transform 1 0 3772 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_32
timestamp -3599
transform 1 0 4048 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_35
timestamp -3599
transform 1 0 4324 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_38
timestamp -3599
transform 1 0 4600 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_41
timestamp -3599
transform 1 0 4876 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_44
timestamp -3599
transform 1 0 5152 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_47
timestamp -3599
transform 1 0 5428 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_50
timestamp -3599
transform 1 0 5704 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp -3599
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_57
timestamp -3599
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_60
timestamp -3599
transform 1 0 6624 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_63
timestamp -3599
transform 1 0 6900 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_66
timestamp -3599
transform 1 0 7176 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_69
timestamp -3599
transform 1 0 7452 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp -3599
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_6
timestamp -3599
transform 1 0 1656 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_9
timestamp -3599
transform 1 0 1932 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_12
timestamp -3599
transform 1 0 2208 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_15
timestamp -3599
transform 1 0 2484 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_21
timestamp -3599
transform 1 0 3036 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_24
timestamp -3599
transform 1 0 3312 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp -3599
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_29
timestamp -3599
transform 1 0 3772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_32
timestamp -3599
transform 1 0 4048 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_35
timestamp -3599
transform 1 0 4324 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_38
timestamp -3599
transform 1 0 4600 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_41
timestamp -3599
transform 1 0 4876 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_44
timestamp -3599
transform 1 0 5152 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_47
timestamp -3599
transform 1 0 5428 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_50
timestamp -3599
transform 1 0 5704 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_53
timestamp -3599
transform 1 0 5980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_56
timestamp -3599
transform 1 0 6256 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_59
timestamp -3599
transform 1 0 6532 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_62
timestamp -3599
transform 1 0 6808 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_65
timestamp -3599
transform 1 0 7084 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_69
timestamp -3599
transform 1 0 7452 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_3
timestamp -3599
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_6
timestamp -3599
transform 1 0 1656 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_9
timestamp -3599
transform 1 0 1932 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_12
timestamp -3599
transform 1 0 2208 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_15
timestamp -3599
transform 1 0 2484 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_19
timestamp -3599
transform 1 0 2852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_22
timestamp -3599
transform 1 0 3128 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_25
timestamp -3599
transform 1 0 3404 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_28
timestamp -3599
transform 1 0 3680 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_31
timestamp -3599
transform 1 0 3956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_34
timestamp -3599
transform 1 0 4232 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_37
timestamp -3599
transform 1 0 4508 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_40
timestamp -3599
transform 1 0 4784 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_43
timestamp -3599
transform 1 0 5060 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_46
timestamp -3599
transform 1 0 5336 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_49
timestamp -3599
transform 1 0 5612 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_52
timestamp -3599
transform 1 0 5888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp -3599
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_57
timestamp -3599
transform 1 0 6348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_60
timestamp -3599
transform 1 0 6624 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_63
timestamp -3599
transform 1 0 6900 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_66
timestamp -3599
transform 1 0 7176 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_69
timestamp -3599
transform 1 0 7452 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_3
timestamp -3599
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_6
timestamp -3599
transform 1 0 1656 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_9
timestamp -3599
transform 1 0 1932 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_12
timestamp -3599
transform 1 0 2208 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_17
timestamp -3599
transform 1 0 2668 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_20
timestamp -3599
transform 1 0 2944 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_23
timestamp -3599
transform 1 0 3220 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp -3599
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_29
timestamp -3599
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_32
timestamp -3599
transform 1 0 4048 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_35
timestamp -3599
transform 1 0 4324 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_38
timestamp -3599
transform 1 0 4600 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_41
timestamp -3599
transform 1 0 4876 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_44
timestamp -3599
transform 1 0 5152 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_47
timestamp -3599
transform 1 0 5428 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_50
timestamp -3599
transform 1 0 5704 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_53
timestamp -3599
transform 1 0 5980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_56
timestamp -3599
transform 1 0 6256 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_59
timestamp -3599
transform 1 0 6532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_62
timestamp -3599
transform 1 0 6808 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_65
timestamp -3599
transform 1 0 7084 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_68
timestamp -3599
transform 1 0 7360 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_3
timestamp -3599
transform 1 0 1380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_9
timestamp -3599
transform 1 0 1932 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_12
timestamp -3599
transform 1 0 2208 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_15
timestamp -3599
transform 1 0 2484 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_18
timestamp -3599
transform 1 0 2760 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_21
timestamp -3599
transform 1 0 3036 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_24
timestamp -3599
transform 1 0 3312 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_27
timestamp -3599
transform 1 0 3588 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_30
timestamp -3599
transform 1 0 3864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_33
timestamp -3599
transform 1 0 4140 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_36
timestamp -3599
transform 1 0 4416 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_39
timestamp -3599
transform 1 0 4692 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_42
timestamp -3599
transform 1 0 4968 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_45
timestamp -3599
transform 1 0 5244 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_48
timestamp -3599
transform 1 0 5520 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_51
timestamp -3599
transform 1 0 5796 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp -3599
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_57
timestamp -3599
transform 1 0 6348 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_60
timestamp -3599
transform 1 0 6624 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_63
timestamp -3599
transform 1 0 6900 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_66
timestamp -3599
transform 1 0 7176 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_69
timestamp -3599
transform 1 0 7452 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_3
timestamp -3599
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_6
timestamp -3599
transform 1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_9
timestamp -3599
transform 1 0 1932 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_13
timestamp -3599
transform 1 0 2300 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_16
timestamp -3599
transform 1 0 2576 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_19
timestamp -3599
transform 1 0 2852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_22
timestamp -3599
transform 1 0 3128 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_25
timestamp -3599
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_29
timestamp -3599
transform 1 0 3772 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_32
timestamp -3599
transform 1 0 4048 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_35
timestamp -3599
transform 1 0 4324 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_38
timestamp -3599
transform 1 0 4600 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_41
timestamp -3599
transform 1 0 4876 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_44
timestamp -3599
transform 1 0 5152 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_47
timestamp -3599
transform 1 0 5428 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_50
timestamp -3599
transform 1 0 5704 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_53
timestamp -3599
transform 1 0 5980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_56
timestamp -3599
transform 1 0 6256 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_59
timestamp -3599
transform 1 0 6532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_62
timestamp -3599
transform 1 0 6808 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_65
timestamp -3599
transform 1 0 7084 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_68
timestamp -3599
transform 1 0 7360 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_71
timestamp -3599
transform 1 0 7636 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_3
timestamp -3599
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_6
timestamp -3599
transform 1 0 1656 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_9
timestamp -3599
transform 1 0 1932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_12
timestamp -3599
transform 1 0 2208 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_15
timestamp -3599
transform 1 0 2484 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_18
timestamp -3599
transform 1 0 2760 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_21
timestamp -3599
transform 1 0 3036 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_24
timestamp -3599
transform 1 0 3312 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_27
timestamp -3599
transform 1 0 3588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_30
timestamp -3599
transform 1 0 3864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_33
timestamp -3599
transform 1 0 4140 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_36
timestamp -3599
transform 1 0 4416 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_39
timestamp -3599
transform 1 0 4692 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_42
timestamp -3599
transform 1 0 4968 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_45
timestamp -3599
transform 1 0 5244 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_48
timestamp -3599
transform 1 0 5520 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_51
timestamp -3599
transform 1 0 5796 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp -3599
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_57
timestamp -3599
transform 1 0 6348 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_60
timestamp -3599
transform 1 0 6624 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_63
timestamp -3599
transform 1 0 6900 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_66
timestamp -3599
transform 1 0 7176 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_69
timestamp -3599
transform 1 0 7452 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp -3599
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_8
timestamp -3599
transform 1 0 1840 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_11
timestamp -3599
transform 1 0 2116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_14
timestamp -3599
transform 1 0 2392 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_17
timestamp -3599
transform 1 0 2668 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_20
timestamp -3599
transform 1 0 2944 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_23
timestamp -3599
transform 1 0 3220 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp -3599
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_29
timestamp -3599
transform 1 0 3772 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_32
timestamp -3599
transform 1 0 4048 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_35
timestamp -3599
transform 1 0 4324 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_38
timestamp -3599
transform 1 0 4600 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_41
timestamp -3599
transform 1 0 4876 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_44
timestamp -3599
transform 1 0 5152 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_47
timestamp -3599
transform 1 0 5428 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_50
timestamp -3599
transform 1 0 5704 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_53
timestamp -3599
transform 1 0 5980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_56
timestamp -3599
transform 1 0 6256 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_59
timestamp -3599
transform 1 0 6532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_62
timestamp -3599
transform 1 0 6808 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_65
timestamp -3599
transform 1 0 7084 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_68
timestamp -3599
transform 1 0 7360 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_3
timestamp -3599
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_6
timestamp -3599
transform 1 0 1656 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_9
timestamp -3599
transform 1 0 1932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_12
timestamp -3599
transform 1 0 2208 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_15
timestamp -3599
transform 1 0 2484 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_18
timestamp -3599
transform 1 0 2760 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_21
timestamp -3599
transform 1 0 3036 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_24
timestamp -3599
transform 1 0 3312 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_27
timestamp -3599
transform 1 0 3588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_30
timestamp -3599
transform 1 0 3864 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_33
timestamp -3599
transform 1 0 4140 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_36
timestamp -3599
transform 1 0 4416 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_39
timestamp -3599
transform 1 0 4692 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_42
timestamp -3599
transform 1 0 4968 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_45
timestamp -3599
transform 1 0 5244 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_48
timestamp -3599
transform 1 0 5520 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_51
timestamp -3599
transform 1 0 5796 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp -3599
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_57
timestamp -3599
transform 1 0 6348 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_60
timestamp -3599
transform 1 0 6624 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_63
timestamp -3599
transform 1 0 6900 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_66
timestamp -3599
transform 1 0 7176 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_69
timestamp -3599
transform 1 0 7452 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_3
timestamp -3599
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_6
timestamp -3599
transform 1 0 1656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_9
timestamp -3599
transform 1 0 1932 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_13
timestamp -3599
transform 1 0 2300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_16
timestamp -3599
transform 1 0 2576 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_19
timestamp -3599
transform 1 0 2852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_22
timestamp -3599
transform 1 0 3128 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_25
timestamp -3599
transform 1 0 3404 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_29
timestamp -3599
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_32
timestamp -3599
transform 1 0 4048 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_35
timestamp -3599
transform 1 0 4324 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_38
timestamp -3599
transform 1 0 4600 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_41
timestamp -3599
transform 1 0 4876 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_44
timestamp -3599
transform 1 0 5152 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_47
timestamp -3599
transform 1 0 5428 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_50
timestamp -3599
transform 1 0 5704 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_53
timestamp -3599
transform 1 0 5980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_56
timestamp -3599
transform 1 0 6256 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_59
timestamp -3599
transform 1 0 6532 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_62
timestamp -3599
transform 1 0 6808 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_65
timestamp -3599
transform 1 0 7084 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_68
timestamp -3599
transform 1 0 7360 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_71
timestamp -3599
transform 1 0 7636 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_3
timestamp -3599
transform 1 0 1380 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_6
timestamp -3599
transform 1 0 1656 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_9
timestamp -3599
transform 1 0 1932 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_12
timestamp -3599
transform 1 0 2208 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_17
timestamp -3599
transform 1 0 2668 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_20
timestamp -3599
transform 1 0 2944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_23
timestamp -3599
transform 1 0 3220 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_26
timestamp -3599
transform 1 0 3496 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_29
timestamp -3599
transform 1 0 3772 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_32
timestamp -3599
transform 1 0 4048 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_35
timestamp -3599
transform 1 0 4324 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_38
timestamp -3599
transform 1 0 4600 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_41
timestamp -3599
transform 1 0 4876 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_44
timestamp -3599
transform 1 0 5152 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_47
timestamp -3599
transform 1 0 5428 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_50
timestamp -3599
transform 1 0 5704 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp -3599
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_57
timestamp -3599
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_60
timestamp -3599
transform 1 0 6624 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_63
timestamp -3599
transform 1 0 6900 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_66
timestamp -3599
transform 1 0 7176 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_69
timestamp -3599
transform 1 0 7452 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_3
timestamp -3599
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_6
timestamp -3599
transform 1 0 1656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_9
timestamp -3599
transform 1 0 1932 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_12
timestamp -3599
transform 1 0 2208 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_15
timestamp -3599
transform 1 0 2484 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_18
timestamp -3599
transform 1 0 2760 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_21
timestamp -3599
transform 1 0 3036 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_24
timestamp -3599
transform 1 0 3312 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp -3599
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_29
timestamp -3599
transform 1 0 3772 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_32
timestamp -3599
transform 1 0 4048 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_35
timestamp -3599
transform 1 0 4324 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_38
timestamp -3599
transform 1 0 4600 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_41
timestamp -3599
transform 1 0 4876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_44
timestamp -3599
transform 1 0 5152 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_47
timestamp -3599
transform 1 0 5428 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_50
timestamp -3599
transform 1 0 5704 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp -3599
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_56
timestamp -3599
transform 1 0 6256 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_59
timestamp -3599
transform 1 0 6532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_62
timestamp -3599
transform 1 0 6808 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_65
timestamp -3599
transform 1 0 7084 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_68
timestamp -3599
transform 1 0 7360 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_3
timestamp -3599
transform 1 0 1380 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_6
timestamp -3599
transform 1 0 1656 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_9
timestamp -3599
transform 1 0 1932 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_12
timestamp -3599
transform 1 0 2208 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_15
timestamp -3599
transform 1 0 2484 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_18
timestamp -3599
transform 1 0 2760 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_21
timestamp -3599
transform 1 0 3036 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_24
timestamp -3599
transform 1 0 3312 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_27
timestamp -3599
transform 1 0 3588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_30
timestamp -3599
transform 1 0 3864 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_33
timestamp -3599
transform 1 0 4140 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_36
timestamp -3599
transform 1 0 4416 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_39
timestamp -3599
transform 1 0 4692 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_42
timestamp -3599
transform 1 0 4968 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_45
timestamp -3599
transform 1 0 5244 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_48
timestamp -3599
transform 1 0 5520 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_51
timestamp -3599
transform 1 0 5796 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp -3599
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_57
timestamp -3599
transform 1 0 6348 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_60
timestamp -3599
transform 1 0 6624 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_63
timestamp -3599
transform 1 0 6900 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_66
timestamp -3599
transform 1 0 7176 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_3
timestamp -3599
transform 1 0 1380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_6
timestamp -3599
transform 1 0 1656 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_9
timestamp -3599
transform 1 0 1932 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_12
timestamp -3599
transform 1 0 2208 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_15
timestamp -3599
transform 1 0 2484 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_20
timestamp -3599
transform 1 0 2944 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_23
timestamp -3599
transform 1 0 3220 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp -3599
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_29
timestamp -3599
transform 1 0 3772 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_32
timestamp -3599
transform 1 0 4048 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_35
timestamp -3599
transform 1 0 4324 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_38
timestamp -3599
transform 1 0 4600 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_41
timestamp -3599
transform 1 0 4876 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_44
timestamp -3599
transform 1 0 5152 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_47
timestamp -3599
transform 1 0 5428 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_50
timestamp -3599
transform 1 0 5704 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_53
timestamp -3599
transform 1 0 5980 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_56
timestamp -3599
transform 1 0 6256 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_59
timestamp -3599
transform 1 0 6532 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_62
timestamp -3599
transform 1 0 6808 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_65
timestamp -3599
transform 1 0 7084 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_68
timestamp -3599
transform 1 0 7360 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_3
timestamp -3599
transform 1 0 1380 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_6
timestamp -3599
transform 1 0 1656 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_9
timestamp -3599
transform 1 0 1932 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_12
timestamp -3599
transform 1 0 2208 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_15
timestamp -3599
transform 1 0 2484 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_18
timestamp -3599
transform 1 0 2760 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_21
timestamp -3599
transform 1 0 3036 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_24
timestamp -3599
transform 1 0 3312 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_27
timestamp -3599
transform 1 0 3588 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_30
timestamp -3599
transform 1 0 3864 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_33
timestamp -3599
transform 1 0 4140 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_36
timestamp -3599
transform 1 0 4416 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_39
timestamp -3599
transform 1 0 4692 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_42
timestamp -3599
transform 1 0 4968 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_45
timestamp -3599
transform 1 0 5244 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_48
timestamp -3599
transform 1 0 5520 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_51
timestamp -3599
transform 1 0 5796 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp -3599
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_57
timestamp -3599
transform 1 0 6348 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_60
timestamp -3599
transform 1 0 6624 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_63
timestamp -3599
transform 1 0 6900 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_66
timestamp -3599
transform 1 0 7176 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_69
timestamp -3599
transform 1 0 7452 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_3
timestamp -3599
transform 1 0 1380 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_6
timestamp -3599
transform 1 0 1656 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_9
timestamp -3599
transform 1 0 1932 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_12
timestamp -3599
transform 1 0 2208 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_15
timestamp -3599
transform 1 0 2484 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_21
timestamp -3599
transform 1 0 3036 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_24
timestamp -3599
transform 1 0 3312 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp -3599
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_29
timestamp -3599
transform 1 0 3772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_32
timestamp -3599
transform 1 0 4048 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_35
timestamp -3599
transform 1 0 4324 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_38
timestamp -3599
transform 1 0 4600 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_41
timestamp -3599
transform 1 0 4876 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_44
timestamp -3599
transform 1 0 5152 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_47
timestamp -3599
transform 1 0 5428 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_50
timestamp -3599
transform 1 0 5704 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_53
timestamp -3599
transform 1 0 5980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_56
timestamp -3599
transform 1 0 6256 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_59
timestamp -3599
transform 1 0 6532 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_62
timestamp -3599
transform 1 0 6808 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_65
timestamp -3599
transform 1 0 7084 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_68
timestamp -3599
transform 1 0 7360 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_3
timestamp -3599
transform 1 0 1380 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_6
timestamp -3599
transform 1 0 1656 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_9
timestamp -3599
transform 1 0 1932 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_12
timestamp -3599
transform 1 0 2208 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_15
timestamp -3599
transform 1 0 2484 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_18
timestamp -3599
transform 1 0 2760 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_21
timestamp -3599
transform 1 0 3036 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_24
timestamp -3599
transform 1 0 3312 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_27
timestamp -3599
transform 1 0 3588 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_30
timestamp -3599
transform 1 0 3864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_33
timestamp -3599
transform 1 0 4140 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_36
timestamp -3599
transform 1 0 4416 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_39
timestamp -3599
transform 1 0 4692 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_42
timestamp -3599
transform 1 0 4968 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_45
timestamp -3599
transform 1 0 5244 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_48
timestamp -3599
transform 1 0 5520 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_51
timestamp -3599
transform 1 0 5796 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_54
timestamp -3599
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_57
timestamp -3599
transform 1 0 6348 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_60
timestamp -3599
transform 1 0 6624 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_63
timestamp -3599
transform 1 0 6900 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_66
timestamp -3599
transform 1 0 7176 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_69_69
timestamp -3599
transform 1 0 7452 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_3
timestamp -3599
transform 1 0 1380 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_6
timestamp -3599
transform 1 0 1656 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_9
timestamp -3599
transform 1 0 1932 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_13
timestamp -3599
transform 1 0 2300 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_16
timestamp -3599
transform 1 0 2576 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_19
timestamp -3599
transform 1 0 2852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_22
timestamp -3599
transform 1 0 3128 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_25
timestamp -3599
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_29
timestamp -3599
transform 1 0 3772 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_32
timestamp -3599
transform 1 0 4048 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_35
timestamp -3599
transform 1 0 4324 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_38
timestamp -3599
transform 1 0 4600 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_41
timestamp -3599
transform 1 0 4876 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_44
timestamp -3599
transform 1 0 5152 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_47
timestamp -3599
transform 1 0 5428 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_50
timestamp -3599
transform 1 0 5704 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_53
timestamp -3599
transform 1 0 5980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_56
timestamp -3599
transform 1 0 6256 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_59
timestamp -3599
transform 1 0 6532 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_62
timestamp -3599
transform 1 0 6808 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_65
timestamp -3599
transform 1 0 7084 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_68
timestamp -3599
transform 1 0 7360 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_74
timestamp -3599
transform 1 0 7912 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_77
timestamp -3599
transform 1 0 8188 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_3
timestamp -3599
transform 1 0 1380 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_6
timestamp -3599
transform 1 0 1656 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_9
timestamp -3599
transform 1 0 1932 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_12
timestamp -3599
transform 1 0 2208 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_15
timestamp -3599
transform 1 0 2484 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_18
timestamp -3599
transform 1 0 2760 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_21
timestamp -3599
transform 1 0 3036 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_24
timestamp -3599
transform 1 0 3312 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_27
timestamp -3599
transform 1 0 3588 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_30
timestamp -3599
transform 1 0 3864 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_33
timestamp -3599
transform 1 0 4140 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_36
timestamp -3599
transform 1 0 4416 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_39
timestamp -3599
transform 1 0 4692 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_42
timestamp -3599
transform 1 0 4968 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_45
timestamp -3599
transform 1 0 5244 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_48
timestamp -3599
transform 1 0 5520 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_51
timestamp -3599
transform 1 0 5796 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp -3599
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_57
timestamp -3599
transform 1 0 6348 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_60
timestamp -3599
transform 1 0 6624 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_63
timestamp -3599
transform 1 0 6900 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_66
timestamp -3599
transform 1 0 7176 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_69
timestamp -3599
transform 1 0 7452 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_71_75
timestamp -3599
transform 1 0 8004 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_10
timestamp -3599
transform 1 0 2024 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_13
timestamp -3599
transform 1 0 2300 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_16
timestamp -3599
transform 1 0 2576 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_19
timestamp -3599
transform 1 0 2852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_22
timestamp -3599
transform 1 0 3128 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_25
timestamp -3599
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_29
timestamp -3599
transform 1 0 3772 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_32
timestamp -3599
transform 1 0 4048 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_35
timestamp -3599
transform 1 0 4324 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_38
timestamp -3599
transform 1 0 4600 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_41
timestamp -3599
transform 1 0 4876 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_44
timestamp -3599
transform 1 0 5152 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_47
timestamp -3599
transform 1 0 5428 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_50
timestamp -3599
transform 1 0 5704 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_53
timestamp -3599
transform 1 0 5980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_56
timestamp -3599
transform 1 0 6256 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_59
timestamp -3599
transform 1 0 6532 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_62
timestamp -3599
transform 1 0 6808 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_65
timestamp -3599
transform 1 0 7084 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_68
timestamp -3599
transform 1 0 7360 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_11
timestamp -3599
transform 1 0 2116 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_29
timestamp -3599
transform 1 0 3772 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_73_36
timestamp -3599
transform 1 0 4416 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_41
timestamp -3599
transform 1 0 4876 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_46
timestamp -3599
transform 1 0 5336 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_51
timestamp -3599
transform 1 0 5796 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_61
timestamp -3599
transform 1 0 6716 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_66
timestamp -3599
transform 1 0 7176 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_71
timestamp -3599
transform 1 0 7636 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 7728 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 8096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform -1 0 8096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 8096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 7728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 8096 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 7728 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 8096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 7728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 8096 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 7728 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 8096 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 7728 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 8096 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 7728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 8096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 7728 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 8096 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 7728 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 8096 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 8096 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 8096 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 7728 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 7728 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 8096 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 7728 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 8096 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 7728 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 8096 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 7728 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 8096 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 7728 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform 1 0 7728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform 1 0 8096 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform 1 0 7728 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform 1 0 8096 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform 1 0 7728 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 8096 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 7728 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 8096 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 7728 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform 1 0 8096 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform 1 0 7728 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 8096 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 7728 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 8096 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform -1 0 8096 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform 1 0 8096 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform 1 0 8096 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform 1 0 7728 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform 1 0 8096 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 7728 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 8096 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 7728 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 8096 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 7728 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 8096 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 7728 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 7728 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 8096 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 7728 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 8096 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 7728 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 8096 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 7728 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 8096 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 7728 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 8096 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 7728 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 8096 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 8096 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 7728 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 7728 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 8096 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 7728 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 8096 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 7728 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 8096 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 7728 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform -1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform -1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 5888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 6348 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 6808 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 7268 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 7728 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 8096 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform 1 0 8096 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 7728 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform 1 0 8096 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 2208 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 2576 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 3312 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 3680 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform 1 0 4048 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 4876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform 1 0 4968 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output101
timestamp -3599
transform -1 0 2024 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_74
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_75
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_76
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 8740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_77
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_78
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 8740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_79
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_80
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 8740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_81
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_82
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 8740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_83
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 8740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_84
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 8740 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_85
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 8740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_86
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 8740 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_87
timestamp -3599
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3599
transform -1 0 8740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_88
timestamp -3599
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -3599
transform -1 0 8740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_89
timestamp -3599
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -3599
transform -1 0 8740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_90
timestamp -3599
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -3599
transform -1 0 8740 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_91
timestamp -3599
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -3599
transform -1 0 8740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_92
timestamp -3599
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -3599
transform -1 0 8740 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_93
timestamp -3599
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -3599
transform -1 0 8740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_94
timestamp -3599
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -3599
transform -1 0 8740 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_95
timestamp -3599
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -3599
transform -1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_96
timestamp -3599
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -3599
transform -1 0 8740 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_97
timestamp -3599
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -3599
transform -1 0 8740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_98
timestamp -3599
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -3599
transform -1 0 8740 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_99
timestamp -3599
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -3599
transform -1 0 8740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_100
timestamp -3599
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -3599
transform -1 0 8740 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_101
timestamp -3599
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -3599
transform -1 0 8740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_102
timestamp -3599
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -3599
transform -1 0 8740 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_103
timestamp -3599
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -3599
transform -1 0 8740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_104
timestamp -3599
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -3599
transform -1 0 8740 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_105
timestamp -3599
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -3599
transform -1 0 8740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_106
timestamp -3599
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -3599
transform -1 0 8740 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_107
timestamp -3599
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -3599
transform -1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_108
timestamp -3599
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp -3599
transform -1 0 8740 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_109
timestamp -3599
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp -3599
transform -1 0 8740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_110
timestamp -3599
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp -3599
transform -1 0 8740 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_111
timestamp -3599
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp -3599
transform -1 0 8740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_112
timestamp -3599
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp -3599
transform -1 0 8740 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_113
timestamp -3599
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp -3599
transform -1 0 8740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_114
timestamp -3599
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp -3599
transform -1 0 8740 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_115
timestamp -3599
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp -3599
transform -1 0 8740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_116
timestamp -3599
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp -3599
transform -1 0 8740 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_117
timestamp -3599
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp -3599
transform -1 0 8740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_118
timestamp -3599
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp -3599
transform -1 0 8740 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_119
timestamp -3599
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp -3599
transform -1 0 8740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_120
timestamp -3599
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp -3599
transform -1 0 8740 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_121
timestamp -3599
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp -3599
transform -1 0 8740 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_122
timestamp -3599
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp -3599
transform -1 0 8740 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_123
timestamp -3599
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp -3599
transform -1 0 8740 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_124
timestamp -3599
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp -3599
transform -1 0 8740 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_125
timestamp -3599
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp -3599
transform -1 0 8740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_126
timestamp -3599
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp -3599
transform -1 0 8740 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_127
timestamp -3599
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp -3599
transform -1 0 8740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_128
timestamp -3599
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp -3599
transform -1 0 8740 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_129
timestamp -3599
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp -3599
transform -1 0 8740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_130
timestamp -3599
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp -3599
transform -1 0 8740 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_131
timestamp -3599
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp -3599
transform -1 0 8740 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_132
timestamp -3599
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp -3599
transform -1 0 8740 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_133
timestamp -3599
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp -3599
transform -1 0 8740 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_134
timestamp -3599
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp -3599
transform -1 0 8740 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_135
timestamp -3599
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp -3599
transform -1 0 8740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_136
timestamp -3599
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp -3599
transform -1 0 8740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_137
timestamp -3599
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp -3599
transform -1 0 8740 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_138
timestamp -3599
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp -3599
transform -1 0 8740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_139
timestamp -3599
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp -3599
transform -1 0 8740 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_140
timestamp -3599
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp -3599
transform -1 0 8740 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_141
timestamp -3599
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp -3599
transform -1 0 8740 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_142
timestamp -3599
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp -3599
transform -1 0 8740 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_143
timestamp -3599
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp -3599
transform -1 0 8740 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_144
timestamp -3599
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp -3599
transform -1 0 8740 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_145
timestamp -3599
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp -3599
transform -1 0 8740 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_146
timestamp -3599
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp -3599
transform -1 0 8740 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_147
timestamp -3599
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp -3599
transform -1 0 8740 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_148
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_149
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_150
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_151
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_152
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_153
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_154
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_155
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_156
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_157
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_158
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_159
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_160
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_161
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_162
timestamp -3599
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp -3599
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_164
timestamp -3599
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp -3599
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_166
timestamp -3599
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_167
timestamp -3599
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_168
timestamp -3599
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp -3599
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_170
timestamp -3599
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_171
timestamp -3599
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_172
timestamp -3599
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_173
timestamp -3599
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_174
timestamp -3599
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_175
timestamp -3599
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_176
timestamp -3599
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_177
timestamp -3599
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_178
timestamp -3599
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_179
timestamp -3599
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_180
timestamp -3599
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_181
timestamp -3599
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_182
timestamp -3599
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_183
timestamp -3599
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_184
timestamp -3599
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_185
timestamp -3599
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_186
timestamp -3599
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_187
timestamp -3599
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_188
timestamp -3599
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_189
timestamp -3599
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_190
timestamp -3599
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_191
timestamp -3599
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_192
timestamp -3599
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_193
timestamp -3599
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_194
timestamp -3599
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_195
timestamp -3599
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_196
timestamp -3599
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_197
timestamp -3599
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_198
timestamp -3599
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_199
timestamp -3599
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_200
timestamp -3599
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_201
timestamp -3599
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_202
timestamp -3599
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_203
timestamp -3599
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_204
timestamp -3599
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_205
timestamp -3599
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_206
timestamp -3599
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_207
timestamp -3599
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_208
timestamp -3599
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_209
timestamp -3599
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_210
timestamp -3599
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_211
timestamp -3599
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_212
timestamp -3599
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_213
timestamp -3599
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_214
timestamp -3599
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_215
timestamp -3599
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_216
timestamp -3599
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_217
timestamp -3599
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_218
timestamp -3599
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_219
timestamp -3599
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_220
timestamp -3599
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_221
timestamp -3599
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_222
timestamp -3599
transform 1 0 3680 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_223
timestamp -3599
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
<< labels >>
flabel metal3 s 9724 18232 9844 18352 0 FreeSans 480 0 0 0 E1BEG[0]
port 0 nsew signal output
flabel metal3 s 9724 18504 9844 18624 0 FreeSans 480 0 0 0 E1BEG[1]
port 1 nsew signal output
flabel metal3 s 9724 18776 9844 18896 0 FreeSans 480 0 0 0 E1BEG[2]
port 2 nsew signal output
flabel metal3 s 9724 19048 9844 19168 0 FreeSans 480 0 0 0 E1BEG[3]
port 3 nsew signal output
flabel metal3 s 9724 19320 9844 19440 0 FreeSans 480 0 0 0 E2BEG[0]
port 4 nsew signal output
flabel metal3 s 9724 19592 9844 19712 0 FreeSans 480 0 0 0 E2BEG[1]
port 5 nsew signal output
flabel metal3 s 9724 19864 9844 19984 0 FreeSans 480 0 0 0 E2BEG[2]
port 6 nsew signal output
flabel metal3 s 9724 20136 9844 20256 0 FreeSans 480 0 0 0 E2BEG[3]
port 7 nsew signal output
flabel metal3 s 9724 20408 9844 20528 0 FreeSans 480 0 0 0 E2BEG[4]
port 8 nsew signal output
flabel metal3 s 9724 20680 9844 20800 0 FreeSans 480 0 0 0 E2BEG[5]
port 9 nsew signal output
flabel metal3 s 9724 20952 9844 21072 0 FreeSans 480 0 0 0 E2BEG[6]
port 10 nsew signal output
flabel metal3 s 9724 21224 9844 21344 0 FreeSans 480 0 0 0 E2BEG[7]
port 11 nsew signal output
flabel metal3 s 9724 21496 9844 21616 0 FreeSans 480 0 0 0 E2BEGb[0]
port 12 nsew signal output
flabel metal3 s 9724 21768 9844 21888 0 FreeSans 480 0 0 0 E2BEGb[1]
port 13 nsew signal output
flabel metal3 s 9724 22040 9844 22160 0 FreeSans 480 0 0 0 E2BEGb[2]
port 14 nsew signal output
flabel metal3 s 9724 22312 9844 22432 0 FreeSans 480 0 0 0 E2BEGb[3]
port 15 nsew signal output
flabel metal3 s 9724 22584 9844 22704 0 FreeSans 480 0 0 0 E2BEGb[4]
port 16 nsew signal output
flabel metal3 s 9724 22856 9844 22976 0 FreeSans 480 0 0 0 E2BEGb[5]
port 17 nsew signal output
flabel metal3 s 9724 23128 9844 23248 0 FreeSans 480 0 0 0 E2BEGb[6]
port 18 nsew signal output
flabel metal3 s 9724 23400 9844 23520 0 FreeSans 480 0 0 0 E2BEGb[7]
port 19 nsew signal output
flabel metal3 s 9724 28024 9844 28144 0 FreeSans 480 0 0 0 E6BEG[0]
port 20 nsew signal output
flabel metal3 s 9724 30744 9844 30864 0 FreeSans 480 0 0 0 E6BEG[10]
port 21 nsew signal output
flabel metal3 s 9724 31016 9844 31136 0 FreeSans 480 0 0 0 E6BEG[11]
port 22 nsew signal output
flabel metal3 s 9724 28296 9844 28416 0 FreeSans 480 0 0 0 E6BEG[1]
port 23 nsew signal output
flabel metal3 s 9724 28568 9844 28688 0 FreeSans 480 0 0 0 E6BEG[2]
port 24 nsew signal output
flabel metal3 s 9724 28840 9844 28960 0 FreeSans 480 0 0 0 E6BEG[3]
port 25 nsew signal output
flabel metal3 s 9724 29112 9844 29232 0 FreeSans 480 0 0 0 E6BEG[4]
port 26 nsew signal output
flabel metal3 s 9724 29384 9844 29504 0 FreeSans 480 0 0 0 E6BEG[5]
port 27 nsew signal output
flabel metal3 s 9724 29656 9844 29776 0 FreeSans 480 0 0 0 E6BEG[6]
port 28 nsew signal output
flabel metal3 s 9724 29928 9844 30048 0 FreeSans 480 0 0 0 E6BEG[7]
port 29 nsew signal output
flabel metal3 s 9724 30200 9844 30320 0 FreeSans 480 0 0 0 E6BEG[8]
port 30 nsew signal output
flabel metal3 s 9724 30472 9844 30592 0 FreeSans 480 0 0 0 E6BEG[9]
port 31 nsew signal output
flabel metal3 s 9724 23672 9844 23792 0 FreeSans 480 0 0 0 EE4BEG[0]
port 32 nsew signal output
flabel metal3 s 9724 26392 9844 26512 0 FreeSans 480 0 0 0 EE4BEG[10]
port 33 nsew signal output
flabel metal3 s 9724 26664 9844 26784 0 FreeSans 480 0 0 0 EE4BEG[11]
port 34 nsew signal output
flabel metal3 s 9724 26936 9844 27056 0 FreeSans 480 0 0 0 EE4BEG[12]
port 35 nsew signal output
flabel metal3 s 9724 27208 9844 27328 0 FreeSans 480 0 0 0 EE4BEG[13]
port 36 nsew signal output
flabel metal3 s 9724 27480 9844 27600 0 FreeSans 480 0 0 0 EE4BEG[14]
port 37 nsew signal output
flabel metal3 s 9724 27752 9844 27872 0 FreeSans 480 0 0 0 EE4BEG[15]
port 38 nsew signal output
flabel metal3 s 9724 23944 9844 24064 0 FreeSans 480 0 0 0 EE4BEG[1]
port 39 nsew signal output
flabel metal3 s 9724 24216 9844 24336 0 FreeSans 480 0 0 0 EE4BEG[2]
port 40 nsew signal output
flabel metal3 s 9724 24488 9844 24608 0 FreeSans 480 0 0 0 EE4BEG[3]
port 41 nsew signal output
flabel metal3 s 9724 24760 9844 24880 0 FreeSans 480 0 0 0 EE4BEG[4]
port 42 nsew signal output
flabel metal3 s 9724 25032 9844 25152 0 FreeSans 480 0 0 0 EE4BEG[5]
port 43 nsew signal output
flabel metal3 s 9724 25304 9844 25424 0 FreeSans 480 0 0 0 EE4BEG[6]
port 44 nsew signal output
flabel metal3 s 9724 25576 9844 25696 0 FreeSans 480 0 0 0 EE4BEG[7]
port 45 nsew signal output
flabel metal3 s 9724 25848 9844 25968 0 FreeSans 480 0 0 0 EE4BEG[8]
port 46 nsew signal output
flabel metal3 s 9724 26120 9844 26240 0 FreeSans 480 0 0 0 EE4BEG[9]
port 47 nsew signal output
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 48 nsew signal input
flabel metal3 s 0 14968 120 15088 0 FreeSans 480 0 0 0 FrameData[10]
port 49 nsew signal input
flabel metal3 s 0 16328 120 16448 0 FreeSans 480 0 0 0 FrameData[11]
port 50 nsew signal input
flabel metal3 s 0 17688 120 17808 0 FreeSans 480 0 0 0 FrameData[12]
port 51 nsew signal input
flabel metal3 s 0 19048 120 19168 0 FreeSans 480 0 0 0 FrameData[13]
port 52 nsew signal input
flabel metal3 s 0 20408 120 20528 0 FreeSans 480 0 0 0 FrameData[14]
port 53 nsew signal input
flabel metal3 s 0 21768 120 21888 0 FreeSans 480 0 0 0 FrameData[15]
port 54 nsew signal input
flabel metal3 s 0 23128 120 23248 0 FreeSans 480 0 0 0 FrameData[16]
port 55 nsew signal input
flabel metal3 s 0 24488 120 24608 0 FreeSans 480 0 0 0 FrameData[17]
port 56 nsew signal input
flabel metal3 s 0 25848 120 25968 0 FreeSans 480 0 0 0 FrameData[18]
port 57 nsew signal input
flabel metal3 s 0 27208 120 27328 0 FreeSans 480 0 0 0 FrameData[19]
port 58 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[1]
port 59 nsew signal input
flabel metal3 s 0 28568 120 28688 0 FreeSans 480 0 0 0 FrameData[20]
port 60 nsew signal input
flabel metal3 s 0 29928 120 30048 0 FreeSans 480 0 0 0 FrameData[21]
port 61 nsew signal input
flabel metal3 s 0 31288 120 31408 0 FreeSans 480 0 0 0 FrameData[22]
port 62 nsew signal input
flabel metal3 s 0 32648 120 32768 0 FreeSans 480 0 0 0 FrameData[23]
port 63 nsew signal input
flabel metal3 s 0 34008 120 34128 0 FreeSans 480 0 0 0 FrameData[24]
port 64 nsew signal input
flabel metal3 s 0 35368 120 35488 0 FreeSans 480 0 0 0 FrameData[25]
port 65 nsew signal input
flabel metal3 s 0 36728 120 36848 0 FreeSans 480 0 0 0 FrameData[26]
port 66 nsew signal input
flabel metal3 s 0 38088 120 38208 0 FreeSans 480 0 0 0 FrameData[27]
port 67 nsew signal input
flabel metal3 s 0 39448 120 39568 0 FreeSans 480 0 0 0 FrameData[28]
port 68 nsew signal input
flabel metal3 s 0 40808 120 40928 0 FreeSans 480 0 0 0 FrameData[29]
port 69 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[2]
port 70 nsew signal input
flabel metal3 s 0 42168 120 42288 0 FreeSans 480 0 0 0 FrameData[30]
port 71 nsew signal input
flabel metal3 s 0 43528 120 43648 0 FreeSans 480 0 0 0 FrameData[31]
port 72 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[3]
port 73 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[4]
port 74 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[5]
port 75 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[6]
port 76 nsew signal input
flabel metal3 s 0 10888 120 11008 0 FreeSans 480 0 0 0 FrameData[7]
port 77 nsew signal input
flabel metal3 s 0 12248 120 12368 0 FreeSans 480 0 0 0 FrameData[8]
port 78 nsew signal input
flabel metal3 s 0 13608 120 13728 0 FreeSans 480 0 0 0 FrameData[9]
port 79 nsew signal input
flabel metal3 s 9724 31288 9844 31408 0 FreeSans 480 0 0 0 FrameData_O[0]
port 80 nsew signal output
flabel metal3 s 9724 34008 9844 34128 0 FreeSans 480 0 0 0 FrameData_O[10]
port 81 nsew signal output
flabel metal3 s 9724 34280 9844 34400 0 FreeSans 480 0 0 0 FrameData_O[11]
port 82 nsew signal output
flabel metal3 s 9724 34552 9844 34672 0 FreeSans 480 0 0 0 FrameData_O[12]
port 83 nsew signal output
flabel metal3 s 9724 34824 9844 34944 0 FreeSans 480 0 0 0 FrameData_O[13]
port 84 nsew signal output
flabel metal3 s 9724 35096 9844 35216 0 FreeSans 480 0 0 0 FrameData_O[14]
port 85 nsew signal output
flabel metal3 s 9724 35368 9844 35488 0 FreeSans 480 0 0 0 FrameData_O[15]
port 86 nsew signal output
flabel metal3 s 9724 35640 9844 35760 0 FreeSans 480 0 0 0 FrameData_O[16]
port 87 nsew signal output
flabel metal3 s 9724 35912 9844 36032 0 FreeSans 480 0 0 0 FrameData_O[17]
port 88 nsew signal output
flabel metal3 s 9724 36184 9844 36304 0 FreeSans 480 0 0 0 FrameData_O[18]
port 89 nsew signal output
flabel metal3 s 9724 36456 9844 36576 0 FreeSans 480 0 0 0 FrameData_O[19]
port 90 nsew signal output
flabel metal3 s 9724 31560 9844 31680 0 FreeSans 480 0 0 0 FrameData_O[1]
port 91 nsew signal output
flabel metal3 s 9724 36728 9844 36848 0 FreeSans 480 0 0 0 FrameData_O[20]
port 92 nsew signal output
flabel metal3 s 9724 37000 9844 37120 0 FreeSans 480 0 0 0 FrameData_O[21]
port 93 nsew signal output
flabel metal3 s 9724 37272 9844 37392 0 FreeSans 480 0 0 0 FrameData_O[22]
port 94 nsew signal output
flabel metal3 s 9724 37544 9844 37664 0 FreeSans 480 0 0 0 FrameData_O[23]
port 95 nsew signal output
flabel metal3 s 9724 37816 9844 37936 0 FreeSans 480 0 0 0 FrameData_O[24]
port 96 nsew signal output
flabel metal3 s 9724 38088 9844 38208 0 FreeSans 480 0 0 0 FrameData_O[25]
port 97 nsew signal output
flabel metal3 s 9724 38360 9844 38480 0 FreeSans 480 0 0 0 FrameData_O[26]
port 98 nsew signal output
flabel metal3 s 9724 38632 9844 38752 0 FreeSans 480 0 0 0 FrameData_O[27]
port 99 nsew signal output
flabel metal3 s 9724 38904 9844 39024 0 FreeSans 480 0 0 0 FrameData_O[28]
port 100 nsew signal output
flabel metal3 s 9724 39176 9844 39296 0 FreeSans 480 0 0 0 FrameData_O[29]
port 101 nsew signal output
flabel metal3 s 9724 31832 9844 31952 0 FreeSans 480 0 0 0 FrameData_O[2]
port 102 nsew signal output
flabel metal3 s 9724 39448 9844 39568 0 FreeSans 480 0 0 0 FrameData_O[30]
port 103 nsew signal output
flabel metal3 s 9724 39720 9844 39840 0 FreeSans 480 0 0 0 FrameData_O[31]
port 104 nsew signal output
flabel metal3 s 9724 32104 9844 32224 0 FreeSans 480 0 0 0 FrameData_O[3]
port 105 nsew signal output
flabel metal3 s 9724 32376 9844 32496 0 FreeSans 480 0 0 0 FrameData_O[4]
port 106 nsew signal output
flabel metal3 s 9724 32648 9844 32768 0 FreeSans 480 0 0 0 FrameData_O[5]
port 107 nsew signal output
flabel metal3 s 9724 32920 9844 33040 0 FreeSans 480 0 0 0 FrameData_O[6]
port 108 nsew signal output
flabel metal3 s 9724 33192 9844 33312 0 FreeSans 480 0 0 0 FrameData_O[7]
port 109 nsew signal output
flabel metal3 s 9724 33464 9844 33584 0 FreeSans 480 0 0 0 FrameData_O[8]
port 110 nsew signal output
flabel metal3 s 9724 33736 9844 33856 0 FreeSans 480 0 0 0 FrameData_O[9]
port 111 nsew signal output
flabel metal2 s 754 0 810 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 112 nsew signal input
flabel metal2 s 5354 0 5410 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 113 nsew signal input
flabel metal2 s 5814 0 5870 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 114 nsew signal input
flabel metal2 s 6274 0 6330 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 115 nsew signal input
flabel metal2 s 6734 0 6790 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 116 nsew signal input
flabel metal2 s 7194 0 7250 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 117 nsew signal input
flabel metal2 s 7654 0 7710 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 118 nsew signal input
flabel metal2 s 8114 0 8170 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 119 nsew signal input
flabel metal2 s 8574 0 8630 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 120 nsew signal input
flabel metal2 s 9034 0 9090 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 121 nsew signal input
flabel metal2 s 9494 0 9550 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 122 nsew signal input
flabel metal2 s 1214 0 1270 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 123 nsew signal input
flabel metal2 s 1674 0 1730 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 124 nsew signal input
flabel metal2 s 2134 0 2190 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 125 nsew signal input
flabel metal2 s 2594 0 2650 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 126 nsew signal input
flabel metal2 s 3054 0 3110 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 127 nsew signal input
flabel metal2 s 3514 0 3570 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 128 nsew signal input
flabel metal2 s 3974 0 4030 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 129 nsew signal input
flabel metal2 s 4434 0 4490 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 130 nsew signal input
flabel metal2 s 4894 0 4950 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 131 nsew signal input
flabel metal2 s 754 44960 810 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 132 nsew signal output
flabel metal2 s 5354 44960 5410 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 133 nsew signal output
flabel metal2 s 5814 44960 5870 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 134 nsew signal output
flabel metal2 s 6274 44960 6330 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 135 nsew signal output
flabel metal2 s 6734 44960 6790 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 136 nsew signal output
flabel metal2 s 7194 44960 7250 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 137 nsew signal output
flabel metal2 s 7654 44960 7710 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 138 nsew signal output
flabel metal2 s 8114 44960 8170 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 139 nsew signal output
flabel metal2 s 8574 44960 8630 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 140 nsew signal output
flabel metal2 s 9034 44960 9090 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 141 nsew signal output
flabel metal2 s 9494 44960 9550 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 142 nsew signal output
flabel metal2 s 1214 44960 1270 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 143 nsew signal output
flabel metal2 s 1674 44960 1730 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 144 nsew signal output
flabel metal2 s 2134 44960 2190 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 145 nsew signal output
flabel metal2 s 2594 44960 2650 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 146 nsew signal output
flabel metal2 s 3054 44960 3110 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 147 nsew signal output
flabel metal2 s 3514 44960 3570 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 148 nsew signal output
flabel metal2 s 3974 44960 4030 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 149 nsew signal output
flabel metal2 s 4434 44960 4490 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 150 nsew signal output
flabel metal2 s 4894 44960 4950 45016 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 151 nsew signal output
flabel metal2 s 294 0 350 56 0 FreeSans 224 0 0 0 UserCLK
port 152 nsew signal input
flabel metal2 s 294 44960 350 45016 0 FreeSans 224 0 0 0 UserCLKo
port 153 nsew signal output
flabel metal4 s 3004 0 3324 45016 0 FreeSans 1920 90 0 0 VGND
port 154 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 154 nsew ground bidirectional
flabel metal4 s 3004 44956 3324 45016 0 FreeSans 480 0 0 0 VGND
port 154 nsew ground bidirectional
flabel metal4 s 1944 0 2264 45016 0 FreeSans 1920 90 0 0 VPWR
port 155 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 155 nsew power bidirectional
flabel metal4 s 1944 44956 2264 45016 0 FreeSans 480 0 0 0 VPWR
port 155 nsew power bidirectional
flabel metal4 s 7944 0 8264 45016 0 FreeSans 1920 90 0 0 VPWR
port 155 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 155 nsew power bidirectional
flabel metal4 s 7944 44956 8264 45016 0 FreeSans 480 0 0 0 VPWR
port 155 nsew power bidirectional
flabel metal3 s 9724 5176 9844 5296 0 FreeSans 480 0 0 0 W1END[0]
port 156 nsew signal input
flabel metal3 s 9724 5448 9844 5568 0 FreeSans 480 0 0 0 W1END[1]
port 157 nsew signal input
flabel metal3 s 9724 5720 9844 5840 0 FreeSans 480 0 0 0 W1END[2]
port 158 nsew signal input
flabel metal3 s 9724 5992 9844 6112 0 FreeSans 480 0 0 0 W1END[3]
port 159 nsew signal input
flabel metal3 s 9724 8440 9844 8560 0 FreeSans 480 0 0 0 W2END[0]
port 160 nsew signal input
flabel metal3 s 9724 8712 9844 8832 0 FreeSans 480 0 0 0 W2END[1]
port 161 nsew signal input
flabel metal3 s 9724 8984 9844 9104 0 FreeSans 480 0 0 0 W2END[2]
port 162 nsew signal input
flabel metal3 s 9724 9256 9844 9376 0 FreeSans 480 0 0 0 W2END[3]
port 163 nsew signal input
flabel metal3 s 9724 9528 9844 9648 0 FreeSans 480 0 0 0 W2END[4]
port 164 nsew signal input
flabel metal3 s 9724 9800 9844 9920 0 FreeSans 480 0 0 0 W2END[5]
port 165 nsew signal input
flabel metal3 s 9724 10072 9844 10192 0 FreeSans 480 0 0 0 W2END[6]
port 166 nsew signal input
flabel metal3 s 9724 10344 9844 10464 0 FreeSans 480 0 0 0 W2END[7]
port 167 nsew signal input
flabel metal3 s 9724 6264 9844 6384 0 FreeSans 480 0 0 0 W2MID[0]
port 168 nsew signal input
flabel metal3 s 9724 6536 9844 6656 0 FreeSans 480 0 0 0 W2MID[1]
port 169 nsew signal input
flabel metal3 s 9724 6808 9844 6928 0 FreeSans 480 0 0 0 W2MID[2]
port 170 nsew signal input
flabel metal3 s 9724 7080 9844 7200 0 FreeSans 480 0 0 0 W2MID[3]
port 171 nsew signal input
flabel metal3 s 9724 7352 9844 7472 0 FreeSans 480 0 0 0 W2MID[4]
port 172 nsew signal input
flabel metal3 s 9724 7624 9844 7744 0 FreeSans 480 0 0 0 W2MID[5]
port 173 nsew signal input
flabel metal3 s 9724 7896 9844 8016 0 FreeSans 480 0 0 0 W2MID[6]
port 174 nsew signal input
flabel metal3 s 9724 8168 9844 8288 0 FreeSans 480 0 0 0 W2MID[7]
port 175 nsew signal input
flabel metal3 s 9724 14968 9844 15088 0 FreeSans 480 0 0 0 W6END[0]
port 176 nsew signal input
flabel metal3 s 9724 17688 9844 17808 0 FreeSans 480 0 0 0 W6END[10]
port 177 nsew signal input
flabel metal3 s 9724 17960 9844 18080 0 FreeSans 480 0 0 0 W6END[11]
port 178 nsew signal input
flabel metal3 s 9724 15240 9844 15360 0 FreeSans 480 0 0 0 W6END[1]
port 179 nsew signal input
flabel metal3 s 9724 15512 9844 15632 0 FreeSans 480 0 0 0 W6END[2]
port 180 nsew signal input
flabel metal3 s 9724 15784 9844 15904 0 FreeSans 480 0 0 0 W6END[3]
port 181 nsew signal input
flabel metal3 s 9724 16056 9844 16176 0 FreeSans 480 0 0 0 W6END[4]
port 182 nsew signal input
flabel metal3 s 9724 16328 9844 16448 0 FreeSans 480 0 0 0 W6END[5]
port 183 nsew signal input
flabel metal3 s 9724 16600 9844 16720 0 FreeSans 480 0 0 0 W6END[6]
port 184 nsew signal input
flabel metal3 s 9724 16872 9844 16992 0 FreeSans 480 0 0 0 W6END[7]
port 185 nsew signal input
flabel metal3 s 9724 17144 9844 17264 0 FreeSans 480 0 0 0 W6END[8]
port 186 nsew signal input
flabel metal3 s 9724 17416 9844 17536 0 FreeSans 480 0 0 0 W6END[9]
port 187 nsew signal input
flabel metal3 s 9724 10616 9844 10736 0 FreeSans 480 0 0 0 WW4END[0]
port 188 nsew signal input
flabel metal3 s 9724 13336 9844 13456 0 FreeSans 480 0 0 0 WW4END[10]
port 189 nsew signal input
flabel metal3 s 9724 13608 9844 13728 0 FreeSans 480 0 0 0 WW4END[11]
port 190 nsew signal input
flabel metal3 s 9724 13880 9844 14000 0 FreeSans 480 0 0 0 WW4END[12]
port 191 nsew signal input
flabel metal3 s 9724 14152 9844 14272 0 FreeSans 480 0 0 0 WW4END[13]
port 192 nsew signal input
flabel metal3 s 9724 14424 9844 14544 0 FreeSans 480 0 0 0 WW4END[14]
port 193 nsew signal input
flabel metal3 s 9724 14696 9844 14816 0 FreeSans 480 0 0 0 WW4END[15]
port 194 nsew signal input
flabel metal3 s 9724 10888 9844 11008 0 FreeSans 480 0 0 0 WW4END[1]
port 195 nsew signal input
flabel metal3 s 9724 11160 9844 11280 0 FreeSans 480 0 0 0 WW4END[2]
port 196 nsew signal input
flabel metal3 s 9724 11432 9844 11552 0 FreeSans 480 0 0 0 WW4END[3]
port 197 nsew signal input
flabel metal3 s 9724 11704 9844 11824 0 FreeSans 480 0 0 0 WW4END[4]
port 198 nsew signal input
flabel metal3 s 9724 11976 9844 12096 0 FreeSans 480 0 0 0 WW4END[5]
port 199 nsew signal input
flabel metal3 s 9724 12248 9844 12368 0 FreeSans 480 0 0 0 WW4END[6]
port 200 nsew signal input
flabel metal3 s 9724 12520 9844 12640 0 FreeSans 480 0 0 0 WW4END[7]
port 201 nsew signal input
flabel metal3 s 9724 12792 9844 12912 0 FreeSans 480 0 0 0 WW4END[8]
port 202 nsew signal input
flabel metal3 s 9724 13064 9844 13184 0 FreeSans 480 0 0 0 WW4END[9]
port 203 nsew signal input
rlabel metal1 4922 42432 4922 42432 0 VGND
rlabel metal1 4922 41888 4922 41888 0 VPWR
rlabel metal3 8856 18292 8856 18292 0 E1BEG[0]
rlabel metal3 9040 18564 9040 18564 0 E1BEG[1]
rlabel metal3 9270 18836 9270 18836 0 E1BEG[2]
rlabel metal3 9408 19108 9408 19108 0 E1BEG[3]
rlabel metal3 8856 19380 8856 19380 0 E2BEG[0]
rlabel metal3 9040 19652 9040 19652 0 E2BEG[1]
rlabel metal3 8810 19924 8810 19924 0 E2BEG[2]
rlabel metal3 9408 20196 9408 20196 0 E2BEG[3]
rlabel metal3 9316 20468 9316 20468 0 E2BEG[4]
rlabel metal3 9040 20740 9040 20740 0 E2BEG[5]
rlabel metal3 8810 21012 8810 21012 0 E2BEG[6]
rlabel metal3 9408 21284 9408 21284 0 E2BEG[7]
rlabel metal3 8856 21556 8856 21556 0 E2BEGb[0]
rlabel metal3 9040 21828 9040 21828 0 E2BEGb[1]
rlabel metal3 8810 22100 8810 22100 0 E2BEGb[2]
rlabel metal3 9408 22372 9408 22372 0 E2BEGb[3]
rlabel metal3 8856 22644 8856 22644 0 E2BEGb[4]
rlabel metal3 9040 22916 9040 22916 0 E2BEGb[5]
rlabel metal3 9316 23188 9316 23188 0 E2BEGb[6]
rlabel metal3 9408 23460 9408 23460 0 E2BEGb[7]
rlabel metal3 9040 28084 9040 28084 0 E6BEG[0]
rlabel metal3 9040 30804 9040 30804 0 E6BEG[10]
rlabel metal3 9316 31076 9316 31076 0 E6BEG[11]
rlabel metal3 8856 28356 8856 28356 0 E6BEG[1]
rlabel metal3 9040 28628 9040 28628 0 E6BEG[2]
rlabel metal3 9362 28900 9362 28900 0 E6BEG[3]
rlabel metal3 9040 29172 9040 29172 0 E6BEG[4]
rlabel metal3 8856 29444 8856 29444 0 E6BEG[5]
rlabel metal3 9040 29716 9040 29716 0 E6BEG[6]
rlabel metal3 9316 29988 9316 29988 0 E6BEG[7]
rlabel metal3 9040 30260 9040 30260 0 E6BEG[8]
rlabel metal3 8856 30532 8856 30532 0 E6BEG[9]
rlabel metal3 8856 23732 8856 23732 0 EE4BEG[0]
rlabel metal3 9040 26452 9040 26452 0 EE4BEG[10]
rlabel metal3 9316 26724 9316 26724 0 EE4BEG[11]
rlabel metal3 9040 26996 9040 26996 0 EE4BEG[12]
rlabel metal3 8856 27268 8856 27268 0 EE4BEG[13]
rlabel metal3 9040 27540 9040 27540 0 EE4BEG[14]
rlabel metal3 9316 27812 9316 27812 0 EE4BEG[15]
rlabel metal3 9040 24004 9040 24004 0 EE4BEG[1]
rlabel metal3 8810 24276 8810 24276 0 EE4BEG[2]
rlabel metal3 9408 24548 9408 24548 0 EE4BEG[3]
rlabel metal3 9040 24820 9040 24820 0 EE4BEG[4]
rlabel metal3 8856 25092 8856 25092 0 EE4BEG[5]
rlabel metal3 9040 25364 9040 25364 0 EE4BEG[6]
rlabel metal3 9431 25636 9431 25636 0 EE4BEG[7]
rlabel metal3 9040 25908 9040 25908 0 EE4BEG[8]
rlabel metal3 9270 26180 9270 26180 0 EE4BEG[9]
rlabel metal3 390 1428 390 1428 0 FrameData[0]
rlabel metal3 436 15028 436 15028 0 FrameData[10]
rlabel metal1 1242 17646 1242 17646 0 FrameData[11]
rlabel metal3 620 17748 620 17748 0 FrameData[12]
rlabel metal3 436 19108 436 19108 0 FrameData[13]
rlabel metal3 528 20468 528 20468 0 FrameData[14]
rlabel metal3 804 21828 804 21828 0 FrameData[15]
rlabel metal3 206 23188 206 23188 0 FrameData[16]
rlabel metal3 482 24548 482 24548 0 FrameData[17]
rlabel metal3 666 25908 666 25908 0 FrameData[18]
rlabel metal3 1264 27268 1264 27268 0 FrameData[19]
rlabel metal1 874 30226 874 30226 0 FrameData[1]
rlabel metal3 712 28628 712 28628 0 FrameData[20]
rlabel metal1 2024 38318 2024 38318 0 FrameData[21]
rlabel via2 114 31348 114 31348 0 FrameData[22]
rlabel metal3 1425 32708 1425 32708 0 FrameData[23]
rlabel metal1 1150 40494 1150 40494 0 FrameData[24]
rlabel metal3 919 35428 919 35428 0 FrameData[25]
rlabel metal2 7498 37315 7498 37315 0 FrameData[26]
rlabel metal3 1425 38148 1425 38148 0 FrameData[27]
rlabel metal2 5566 39457 5566 39457 0 FrameData[28]
rlabel metal3 919 40868 919 40868 0 FrameData[29]
rlabel metal1 1518 30158 1518 30158 0 FrameData[2]
rlabel metal2 7498 41905 7498 41905 0 FrameData[30]
rlabel metal3 3748 43588 3748 43588 0 FrameData[31]
rlabel metal1 1150 31314 1150 31314 0 FrameData[3]
rlabel metal3 1448 6868 1448 6868 0 FrameData[4]
rlabel metal1 1564 32402 1564 32402 0 FrameData[5]
rlabel metal1 1518 32878 1518 32878 0 FrameData[6]
rlabel metal2 828 16116 828 16116 0 FrameData[7]
rlabel metal1 1242 13294 1242 13294 0 FrameData[8]
rlabel metal3 574 13668 574 13668 0 FrameData[9]
rlabel metal2 8326 31501 8326 31501 0 FrameData_O[0]
rlabel metal3 9040 34068 9040 34068 0 FrameData_O[10]
rlabel metal3 9316 34340 9316 34340 0 FrameData_O[11]
rlabel metal3 9040 34612 9040 34612 0 FrameData_O[12]
rlabel metal3 8856 34884 8856 34884 0 FrameData_O[13]
rlabel metal3 9040 35156 9040 35156 0 FrameData_O[14]
rlabel metal3 9316 35428 9316 35428 0 FrameData_O[15]
rlabel metal3 9040 35700 9040 35700 0 FrameData_O[16]
rlabel metal3 8856 35972 8856 35972 0 FrameData_O[17]
rlabel metal3 9040 36244 9040 36244 0 FrameData_O[18]
rlabel metal3 9316 36516 9316 36516 0 FrameData_O[19]
rlabel metal1 8418 31926 8418 31926 0 FrameData_O[1]
rlabel metal3 9040 36788 9040 36788 0 FrameData_O[20]
rlabel metal3 8856 37060 8856 37060 0 FrameData_O[21]
rlabel metal3 9040 37332 9040 37332 0 FrameData_O[22]
rlabel metal3 9316 37604 9316 37604 0 FrameData_O[23]
rlabel metal3 9040 37876 9040 37876 0 FrameData_O[24]
rlabel metal3 8856 38148 8856 38148 0 FrameData_O[25]
rlabel metal3 9040 38420 9040 38420 0 FrameData_O[26]
rlabel metal3 9316 38692 9316 38692 0 FrameData_O[27]
rlabel metal3 9040 38964 9040 38964 0 FrameData_O[28]
rlabel metal3 8856 39236 8856 39236 0 FrameData_O[29]
rlabel metal3 9040 31892 9040 31892 0 FrameData_O[2]
rlabel metal3 9040 39508 9040 39508 0 FrameData_O[30]
rlabel metal3 9316 39780 9316 39780 0 FrameData_O[31]
rlabel metal3 9316 32164 9316 32164 0 FrameData_O[3]
rlabel metal3 9040 32436 9040 32436 0 FrameData_O[4]
rlabel metal3 8856 32708 8856 32708 0 FrameData_O[5]
rlabel metal3 9040 32980 9040 32980 0 FrameData_O[6]
rlabel metal3 9316 33252 9316 33252 0 FrameData_O[7]
rlabel metal3 9040 33524 9040 33524 0 FrameData_O[8]
rlabel metal3 8856 33796 8856 33796 0 FrameData_O[9]
rlabel metal2 782 1401 782 1401 0 FrameStrobe[0]
rlabel metal2 5382 10238 5382 10238 0 FrameStrobe[10]
rlabel metal2 5842 1075 5842 1075 0 FrameStrobe[11]
rlabel metal2 6302 242 6302 242 0 FrameStrobe[12]
rlabel metal2 6762 1738 6762 1738 0 FrameStrobe[13]
rlabel metal2 7222 599 7222 599 0 FrameStrobe[14]
rlabel via2 7682 55 7682 55 0 FrameStrobe[15]
rlabel metal2 8142 55 8142 55 0 FrameStrobe[16]
rlabel metal2 5474 11968 5474 11968 0 FrameStrobe[17]
rlabel metal2 9062 531 9062 531 0 FrameStrobe[18]
rlabel via3 6739 21012 6739 21012 0 FrameStrobe[19]
rlabel metal1 1656 16082 1656 16082 0 FrameStrobe[1]
rlabel metal2 1702 55 1702 55 0 FrameStrobe[2]
rlabel metal1 2254 25874 2254 25874 0 FrameStrobe[3]
rlabel metal1 2070 19822 2070 19822 0 FrameStrobe[4]
rlabel metal2 3082 667 3082 667 0 FrameStrobe[5]
rlabel metal1 3680 19346 3680 19346 0 FrameStrobe[6]
rlabel metal1 3864 21318 3864 21318 0 FrameStrobe[7]
rlabel metal1 4600 19822 4600 19822 0 FrameStrobe[8]
rlabel metal1 4830 16082 4830 16082 0 FrameStrobe[9]
rlabel metal1 1150 41718 1150 41718 0 FrameStrobe_O[0]
rlabel metal1 5474 42330 5474 42330 0 FrameStrobe_O[10]
rlabel metal1 5980 42330 5980 42330 0 FrameStrobe_O[11]
rlabel metal1 6440 42330 6440 42330 0 FrameStrobe_O[12]
rlabel metal2 6762 43652 6762 43652 0 FrameStrobe_O[13]
rlabel metal1 7360 42330 7360 42330 0 FrameStrobe_O[14]
rlabel metal1 7820 42330 7820 42330 0 FrameStrobe_O[15]
rlabel metal1 8234 42330 8234 42330 0 FrameStrobe_O[16]
rlabel metal1 8464 41786 8464 41786 0 FrameStrobe_O[17]
rlabel metal1 8510 41718 8510 41718 0 FrameStrobe_O[18]
rlabel metal1 8924 41242 8924 41242 0 FrameStrobe_O[19]
rlabel metal1 1380 42330 1380 42330 0 FrameStrobe_O[1]
rlabel metal1 1840 42330 1840 42330 0 FrameStrobe_O[2]
rlabel metal1 2300 42330 2300 42330 0 FrameStrobe_O[3]
rlabel metal1 2714 42330 2714 42330 0 FrameStrobe_O[4]
rlabel metal1 2990 42330 2990 42330 0 FrameStrobe_O[5]
rlabel metal1 3496 42330 3496 42330 0 FrameStrobe_O[6]
rlabel metal1 4140 42330 4140 42330 0 FrameStrobe_O[7]
rlabel metal1 4554 42330 4554 42330 0 FrameStrobe_O[8]
rlabel metal1 5060 42330 5060 42330 0 FrameStrobe_O[9]
rlabel metal1 1012 20910 1012 20910 0 UserCLK
rlabel metal1 1058 41786 1058 41786 0 UserCLKo
rlabel metal3 8764 5236 8764 5236 0 W1END[0]
rlabel metal3 8810 5508 8810 5508 0 W1END[1]
rlabel metal2 6394 4403 6394 4403 0 W1END[2]
rlabel metal2 5934 4607 5934 4607 0 W1END[3]
rlabel metal3 9615 8500 9615 8500 0 W2END[0]
rlabel metal3 8442 8772 8442 8772 0 W2END[1]
rlabel metal3 8350 9044 8350 9044 0 W2END[2]
rlabel metal3 9086 9316 9086 9316 0 W2END[3]
rlabel metal3 9040 9588 9040 9588 0 W2END[4]
rlabel metal1 6325 12206 6325 12206 0 W2END[5]
rlabel metal3 9270 10132 9270 10132 0 W2END[6]
rlabel metal3 9362 10404 9362 10404 0 W2END[7]
rlabel via2 9730 6324 9730 6324 0 W2MID[0]
rlabel metal3 8534 6596 8534 6596 0 W2MID[1]
rlabel metal2 6762 5729 6762 5729 0 W2MID[2]
rlabel metal2 5842 6477 5842 6477 0 W2MID[3]
rlabel metal3 8488 7412 8488 7412 0 W2MID[4]
rlabel metal1 7912 6766 7912 6766 0 W2MID[5]
rlabel metal3 8396 7956 8396 7956 0 W2MID[6]
rlabel metal3 9086 8228 9086 8228 0 W2MID[7]
rlabel metal1 8188 18326 8188 18326 0 W6END[0]
rlabel metal3 9086 17748 9086 17748 0 W6END[10]
rlabel metal3 9362 18020 9362 18020 0 W6END[11]
rlabel metal2 6486 17391 6486 17391 0 W6END[1]
rlabel metal2 5106 18003 5106 18003 0 W6END[2]
rlabel metal2 6762 18513 6762 18513 0 W6END[3]
rlabel metal3 4669 16116 4669 16116 0 W6END[4]
rlabel metal3 7384 16388 7384 16388 0 W6END[5]
rlabel metal3 9454 16660 9454 16660 0 W6END[6]
rlabel metal3 9546 16932 9546 16932 0 W6END[7]
rlabel metal3 9638 17204 9638 17204 0 W6END[8]
rlabel metal3 9224 17476 9224 17476 0 W6END[9]
rlabel metal3 8143 10676 8143 10676 0 WW4END[0]
rlabel metal3 9270 13396 9270 13396 0 WW4END[10]
rlabel metal1 6647 16082 6647 16082 0 WW4END[11]
rlabel metal3 9592 13940 9592 13940 0 WW4END[12]
rlabel metal1 6946 17102 6946 17102 0 WW4END[13]
rlabel metal1 7176 17646 7176 17646 0 WW4END[14]
rlabel metal1 8004 18258 8004 18258 0 WW4END[15]
rlabel metal3 3243 11084 3243 11084 0 WW4END[1]
rlabel metal3 8947 20604 8947 20604 0 WW4END[2]
rlabel metal3 9224 11492 9224 11492 0 WW4END[3]
rlabel metal3 9615 11764 9615 11764 0 WW4END[4]
rlabel metal3 9684 12036 9684 12036 0 WW4END[5]
rlabel metal3 9270 12308 9270 12308 0 WW4END[6]
rlabel metal3 9638 12580 9638 12580 0 WW4END[7]
rlabel metal1 6831 14382 6831 14382 0 WW4END[8]
rlabel metal3 9132 13124 9132 13124 0 WW4END[9]
rlabel metal2 6118 10880 6118 10880 0 net1
rlabel via3 6187 13804 6187 13804 0 net10
rlabel via3 5037 41412 5037 41412 0 net100
rlabel metal1 1932 41582 1932 41582 0 net101
rlabel metal2 3818 12716 3818 12716 0 net11
rlabel metal1 7544 18938 7544 18938 0 net12
rlabel via3 8395 17612 8395 17612 0 net13
rlabel metal1 6716 20774 6716 20774 0 net14
rlabel metal2 2714 17544 2714 17544 0 net15
rlabel metal1 6992 22542 6992 22542 0 net16
rlabel metal2 6992 17204 6992 17204 0 net17
rlabel metal3 7291 17884 7291 17884 0 net18
rlabel metal1 6256 9146 6256 9146 0 net19
rlabel metal1 6440 3162 6440 3162 0 net2
rlabel metal1 7774 23290 7774 23290 0 net20
rlabel metal1 7912 28186 7912 28186 0 net21
rlabel metal1 7406 31246 7406 31246 0 net22
rlabel via3 7291 22100 7291 22100 0 net23
rlabel metal1 7590 19482 7590 19482 0 net24
rlabel metal1 7774 28730 7774 28730 0 net25
rlabel metal1 7544 29138 7544 29138 0 net26
rlabel metal1 8142 29580 8142 29580 0 net27
rlabel metal2 7774 29818 7774 29818 0 net28
rlabel metal1 8004 30226 8004 30226 0 net29
rlabel metal2 3910 11696 3910 11696 0 net3
rlabel metal2 7406 30940 7406 30940 0 net30
rlabel metal2 6992 22644 6992 22644 0 net31
rlabel metal2 5290 21325 5290 21325 0 net32
rlabel metal1 7268 18394 7268 18394 0 net33
rlabel metal2 7498 25772 7498 25772 0 net34
rlabel metal1 7590 25466 7590 25466 0 net35
rlabel metal2 7222 26690 7222 26690 0 net36
rlabel metal1 7406 26554 7406 26554 0 net37
rlabel metal1 7682 27098 7682 27098 0 net38
rlabel metal1 7728 27642 7728 27642 0 net39
rlabel metal2 5290 11152 5290 11152 0 net4
rlabel metal1 6624 17850 6624 17850 0 net40
rlabel metal1 7084 17306 7084 17306 0 net41
rlabel metal2 7682 24548 7682 24548 0 net42
rlabel metal1 6302 17714 6302 17714 0 net43
rlabel metal2 7636 19244 7636 19244 0 net44
rlabel metal2 6532 20604 6532 20604 0 net45
rlabel metal2 7912 19788 7912 19788 0 net46
rlabel metal1 7866 19210 7866 19210 0 net47
rlabel metal1 7958 13498 7958 13498 0 net48
rlabel metal1 8004 31790 8004 31790 0 net49
rlabel metal1 6256 8602 6256 8602 0 net5
rlabel metal1 2300 15674 2300 15674 0 net50
rlabel metal2 1794 26214 1794 26214 0 net51
rlabel metal1 2668 19482 2668 19482 0 net52
rlabel metal1 2668 21658 2668 21658 0 net53
rlabel metal1 7176 35598 7176 35598 0 net54
rlabel metal2 4370 34646 4370 34646 0 net55
rlabel metal2 5382 35666 5382 35666 0 net56
rlabel metal1 2507 36278 2507 36278 0 net57
rlabel metal1 6072 36686 6072 36686 0 net58
rlabel metal1 2691 36890 2691 36890 0 net59
rlabel metal1 7682 19890 7682 19890 0 net6
rlabel metal1 7636 31790 7636 31790 0 net60
rlabel metal1 6808 37094 6808 37094 0 net61
rlabel metal1 7774 37196 7774 37196 0 net62
rlabel metal1 8142 37876 8142 37876 0 net63
rlabel metal2 7682 36550 7682 36550 0 net64
rlabel metal2 5750 39372 5750 39372 0 net65
rlabel metal1 7728 37434 7728 37434 0 net66
rlabel metal1 7774 37978 7774 37978 0 net67
rlabel metal1 7728 38522 7728 38522 0 net68
rlabel metal1 8142 39372 8142 39372 0 net69
rlabel metal2 7774 13532 7774 13532 0 net7
rlabel metal1 7820 39406 7820 39406 0 net70
rlabel metal1 7682 32334 7682 32334 0 net71
rlabel metal1 7774 41446 7774 41446 0 net72
rlabel metal2 7774 40460 7774 40460 0 net73
rlabel metal1 5014 31450 5014 31450 0 net74
rlabel metal1 3266 31994 3266 31994 0 net75
rlabel metal1 5290 32538 5290 32538 0 net76
rlabel metal2 7866 33286 7866 33286 0 net77
rlabel metal2 7774 33660 7774 33660 0 net78
rlabel metal2 1886 13651 1886 13651 0 net79
rlabel metal3 7705 20332 7705 20332 0 net8
rlabel metal1 2300 14586 2300 14586 0 net80
rlabel via3 1725 41412 1725 41412 0 net81
rlabel metal1 5704 42194 5704 42194 0 net82
rlabel metal1 5382 29002 5382 29002 0 net83
rlabel metal1 5566 42126 5566 42126 0 net84
rlabel via2 3542 19499 3542 19499 0 net85
rlabel metal1 7314 42126 7314 42126 0 net86
rlabel metal1 7774 42092 7774 42092 0 net87
rlabel metal1 7038 42228 7038 42228 0 net88
rlabel metal1 7498 21896 7498 21896 0 net89
rlabel metal3 6187 11628 6187 11628 0 net9
rlabel metal1 7452 41514 7452 41514 0 net90
rlabel metal1 6900 21862 6900 21862 0 net91
rlabel metal3 1633 41684 1633 41684 0 net92
rlabel metal1 1702 23834 1702 23834 0 net93
rlabel metal1 2438 26010 2438 26010 0 net94
rlabel metal2 2622 31110 2622 31110 0 net95
rlabel metal1 3358 42194 3358 42194 0 net96
rlabel metal2 3634 30838 3634 30838 0 net97
rlabel metal1 3956 42194 3956 42194 0 net98
rlabel metal1 4876 42194 4876 42194 0 net99
<< properties >>
string FIXED_BBOX 0 0 9844 45016
<< end >>
