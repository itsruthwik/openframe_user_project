* NGSPICE file created from RegFile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

.subckt RegFile E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2] E1END[3]
+ E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0]
+ E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7] E2END[0] E2END[1]
+ E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0] E2MID[1] E2MID[2]
+ E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1]
+ E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] E6END[0]
+ E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5] E6END[6] E6END[7]
+ E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13] EE4BEG[14]
+ EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6] EE4BEG[7]
+ EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13] EE4END[14]
+ EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6] EE4END[7]
+ EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S1END[0]
+ S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5]
+ S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6]
+ S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7]
+ S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4BEG[0]
+ S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3]
+ S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0] W1BEG[1] W1BEG[2]
+ W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1] W2BEG[2] W2BEG[3]
+ W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2] W2BEGb[3] W2BEGb[4]
+ W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5]
+ W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6]
+ W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4] W6BEG[5]
+ W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11] W6END[1] W6END[2]
+ W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9] WW4BEG[0] WW4BEG[10]
+ WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1] WW4BEG[2] WW4BEG[3]
+ WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9] WW4END[0] WW4END[10]
+ WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1] WW4END[2] WW4END[3]
+ WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2106_ net559 net609 _0935_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__mux2_4
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2037_ net77 net20 Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q VGND VGND VPWR VPWR
+ _0891_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2939_ NN4END[15] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_20_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1270_ _0145_ _0173_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__a21o_1
XFILLER_76_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2724_ net764 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2655_ net770 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1606_ Inst_RegFile_32x4.mem\[4\]\[2\] Inst_RegFile_32x4.mem\[5\]\[2\] net620 VGND
+ VGND VPWR VPWR _0526_ sky130_fd_sc_hd__mux2_1
X_2586_ net775 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1537_ net644 _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__and2b_1
XFILLER_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1468_ Inst_RegFile_32x4.mem\[28\]\[0\] Inst_RegFile_32x4.mem\[29\]\[0\] net624 VGND
+ VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux2_1
XFILLER_86_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1399_ net59 net67 net2 net10 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__mux4_2
XFILLER_67_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold170 Inst_RegFile_32x4.mem\[9\]\[0\] VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold181 Inst_RegFile_32x4.mem\[23\]\[0\] VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout650 AD3 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__buf_8
Xfanout683 net684 VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__clkbuf_4
Xfanout672 net674 VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__buf_2
Xfanout661 AD1 VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__buf_8
Xfanout694 net695 VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2440_ net46 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2371_ net765 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1322_ _0244_ _0234_ _0259_ _0209_ VGND VGND VPWR VPWR Inst_RegFile_32x4.AD_comb\[1\]
+ sky130_fd_sc_hd__a2bb2o_4
X_1253_ net117 net674 net660 net656 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux4_1
XFILLER_76_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1184_ Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q _0128_ VGND VGND VPWR VPWR _0129_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2707_ net749 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput231 net231 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput220 net220 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput242 net242 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__buf_8
Xoutput253 net253 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
X_2638_ net757 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput286 net286 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput275 net275 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput264 net264 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_2
X_2569_ net758 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput297 net297 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__buf_6
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1940_ _0818_ _0817_ _0819_ Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q VGND VGND
+ VPWR VPWR _0820_ sky130_fd_sc_hd__a22o_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1871_ _0756_ _1022_ _0758_ Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q VGND VGND
+ VPWR VPWR _0759_ sky130_fd_sc_hd__o211a_1
X_2423_ net778 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2354_ net54 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1305_ net662 _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__nand2_1
XFILLER_84_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2285_ clknet_4_8_0_UserCLK_regs _0043_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[22\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1236_ Inst_RegFile_32x4.mem\[4\]\[0\] Inst_RegFile_32x4.mem\[5\]\[0\] net394 VGND
+ VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
XFILLER_37_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1167_ Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q _1054_ _1055_ _1058_ VGND VGND
+ VPWR VPWR _1059_ sky130_fd_sc_hd__a31o_1
XFILLER_64_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1098_ Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__inv_2
XFILLER_20_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2070_ _0884_ _0919_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__nor2_4
XFILLER_81_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2972_ S4END[12] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1923_ net402 _0804_ Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q VGND VGND VPWR VPWR
+ _0805_ sky130_fd_sc_hd__mux2_2
XFILLER_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1854_ Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q _0742_ VGND VGND VPWR VPWR _0743_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1785_ net74 net102 net17 Inst_RegFile_switch_matrix.JS2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__mux4_2
X_2406_ net762 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2337_ net40 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2268_ clknet_4_12_0_UserCLK_regs _0026_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[30\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1219_ Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q _0161_ _0158_ _0156_ VGND VGND
+ VPWR VPWR _0162_ sky130_fd_sc_hd__a2bb2o_4
X_2199_ net604 net521 _0959_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__mux2_4
XFILLER_25_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold74 Inst_RegFile_32x4.mem\[18\]\[2\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 Inst_RegFile_32x4.mem\[14\]\[2\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold85 Inst_RegFile_32x4.mem\[8\]\[0\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 Inst_RegFile_32x4.mem\[28\]\[0\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_5 E6END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1570_ Inst_RegFile_32x4.mem\[2\]\[3\] Inst_RegFile_32x4.mem\[3\]\[3\] net622 VGND
+ VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux2_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2122_ net600 net567 _0940_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux2_4
XFILLER_66_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer39 net669 VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__buf_6
XFILLER_66_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2053_ net106 Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q
+ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__o211a_1
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2955_ Inst_RegFile_switch_matrix.JS2BEG7 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_60_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2886_ FrameStrobe[14] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_1
X_1906_ net61 net783 net89 net413 Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q
+ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__mux4_1
X_1837_ _0723_ _0728_ Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.SS4BEG3 sky130_fd_sc_hd__mux2_2
X_1768_ net680 net633 net665 net638 Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__mux4_2
X_1699_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q _0606_ VGND VGND VPWR VPWR _0607_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput120 W2END[2] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_4
Xinput131 W2MID[5] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2740_ clknet_4_11_0_UserCLK_regs _0076_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[19\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2671_ net754 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1622_ _0534_ _0536_ _0539_ _0969_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG4
+ sky130_fd_sc_hd__a22o_4
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1553_ _0471_ _0474_ net645 VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
X_1484_ Inst_RegFile_32x4.mem\[16\]\[0\] Inst_RegFile_32x4.mem\[17\]\[0\] net627 VGND
+ VGND VPWR VPWR _0410_ sky130_fd_sc_hd__mux2_1
XFILLER_86_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2105_ _0930_ _0924_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__nor2_8
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2036_ net76 net104 net132 Inst_RegFile_switch_matrix.JN2BEG3 Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_37_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2938_ NN4END[14] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_20_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2869_ net47 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2723_ net765 net744 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2654_ net771 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1605_ net643 _0524_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__and2b_1
X_2585_ net776 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1536_ _0459_ _0458_ net685 VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__mux2_1
X_1467_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__inv_8
X_1398_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q _0329_ Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__o21a_1
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2019_ _0872_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__inv_1
XFILLER_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold160 Inst_RegFile_32x4.mem\[10\]\[1\] VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 Inst_RegFile_32x4.mem\[29\]\[3\] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 Inst_RegFile_32x4.mem\[23\]\[3\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout651 _0169_ VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__buf_6
Xfanout640 BD3 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__buf_6
Xfanout673 net674 VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__buf_2
Xfanout662 net663 VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__buf_8
Xfanout684 BD0 VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__clkbuf_4
Xfanout695 net696 VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2370_ net766 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1321_ _0251_ _0258_ net393 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__mux2_1
X_1252_ _0183_ _0184_ _1006_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a22o_1
XFILLER_49_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1183_ net75 net18 net103 net131 Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q
+ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__mux4_2
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2706_ net751 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput210 net210 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2637_ net769 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput221 net221 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput232 net232 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput243 Inst_RegFile_switch_matrix.N1BEG3 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__buf_6
Xoutput265 Inst_RegFile_switch_matrix.N4BEG2 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__buf_6
Xoutput276 net276 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput254 net254 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__buf_2
X_2568_ net759 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput287 net287 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput298 net298 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__buf_8
X_2499_ net765 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1519_ _0441_ _0442_ net688 VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__mux2_1
XFILLER_74_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1870_ Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q _0757_ VGND VGND VPWR VPWR _0758_
+ sky130_fd_sc_hd__or2_1
XFILLER_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2422_ net779 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2353_ net752 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1304_ _0241_ _0240_ net675 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_4
X_2284_ clknet_4_10_0_UserCLK_regs _0042_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[22\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1235_ net445 _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__nor2_1
XFILLER_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1166_ Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q _1057_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__o21ai_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1097_ net691 VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__inv_1
X_1999_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _0852_ _0850_ VGND VGND VPWR VPWR
+ _0853_ sky130_fd_sc_hd__a21oi_4
XFILLER_85_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_6_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2971_ S4END[11] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_2
X_1922_ net82 net92 net7 net120 Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q
+ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__mux4_2
X_1853_ _0698_ _0378_ Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q VGND VGND VPWR VPWR
+ _0742_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1784_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__inv_2
XFILLER_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2405_ net763 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2336_ net39 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2267_ clknet_4_13_0_UserCLK_regs _0025_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[30\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1218_ _0159_ _0160_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q VGND VGND VPWR VPWR
+ _0161_ sky130_fd_sc_hd__mux2_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2198_ net608 net490 _0959_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__mux2_4
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1149_ Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q _1041_ VGND VGND VPWR VPWR _1042_
+ sky130_fd_sc_hd__nor2_1
XFILLER_80_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold64 Inst_RegFile_32x4.mem\[4\]\[3\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold75 Inst_RegFile_32x4.mem\[8\]\[2\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 Inst_RegFile_32x4.mem\[14\]\[0\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 Inst_RegFile_32x4.mem\[26\]\[3\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_6 E6END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2121_ net630 net546 _0940_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__mux2_4
X_2052_ Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q _0598_ VGND VGND VPWR VPWR _0903_
+ sky130_fd_sc_hd__nand2_1
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2954_ Inst_RegFile_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_60_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2885_ FrameStrobe[13] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_1
X_1905_ _0683_ _0559_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q VGND VGND VPWR VPWR
+ _0789_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1836_ _0724_ _0725_ _0727_ Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q VGND VGND
+ VPWR VPWR _0728_ sky130_fd_sc_hd__a22o_1
X_1767_ net690 net652 net415 net646 Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__mux4_1
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1698_ net134 net671 net653 net647 Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q
+ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__mux4_1
XFILLER_57_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2319_ net754 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput110 SS4END[0] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_4
Xinput132 W2MID[6] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
Xinput121 W2END[3] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_2
XFILLER_48_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2670_ net757 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1621_ _0537_ _0538_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q VGND VGND VPWR VPWR
+ _0539_ sky130_fd_sc_hd__mux2_1
X_1552_ _0472_ _0473_ net687 VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
X_1483_ _0408_ _0405_ Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q VGND VGND VPWR VPWR
+ _0409_ sky130_fd_sc_hd__mux2_4
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2104_ net601 net462 _0934_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__mux2_4
X_2035_ _0775_ _0827_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q VGND VGND VPWR VPWR
+ _0889_ sky130_fd_sc_hd__mux2_4
XFILLER_54_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2937_ NN4END[13] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_20_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2868_ net46 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
X_1819_ net58 net86 net114 net646 Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q
+ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__mux4_1
X_2799_ Inst_RegFile_switch_matrix.E2BEG3 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_1
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_79_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2722_ net766 net744 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2653_ net772 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1604_ _0523_ _0522_ net685 VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__mux2_1
X_2584_ net777 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1535_ Inst_RegFile_32x4.mem\[0\]\[1\] Inst_RegFile_32x4.mem\[1\]\[1\] net622 VGND
+ VGND VPWR VPWR _0459_ sky130_fd_sc_hd__mux2_1
XFILLER_59_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1466_ _0392_ _0379_ Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q VGND VGND VPWR VPWR
+ _0393_ sky130_fd_sc_hd__mux2_4
X_1397_ net115 net672 net658 net654 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__mux4_1
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2018_ net77 net20 Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q VGND VGND VPWR VPWR
+ _0872_ sky130_fd_sc_hd__mux2_1
XFILLER_82_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold150 Inst_RegFile_32x4.mem\[22\]\[2\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold161 Inst_RegFile_32x4.mem\[29\]\[1\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 Inst_RegFile_32x4.mem\[17\]\[3\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 Inst_RegFile_32x4.mem\[25\]\[2\] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout641 net642 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__buf_8
Xfanout630 net632 VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__clkbuf_4
Xfanout685 net686 VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__clkbuf_4
Xfanout652 net653 VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__buf_8
Xfanout674 AD0 VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__buf_2
Xfanout663 net664 VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__buf_8
XFILLER_73_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout696 net697 VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__buf_2
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1320_ _0254_ _0257_ net664 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__mux2_1
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1251_ _0191_ Inst_RegFile_switch_matrix.JN2BEG5 Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q
+ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_4
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1182_ net433 VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__inv_2
XFILLER_49_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2705_ net752 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput200 net200 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
X_2636_ net780 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput222 net222 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput233 net233 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput244 net244 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__buf_8
Xoutput211 net211 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput277 net277 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput266 net266 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_6
Xoutput255 net255 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__buf_2
X_2567_ net45 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput288 net288 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput299 net299 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__buf_8
X_2498_ net766 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1518_ Inst_RegFile_32x4.mem\[18\]\[1\] Inst_RegFile_32x4.mem\[19\]\[1\] net627 VGND
+ VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux2_1
X_1449_ net82 net782 net118 Inst_RegFile_switch_matrix.JW2BEG4 Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux4_2
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_14_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_14_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2421_ net747 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2352_ net753 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1303_ Inst_RegFile_32x4.mem\[6\]\[1\] Inst_RegFile_32x4.mem\[7\]\[1\] net394 VGND
+ VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_2
X_2283_ clknet_4_10_0_UserCLK_regs _0041_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[22\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1234_ Inst_RegFile_32x4.mem\[2\]\[0\] Inst_RegFile_32x4.mem\[3\]\[0\] net615 VGND
+ VGND VPWR VPWR _0176_ sky130_fd_sc_hd__mux2_1
XFILLER_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1165_ _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__inv_1
XFILLER_37_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1096_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__inv_1
XFILLER_20_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1998_ _0708_ _0851_ Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q VGND VGND VPWR VPWR
+ _0852_ sky130_fd_sc_hd__mux2_2
X_2619_ net774 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2970_ S4END[10] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__buf_2
X_1921_ Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q _1072_ Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q
+ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1852_ _0737_ _0741_ Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.SS4BEG1 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_12_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1783_ _0998_ _0983_ _0979_ _0138_ Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q
+ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__mux4_2
XFILLER_6_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2404_ net764 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2335_ net770 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2266_ clknet_4_13_0_UserCLK_regs _0024_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[30\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1217_ net86 net96 net88 net693 Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q
+ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__mux4_1
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2197_ _0958_ _0886_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__nand2_8
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1148_ _0970_ _0989_ Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q VGND VGND VPWR VPWR
+ _1041_ sky130_fd_sc_hd__mux2_1
XFILLER_37_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1079_ Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__inv_2
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold65 Inst_RegFile_32x4.mem\[18\]\[3\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold98 Inst_RegFile_32x4.mem\[4\]\[0\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 Inst_RegFile_32x4.mem\[10\]\[3\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 Inst_RegFile_32x4.mem\[12\]\[0\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_71_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_7 E6END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2120_ net604 net576 _0940_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__mux2_4
X_2051_ net485 net631 _0888_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_77_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1904_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q _0681_ _0787_ Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q
+ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_60_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2884_ net734 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
X_1835_ _0352_ _0726_ Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q VGND VGND VPWR VPWR
+ _0727_ sky130_fd_sc_hd__mux2_2
X_1766_ _0661_ _0665_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG7 sky130_fd_sc_hd__nand2_2
X_1697_ _0602_ _0600_ _0605_ _1012_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ net757 net734 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2249_ clknet_4_13_0_UserCLK_regs _0007_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[25\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput111 SS4END[1] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_4
Xinput100 S2MID[2] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
Xinput122 W2END[4] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_4
Xinput133 W2MID[7] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1620_ net10 net87 net95 net115 Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__mux4_1
X_1551_ Inst_RegFile_32x4.mem\[30\]\[3\] Inst_RegFile_32x4.mem\[31\]\[3\] net628 VGND
+ VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
X_1482_ net64 net92 _0406_ _0407_ Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q
+ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux4_2
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2103_ net629 net513 _0934_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_65_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ _0887_ _0855_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__nor2_8
X_2936_ NN4END[12] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__buf_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2867_ net760 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_20_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1818_ Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q _0710_ _0712_ VGND VGND VPWR VPWR
+ _0713_ sky130_fd_sc_hd__and3_1
X_2798_ Inst_RegFile_switch_matrix.E2BEG2 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_6
X_1749_ _0646_ _0647_ _0650_ _1018_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG7
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2721_ net767 net746 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2652_ net773 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1603_ Inst_RegFile_32x4.mem\[0\]\[2\] Inst_RegFile_32x4.mem\[1\]\[2\] net622 VGND
+ VGND VPWR VPWR _0523_ sky130_fd_sc_hd__mux2_1
X_2583_ net778 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1534_ Inst_RegFile_32x4.mem\[2\]\[1\] Inst_RegFile_32x4.mem\[3\]\[1\] net622 VGND
+ VGND VPWR VPWR _0458_ sky130_fd_sc_hd__mux2_1
X_1465_ _0985_ _0387_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__a21o_1
X_1396_ _0327_ _0977_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__or2_4
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2017_ Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q _0868_ _0870_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q
+ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__a211o_1
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2919_ N4END[11] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold162 Inst_RegFile_32x4.mem\[16\]\[3\] VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 Inst_RegFile_32x4.mem\[12\]\[1\] VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold140 Inst_RegFile_32x4.mem\[25\]\[0\] VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 Inst_RegFile_32x4.mem\[17\]\[2\] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 Inst_RegFile_32x4.mem\[13\]\[1\] VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout620 net625 VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__buf_8
Xfanout642 BD3 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__buf_8
Xfanout631 net632 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__buf_2
Xfanout675 net677 VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__buf_8
Xfanout664 _0142_ VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__buf_8
Xfanout653 net656 VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__buf_8
Xfanout697 FrameStrobe[9] VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__buf_2
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout686 net687 VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__clkbuf_4
XFILLER_73_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1250_ net62 net90 net24 net118 Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q
+ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux4_2
XFILLER_49_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1181_ _0998_ _0983_ _0980_ _1071_ Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q
+ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__mux4_2
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2704_ net753 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2635_ net50 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput201 net201 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
Xoutput234 net234 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput223 net223 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput212 net212 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput267 net267 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput256 net256 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_8
X_2566_ net762 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput278 net278 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput289 net289 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__buf_2
X_1517_ Inst_RegFile_32x4.mem\[16\]\[1\] Inst_RegFile_32x4.mem\[17\]\[1\] net627 VGND
+ VGND VPWR VPWR _0441_ sky130_fd_sc_hd__mux2_1
X_2497_ net767 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1448_ _0376_ _0373_ Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JW2BEG4 sky130_fd_sc_hd__mux2_4
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1379_ _0312_ _0308_ net651 VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__or3_4
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2420_ net748 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2351_ net754 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2282_ clknet_4_10_0_UserCLK_regs _0040_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[22\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1302_ Inst_RegFile_32x4.mem\[4\]\[1\] Inst_RegFile_32x4.mem\[5\]\[1\] net394 VGND
+ VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_4
XFILLER_84_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1233_ _0174_ net446 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__and2b_1
XFILLER_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1164_ net84 net7 Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q VGND VGND VPWR VPWR
+ _1056_ sky130_fd_sc_hd__mux2_1
XFILLER_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1095_ net15 VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__inv_2
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1997_ net83 net24 net107 Inst_RegFile_switch_matrix.JS2BEG2 Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__mux4_1
XFILLER_9_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2618_ net775 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_7_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2549_ net747 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_85_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1920_ Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q net683 VGND VGND VPWR VPWR _0802_
+ sky130_fd_sc_hd__or2_1
X_1851_ _0739_ _0738_ _0740_ Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q VGND VGND
+ VPWR VPWR _0741_ sky130_fd_sc_hd__a22o_1
X_1782_ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q _0678_ _0679_ VGND VGND VPWR VPWR
+ _0680_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2403_ net765 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2334_ net771 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2265_ clknet_4_7_0_UserCLK_regs _0023_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1216_ net60 net68 net784 net11 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux4_1
X_2196_ _0932_ net437 VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__nor2_8
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1147_ net100 Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q
+ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__o21a_1
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1078_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__inv_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold88 Inst_RegFile_32x4.mem\[16\]\[0\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 Inst_RegFile_32x4.mem\[7\]\[2\] VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 Inst_RegFile_32x4.mem\[26\]\[0\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 Inst_RegFile_32x4.mem\[22\]\[1\] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 E6END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_2_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_2_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2050_ _0682_ _0706_ _0407_ _0901_ Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q
+ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_77_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2952_ Inst_RegFile_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_6
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1903_ Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q net398 VGND VGND VPWR VPWR _0787_
+ sky130_fd_sc_hd__nor2_1
XFILLER_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2883_ net738 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_60_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1834_ net62 net90 net5 net139 Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q
+ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__mux4_2
X_1765_ Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q _0664_ VGND VGND VPWR VPWR _0665_
+ sky130_fd_sc_hd__nand2b_1
X_1696_ _0603_ _0604_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q VGND VGND VPWR VPWR
+ _0605_ sky130_fd_sc_hd__mux2_1
X_2317_ clknet_4_8_0_UserCLK_regs _0075_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[21\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ clknet_4_12_0_UserCLK_regs _0006_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[25\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2179_ net545 net631 _0954_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux2_4
XFILLER_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput101 S2MID[3] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
Xinput112 SS4END[2] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput123 W2END[5] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__buf_2
Xinput134 W6END[0] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1550_ Inst_RegFile_32x4.mem\[28\]\[3\] Inst_RegFile_32x4.mem\[29\]\[3\] net624 VGND
+ VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux2_1
X_1481_ net75 net18 net103 net131 Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux4_2
XFILLER_79_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2102_ net605 net482 _0934_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_65_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2033_ _0884_ _0879_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__or2_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2935_ NN4END[11] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_1
X_2866_ net761 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
X_1817_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q _1045_ _0711_ Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q
+ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_20_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2797_ Inst_RegFile_switch_matrix.E2BEG1 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_6
X_1748_ _0648_ _0649_ _1017_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux2_1
X_1679_ _0586_ _0584_ _0589_ _1008_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG2
+ sky130_fd_sc_hd__a22o_4
XFILLER_85_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2720_ net768 net746 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2651_ net774 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1602_ Inst_RegFile_32x4.mem\[2\]\[2\] Inst_RegFile_32x4.mem\[3\]\[2\] net622 VGND
+ VGND VPWR VPWR _0522_ sky130_fd_sc_hd__mux2_1
X_2582_ net779 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1533_ net417 _0450_ _0452_ _0393_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__o31a_1
X_1464_ _0988_ _0390_ _0389_ Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q VGND VGND
+ VPWR VPWR _0391_ sky130_fd_sc_hd__o211a_1
X_1395_ net648 net636 net668 net447 Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q
+ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__mux4_2
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2016_ Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q _0869_ VGND VGND VPWR VPWR _0870_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_33_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2918_ N4END[10] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_1
X_2849_ net56 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
Xhold141 Inst_RegFile_32x4.mem\[5\]\[1\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold130 Inst_RegFile_32x4.mem\[28\]\[3\] VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 Inst_RegFile_32x4.mem\[31\]\[1\] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 Inst_RegFile_32x4.mem\[23\]\[2\] VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 Inst_RegFile_32x4.mem\[19\]\[1\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 Inst_RegFile_32x4.mem\[21\]\[3\] VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout621 net625 VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__clkbuf_2
Xfanout632 _0902_ VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__clkbuf_2
Xfanout610 net611 VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__buf_2
Xfanout654 net655 VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__buf_8
Xfanout665 net666 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__buf_8
Xfanout643 net644 VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__buf_8
Xfanout676 net677 VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__buf_8
XFILLER_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout698 net700 VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__buf_2
Xfanout687 _0343_ VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__buf_2
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1180_ net436 VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG5 sky130_fd_sc_hd__inv_6
XFILLER_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2703_ net51 net744 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2634_ net49 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput235 net235 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput224 net224 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput202 net202 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput213 net213 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
X_2565_ net44 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput268 net268 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput257 net257 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput246 net246 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__buf_8
X_1516_ _0436_ _0439_ net645 VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__mux2_1
Xoutput279 Inst_RegFile_switch_matrix.NN4BEG0 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__buf_6
XFILLER_59_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2496_ net768 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1447_ _0374_ _0375_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR VPWR
+ _0376_ sky130_fd_sc_hd__mux2_1
XFILLER_67_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1378_ net677 _0309_ net663 _0311_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__o211a_1
XFILLER_55_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2350_ net757 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1301_ net444 _0236_ _0238_ net662 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a211o_1
X_2281_ clknet_4_11_0_UserCLK_regs _0039_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[17\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1232_ Inst_RegFile_32x4.mem\[0\]\[0\] Inst_RegFile_32x4.mem\[1\]\[0\] net615 VGND
+ VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux2_1
XFILLER_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1163_ Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q net108 VGND VGND VPWR VPWR _1055_
+ sky130_fd_sc_hd__or2_1
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1094_ Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__inv_1
XFILLER_52_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1996_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _0849_ VGND VGND VPWR VPWR _0850_
+ sky130_fd_sc_hd__and2b_1
X_2617_ net776 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_7_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2548_ net748 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_75_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2479_ net51 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload0 clknet_4_0_0_UserCLK_regs VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_8
XFILLER_7_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_10_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1850_ _0683_ _0153_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q VGND VGND VPWR VPWR
+ _0740_ sky130_fd_sc_hd__mux2_4
X_1781_ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q _0677_ Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_12_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2402_ net766 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2333_ net772 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2264_ clknet_4_7_0_UserCLK_regs _0022_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1215_ _0157_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__a21boi_2
X_2195_ net601 net461 _0957_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux2_2
X_1146_ _1033_ _1035_ _1038_ _0996_ _0994_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__a221o_2
XFILLER_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1077_ Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__inv_2
XFILLER_52_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1979_ _1029_ _0832_ _0831_ _0830_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold67 Inst_RegFile_32x4.mem\[18\]\[0\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 Inst_RegFile_32x4.mem\[8\]\[3\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 Inst_RegFile_32x4.mem\[10\]\[0\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_9 EE4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2951_ Inst_RegFile_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__buf_6
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1902_ _0782_ _0780_ Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q _0784_ _0786_ VGND
+ VGND VPWR VPWR Inst_RegFile_switch_matrix.EE4BEG2 sky130_fd_sc_hd__a32oi_1
X_2882_ FrameStrobe[10] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_60_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1833_ Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q _1072_ Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__a21oi_1
X_1764_ _0662_ _0663_ Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q VGND VGND VPWR VPWR
+ _0664_ sky130_fd_sc_hd__mux2_1
X_1695_ net92 net108 net120 net137 Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__mux4_1
X_2316_ clknet_4_11_0_UserCLK_regs _0074_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[21\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2247_ clknet_4_13_0_UserCLK_regs _0005_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[25\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2178_ net555 net606 _0954_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__mux2_4
X_1129_ Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__inv_1
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput102 S2MID[4] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput113 SS4END[3] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_2
Xinput124 W2END[6] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xinput135 W6END[1] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ net15 net128 net100 Inst_RegFile_switch_matrix.E2BEG3 Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux4_2
XFILLER_79_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2101_ net611 net502 _0934_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_65_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2032_ _0884_ _0879_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__nor2_8
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2934_ NN4END[10] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__buf_1
XFILLER_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2865_ net763 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_4
X_1816_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q net638 VGND VGND VPWR VPWR _0711_
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2796_ Inst_RegFile_switch_matrix.E2BEG0 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_6
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1747_ net58 net1 net62 net5 Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux4_1
X_1678_ _0587_ _0588_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q VGND VGND VPWR VPWR
+ _0589_ sky130_fd_sc_hd__mux2_1
XFILLER_85_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2650_ net775 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_57_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1601_ _0518_ _0519_ _0520_ net685 net644 VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__o221a_1
X_2581_ net747 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1532_ net417 _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__nand2_1
X_1463_ net99 net127 Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q VGND VGND VPWR VPWR
+ _0390_ sky130_fd_sc_hd__mux2_1
X_1394_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q _0325_ Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q
+ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_66_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2015_ net19 net104 Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q VGND VGND VPWR VPWR
+ _0869_ sky130_fd_sc_hd__mux2_1
XFILLER_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2917_ N4END[9] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_75_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2848_ net55 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_1
X_2779_ clknet_4_6_0_UserCLK_regs _0115_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold153 Inst_RegFile_32x4.mem\[19\]\[2\] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 Inst_RegFile_32x4.mem\[8\]\[1\] VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 Inst_RegFile_32x4.mem\[14\]\[1\] VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold131 Inst_RegFile_32x4.mem\[31\]\[0\] VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 Inst_RegFile_32x4.mem\[21\]\[1\] VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold175 Inst_RegFile_32x4.mem\[13\]\[3\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 Inst_RegFile_32x4.mem\[27\]\[0\] VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout611 _0896_ VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__buf_6
Xfanout622 net624 VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__clkbuf_4
Xfanout633 net635 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__buf_8
Xfanout600 _0918_ VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_84_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout655 net656 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__buf_8
Xfanout666 net669 VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__buf_12
Xfanout644 net645 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__buf_8
Xfanout688 _0343_ VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__clkbuf_4
Xfanout699 net700 VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkbuf_2
Xfanout677 net679 VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__buf_8
XFILLER_85_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2702_ net48 net744 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_30_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2633_ net758 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput225 net225 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput203 net203 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput214 net214 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__buf_2
X_2564_ net43 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput236 net236 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
Xoutput258 net258 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput247 net247 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__buf_2
X_1515_ _0437_ _0438_ net687 VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__mux2_1
Xoutput269 net269 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__buf_2
X_2495_ net37 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1446_ net87 net95 net89 net115 Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux4_1
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1377_ _0310_ net675 VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__nand2b_4
XFILLER_82_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2280_ clknet_4_14_0_UserCLK_regs _0038_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[17\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1300_ net444 _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__nor2_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1231_ net416 _0172_ net393 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1162_ _1048_ _1050_ _1053_ _0992_ _0997_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__a221o_1
X_1093_ net126 VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__inv_1
XFILLER_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1995_ _0683_ _0848_ Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q VGND VGND VPWR VPWR
+ _0849_ sky130_fd_sc_hd__mux2_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2616_ net777 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2547_ net749 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2478_ net48 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1429_ net87 net95 net113 net115 Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux4_1
XFILLER_28_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload1 clknet_4_1_0_UserCLK_regs VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1780_ net419 net649 Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q VGND VGND VPWR VPWR
+ _0678_ sky130_fd_sc_hd__mux2_1
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2401_ net767 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2332_ net773 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2263_ clknet_4_7_0_UserCLK_regs _0021_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1214_ net649 net683 net637 net447 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__mux4_2
XFILLER_65_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2194_ net629 net527 _0957_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__mux2_4
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1145_ _1033_ _1035_ _1038_ _0996_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG5
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1076_ net72 VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1978_ Inst_RegFile_switch_matrix.JW2BEG7 Inst_RegFile_switch_matrix.JS2BEG7 _1028_
+ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__mux2_1
XFILLER_20_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold68 Inst_RegFile_32x4.mem\[6\]\[2\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 Inst_RegFile_32x4.mem\[24\]\[0\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2950_ Inst_RegFile_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_6
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1901_ Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q _0785_ Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__a21oi_1
X_2881_ net697 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_1
X_1832_ Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q net681 VGND VGND VPWR VPWR _0724_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_60_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1763_ net5 net90 net86 net114 Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__mux4_1
X_1694_ net64 net7 net1 net782 Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q
+ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__mux4_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2315_ clknet_4_11_0_UserCLK_regs _0073_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[21\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2246_ clknet_4_9_0_UserCLK_regs _0004_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[25\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2177_ net548 net610 _0954_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_76_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1128_ Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_11_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput103 S2MID[5] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
Xinput114 W1END[0] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_4
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput125 W2END[7] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xinput136 WW4END[0] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2100_ _0923_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__nand2_8
XFILLER_39_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2031_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q _0882_ _0883_ _0880_ _0881_ VGND
+ VGND VPWR VPWR _0885_ sky130_fd_sc_hd__a32o_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2933_ NN4END[9] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_1
X_2864_ net764 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1815_ Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q _0709_ VGND VGND VPWR VPWR _0710_
+ sky130_fd_sc_hd__nand2_1
XFILLER_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1746_ net23 net88 net86 net90 Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__mux4_1
X_1677_ net781 net93 net121 net138 Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q
+ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__mux4_1
XFILLER_85_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2229_ net605 net552 _0965_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_28_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1600_ Inst_RegFile_32x4.mem\[12\]\[2\] Inst_RegFile_32x4.mem\[13\]\[2\] net621 VGND
+ VGND VPWR VPWR _0520_ sky130_fd_sc_hd__mux2_1
X_2580_ net748 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1531_ _0454_ _0453_ net686 VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__mux2_1
X_1462_ Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q _0388_ VGND VGND VPWR VPWR _0389_
+ sky130_fd_sc_hd__or2_1
X_1393_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__inv_1
XFILLER_82_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2014_ net132 Inst_RegFile_switch_matrix.JN2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q
+ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__mux2_1
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2916_ N4END[8] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2847_ net750 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_4
X_2778_ clknet_4_7_0_UserCLK_regs _0114_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold110 Inst_RegFile_32x4.mem\[2\]\[0\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ net646 net680 net665 net427 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__mux4_1
Xhold143 Inst_RegFile_32x4.mem\[7\]\[3\] VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 Inst_RegFile_32x4.mem\[2\]\[2\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 Inst_RegFile_32x4.mem\[1\]\[0\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 Inst_RegFile_32x4.mem\[13\]\[0\] VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 Inst_RegFile_32x4.mem\[13\]\[2\] VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 Inst_RegFile_32x4.mem\[29\]\[0\] VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 Inst_RegFile_32x4.mem\[15\]\[2\] VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 A_ADR0 VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__buf_8
Xfanout623 net624 VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkbuf_2
Xfanout601 _0918_ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__clkbuf_2
Xfanout667 net668 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__buf_2
Xfanout656 AD2 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__buf_8
Xfanout634 net635 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__buf_8
Xfanout645 _0368_ VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__buf_6
Xfanout678 net679 VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__buf_4
Xfanout689 _0324_ VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__buf_4
XFILLER_73_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2701_ net769 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_30_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2632_ net759 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput226 net226 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput204 net204 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput215 net215 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
X_2563_ net765 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput237 net237 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
Xoutput259 net259 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput248 net248 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_8
X_1514_ Inst_RegFile_32x4.mem\[30\]\[1\] Inst_RegFile_32x4.mem\[31\]\[1\] net624 VGND
+ VGND VPWR VPWR _0438_ sky130_fd_sc_hd__mux2_1
XFILLER_4_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2494_ net771 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1445_ net59 net67 net2 net10 Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux4_1
XFILLER_4_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1376_ Inst_RegFile_32x4.mem\[12\]\[3\] Inst_RegFile_32x4.mem\[13\]\[3\] net395 VGND
+ VGND VPWR VPWR _0310_ sky130_fd_sc_hd__mux2_4
XFILLER_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1230_ _0171_ _0170_ net445 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
XFILLER_49_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1161_ _1050_ _1048_ _1053_ _0992_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG3
+ sky130_fd_sc_hd__a22o_4
XFILLER_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1092_ net13 VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__inv_2
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1994_ net75 net18 net103 net131 Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q
+ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__mux4_2
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2615_ net778 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2546_ net751 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2477_ net38 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1428_ net59 net67 net2 net10 Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux4_1
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1359_ Inst_RegFile_32x4.mem\[30\]\[3\] Inst_RegFile_32x4.mem\[31\]\[3\] net619 VGND
+ VGND VPWR VPWR _0293_ sky130_fd_sc_hd__mux2_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3029_ WW4END[4] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__buf_2
XFILLER_70_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload2 clknet_4_2_0_UserCLK_regs VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_59_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2400_ net768 net742 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2331_ net774 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2262_ clknet_4_3_0_UserCLK_regs _0020_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1213_ Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q _0155_ VGND VGND VPWR VPWR _0156_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2193_ net605 net515 _0957_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__mux2_4
X_1144_ _1036_ _1037_ _0995_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__mux2_1
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1075_ Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__inv_1
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1977_ _1028_ _0726_ Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q VGND VGND VPWR VPWR
+ _0831_ sky130_fd_sc_hd__a21oi_1
X_2529_ net767 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_3_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold69 Inst_RegFile_32x4.mem\[3\]\[3\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1900_ net86 net405 Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _0785_ sky130_fd_sc_hd__mux2_1
X_2880_ net701 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_2
X_1831_ net418 net2 net115 net414 Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q
+ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_60_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1762_ net58 net62 net82 net1 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__mux4_1
X_1693_ _1011_ _0601_ Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q VGND VGND VPWR VPWR
+ _0602_ sky130_fd_sc_hd__o21a_1
X_2314_ clknet_4_10_0_UserCLK_regs _0072_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[21\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2245_ clknet_4_15_0_UserCLK_regs _0003_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[24\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2176_ _0942_ _0927_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__nor2_8
X_1127_ Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__inv_1
XFILLER_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput104 S2MID[6] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput126 W2MID[0] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xinput115 W1END[1] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
Xinput137 WW4END[1] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_2
XFILLER_48_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2030_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q _0882_ _0883_ _0880_ _0881_ VGND
+ VGND VPWR VPWR _0884_ sky130_fd_sc_hd__a32oi_4
XFILLER_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2932_ NN4END[8] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__buf_1
X_2863_ net765 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_1
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1814_ net689 _0708_ Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q VGND VGND VPWR VPWR
+ _0709_ sky130_fd_sc_hd__mux2_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1745_ _1017_ _0644_ Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q VGND VGND VPWR VPWR
+ _0647_ sky130_fd_sc_hd__o21a_1
XFILLER_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1676_ net65 net2 net81 net8 Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q
+ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__mux4_1
XFILLER_85_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2228_ net608 net470 _0965_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_28_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2159_ net466 net631 _0950_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux2_4
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1530_ Inst_RegFile_32x4.mem\[12\]\[1\] Inst_RegFile_32x4.mem\[13\]\[1\] net621 VGND
+ VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux2_1
XFILLER_4_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1461_ net71 net14 Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q VGND VGND VPWR VPWR
+ _0388_ sky130_fd_sc_hd__mux2_1
X_1392_ net73 net16 net101 net129 Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q
+ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux4_1
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2013_ _0778_ _0866_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q VGND VGND VPWR VPWR
+ _0867_ sky130_fd_sc_hd__mux2_4
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2915_ N4END[7] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2846_ net54 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__buf_4
Xhold100 Inst_RegFile_32x4.mem\[7\]\[0\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
X_2777_ clknet_4_7_0_UserCLK_regs _0113_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold144 Inst_RegFile_32x4.mem\[24\]\[3\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold133 Inst_RegFile_32x4.mem\[6\]\[0\] VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ net693 net414 net415 net407 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux4_2
Xhold122 Inst_RegFile_32x4.mem\[14\]\[3\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 Inst_RegFile_32x4.mem\[3\]\[0\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 Inst_RegFile_32x4.mem\[19\]\[3\] VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 Inst_RegFile_32x4.mem\[11\]\[1\] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 Inst_RegFile_32x4.mem\[15\]\[1\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ net681 net634 net665 net639 Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q
+ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__mux4_2
Xfanout624 net625 VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__clkbuf_4
Xfanout602 net603 VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__clkbuf_2
Xfanout646 net647 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__buf_4
Xfanout657 net661 VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__buf_8
Xfanout635 BD2 VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__buf_8
Xfanout668 net669 VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__buf_2
Xfanout679 _1062_ VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__buf_6
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2700_ net780 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_30_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2631_ net760 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput205 net205 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput216 net216 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__buf_2
X_2562_ net766 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput238 net238 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput249 net249 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__buf_4
Xoutput227 net227 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
X_1513_ Inst_RegFile_32x4.mem\[28\]\[1\] Inst_RegFile_32x4.mem\[29\]\[1\] net624 VGND
+ VGND VPWR VPWR _0437_ sky130_fd_sc_hd__mux2_1
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2493_ net35 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1444_ _0371_ _0372_ Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR VPWR
+ _0373_ sky130_fd_sc_hd__mux2_4
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1375_ Inst_RegFile_32x4.mem\[14\]\[3\] Inst_RegFile_32x4.mem\[15\]\[3\] net395 VGND
+ VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_2
XFILLER_67_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2829_ EE4END[9] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_1
XFILLER_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1160_ _1051_ _1052_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q VGND VGND VPWR VPWR
+ _1053_ sky130_fd_sc_hd__mux2_1
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1091_ Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__inv_2
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1993_ _0838_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__and2b_2
X_2614_ net779 net720 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2545_ net752 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2476_ net27 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1427_ _0355_ _0356_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q VGND VGND VPWR VPWR
+ _0357_ sky130_fd_sc_hd__mux2_4
X_1358_ _0290_ _0291_ net678 VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__mux2_1
XFILLER_55_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1289_ Inst_RegFile_32x4.mem\[8\]\[1\] Inst_RegFile_32x4.mem\[9\]\[1\] net614 VGND
+ VGND VPWR VPWR _0227_ sky130_fd_sc_hd__mux2_1
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload3 clknet_4_3_0_UserCLK_regs VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_6
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2330_ net775 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2261_ clknet_4_3_0_UserCLK_regs _0019_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[28\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1212_ net138 net673 net659 net413 Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux4_1
XFILLER_77_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2192_ net609 net503 _0957_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__mux2_2
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1143_ net60 net68 net784 net11 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__mux4_1
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1074_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__inv_1
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1976_ _0661_ _0665_ _1028_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__a21o_1
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2528_ net768 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2459_ net774 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_3_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1830_ _0718_ _0721_ Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q _0722_ VGND VGND VPWR
+ VPWR Inst_RegFile_switch_matrix.WW4BEG0 sky130_fd_sc_hd__o22a_1
X_1761_ Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q _0660_ VGND VGND VPWR VPWR _0661_
+ sky130_fd_sc_hd__nand2_4
X_1692_ net680 net427 net665 net638 Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q
+ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__mux4_2
X_2313_ clknet_4_11_0_UserCLK_regs _0071_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[20\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ clknet_4_13_0_UserCLK_regs _0002_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[24\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2175_ net566 net603 _0953_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__mux2_4
XFILLER_65_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1126_ Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__inv_1
XFILLER_53_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1959_ net781 net107 net92 net671 Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S4BEG0 sky130_fd_sc_hd__mux4_1
Xinput105 S2MID[7] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xinput116 W1END[2] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput127 W2MID[1] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xinput138 WW4END[2] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2931_ NN4END[7] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_73_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2862_ net41 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
X_2793_ Inst_RegFile_switch_matrix.E1BEG1 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_6
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1813_ net66 net9 net112 net122 Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q
+ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__mux4_2
X_1744_ Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q _0645_ VGND VGND VPWR VPWR _0646_
+ sky130_fd_sc_hd__or2_1
X_1675_ _0585_ _1007_ Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q VGND VGND VPWR VPWR
+ _0586_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2227_ _0923_ _0937_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_28_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2158_ net463 net606 _0950_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__mux2_4
X_1109_ net98 VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2089_ net550 net631 _0928_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__mux2_4
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1460_ net70 net13 net126 Inst_RegFile_switch_matrix.JW2BEG6 Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__mux4_2
X_1391_ _0201_ _0202_ _0203_ _0975_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q VGND
+ VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_78_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2012_ net8 net113 net138 Inst_RegFile_switch_matrix.JN2BEG2 Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_35_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2914_ N4END[6] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
X_2845_ net53 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
X_2776_ clknet_4_6_0_UserCLK_regs _0112_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold101 Inst_RegFile_32x4.mem\[30\]\[3\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1727_ _0631_ _0628_ Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JW2BEG0 sky130_fd_sc_hd__mux2_4
Xhold112 Inst_RegFile_32x4.mem\[5\]\[0\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 Inst_RegFile_32x4.mem\[9\]\[3\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 Inst_RegFile_32x4.mem\[3\]\[1\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 Inst_RegFile_32x4.mem\[21\]\[0\] VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 Inst_RegFile_32x4.mem\[19\]\[0\] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 Inst_RegFile_32x4.mem\[30\]\[0\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ net690 net670 net661 net647 Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__mux4_1
Xfanout614 net616 VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__clkbuf_4
Xhold178 Inst_RegFile_32x4.mem\[11\]\[3\] VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _0918_ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout636 net637 VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__buf_8
Xfanout658 net660 VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__buf_6
X_1589_ Inst_RegFile_32x4.mem\[20\]\[2\] Inst_RegFile_32x4.mem\[21\]\[2\] net626 VGND
+ VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux2_1
Xfanout647 AD3 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__buf_2
Xfanout625 B_ADR0 VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__buf_6
Xfanout669 BD1 VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__buf_8
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2630_ net761 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_40_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput206 net206 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput217 net217 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__buf_2
X_2561_ net767 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput228 net228 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput239 net239 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
X_1512_ _0435_ _0434_ net688 VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__mux2_1
X_2492_ net34 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1443_ net648 net636 net667 net641 Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__mux4_2
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1374_ net663 _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__and2b_1
XFILLER_82_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2828_ EE4END[8] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_1
X_2759_ clknet_4_2_0_UserCLK_regs _0095_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1090_ net139 VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__inv_1
XFILLER_64_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1992_ _0845_ _0843_ Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q VGND VGND VPWR VPWR
+ _0846_ sky130_fd_sc_hd__mux2_4
XFILLER_9_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload10 clknet_4_11_0_UserCLK_regs VGND VGND VPWR VPWR clkload10/X sky130_fd_sc_hd__clkbuf_8
X_2613_ net747 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2544_ net753 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2475_ net755 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1426_ net648 net428 net431 net641 Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q
+ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux4_2
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1357_ Inst_RegFile_32x4.mem\[24\]\[3\] Inst_RegFile_32x4.mem\[25\]\[3\] net619 VGND
+ VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
XFILLER_83_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1288_ Inst_RegFile_32x4.mem\[10\]\[1\] Inst_RegFile_32x4.mem\[11\]\[1\] net614 VGND
+ VGND VPWR VPWR _0226_ sky130_fd_sc_hd__mux2_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload4 clknet_4_4_0_UserCLK_regs VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__clkinv_2
XFILLER_3_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2260_ clknet_4_12_0_UserCLK_regs _0018_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[28\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1211_ _0153_ _0152_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q VGND VGND VPWR VPWR
+ _0154_ sky130_fd_sc_hd__mux2_4
XFILLER_49_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2191_ _0926_ _0933_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__nand2_4
X_1142_ net25 net86 net88 net96 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__mux4_1
XFILLER_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1975_ net407 Inst_RegFile_switch_matrix.JW2BEG3 _0829_ _0828_ Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N1BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2527_ net770 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2458_ net775 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1409_ _0335_ Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q _0336_ _0339_ VGND VGND
+ VPWR VPWR _0340_ sky130_fd_sc_hd__a31o_1
XFILLER_68_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2389_ net56 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1760_ _0658_ _0659_ Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q VGND VGND VPWR VPWR
+ _0660_ sky130_fd_sc_hd__mux2_4
X_1691_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q _0599_ VGND VGND VPWR VPWR _0600_
+ sky130_fd_sc_hd__or2_1
X_2312_ clknet_4_11_0_UserCLK_regs _0070_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[20\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ clknet_4_13_0_UserCLK_regs _0001_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[24\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2174_ net561 net631 _0953_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_4
XFILLER_65_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1125_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_76_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1958_ net782 net93 net108 net661 Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S4BEG1 sky130_fd_sc_hd__mux4_1
X_1889_ net68 net11 net113 net124 Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q
+ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__mux4_1
Xclkbuf_4_9_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_9_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
Xinput106 S4END[0] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_4
Xinput117 W1END[3] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_2
Xinput128 W2MID[2] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_2
Xinput139 WW4END[3] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_4
XFILLER_56_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_90 net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2930_ NN4END[6] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2861_ net767 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_1
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1812_ _0705_ _0707_ Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.WW4BEG3 sky130_fd_sc_hd__mux2_4
X_1743_ net114 net672 net658 net419 Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__mux4_1
X_1674_ net684 net636 net668 net642 Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q
+ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__mux4_2
XFILLER_85_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2226_ net601 net486 _0964_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__mux2_4
XFILLER_26_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2157_ net459 net610 _0950_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__mux2_4
XFILLER_38_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1108_ Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__inv_1
X_2088_ net539 net606 _0928_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__mux2_4
XFILLER_53_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1390_ Inst_RegFile_32x4.AD_comb\[3\] Inst_RegFile_32x4.AD_reg\[3\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ VGND VGND VPWR VPWR AD3 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_78_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2011_ Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q _0859_ _0862_ _0864_ VGND VGND VPWR
+ VPWR _0865_ sky130_fd_sc_hd__a22o_1
XFILLER_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2913_ N4END[5] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2844_ net52 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_2
X_2775_ clknet_4_5_0_UserCLK_regs _0111_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1726_ _0629_ _0630_ Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR VPWR
+ _0631_ sky130_fd_sc_hd__mux2_1
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold124 Inst_RegFile_32x4.mem\[15\]\[0\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 Inst_RegFile_32x4.mem\[9\]\[2\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 Inst_RegFile_32x4.mem\[3\]\[2\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 Inst_RegFile_32x4.mem\[5\]\[3\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 Inst_RegFile_32x4.mem\[17\]\[0\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 Inst_RegFile_32x4.mem\[9\]\[1\] VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 Inst_RegFile_32x4.mem\[6\]\[1\] VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _0570_ _0567_ Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JW2BEG2 sky130_fd_sc_hd__mux2_4
X_1588_ _0506_ _0507_ net688 VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__mux2_1
Xhold179 Inst_RegFile_32x4.mem\[25\]\[3\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout615 net616 VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__clkbuf_4
Xfanout604 _0900_ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__buf_2
Xfanout648 net650 VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__buf_8
Xfanout637 BD2 VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__buf_8
Xfanout626 B_ADR0 VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__clkbuf_4
Xfanout659 net660 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__buf_4
XFILLER_85_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2209_ net604 net538 _0961_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_84_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput207 net207 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__buf_2
X_2560_ net768 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput229 net229 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput218 net218 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
X_2491_ net774 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1511_ Inst_RegFile_32x4.mem\[24\]\[1\] Inst_RegFile_32x4.mem\[25\]\[1\] net628 VGND
+ VGND VPWR VPWR _0435_ sky130_fd_sc_hd__mux2_1
X_1442_ net139 net672 net658 net654 Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux4_1
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1373_ _0305_ _0306_ net676 VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__mux2_1
XFILLER_67_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3043_ Inst_RegFile_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_2
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2827_ EE4END[7] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_1
X_2758_ clknet_4_0_0_UserCLK_regs _0094_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1709_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q _0615_ Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__o21a_1
X_2689_ net767 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1991_ _0829_ _0844_ _1027_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__mux2_4
XFILLER_9_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2612_ net748 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
Xclkload11 clknet_4_12_0_UserCLK_regs VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__bufinv_16
X_2543_ net51 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_81_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2474_ net756 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1425_ net692 net672 net658 net654 Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux4_1
X_1356_ Inst_RegFile_32x4.mem\[26\]\[3\] Inst_RegFile_32x4.mem\[27\]\[3\] net619 VGND
+ VGND VPWR VPWR _0290_ sky130_fd_sc_hd__mux2_1
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1287_ Inst_RegFile_32x4.AD_comb\[0\] Inst_RegFile_32x4.AD_reg\[0\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ VGND VGND VPWR VPWR AD0 sky130_fd_sc_hd__mux2_4
X_3026_ W6END[11] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload5 clknet_4_5_0_UserCLK_regs VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1210_ net84 net6 net91 net119 Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q
+ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__mux4_2
X_2190_ net531 net602 _0956_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__mux2_2
X_1141_ Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q _1034_ Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__o21a_1
XFILLER_80_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ net646 _0563_ Inst_RegFile_switch_matrix.JW2BEG0 net396 Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N1BEG1
+ sky130_fd_sc_hd__mux4_2
X_2526_ net771 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2457_ net776 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1408_ Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q _0338_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q
+ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2388_ net55 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1339_ Inst_RegFile_32x4.mem\[26\]\[2\] Inst_RegFile_32x4.mem\[27\]\[2\] net619 VGND
+ VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
XFILLER_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3009_ net126 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_54_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput390 net390 VGND VGND VPWR VPWR WW4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_59_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1690_ net691 net670 net407 net646 Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__mux4_1
X_2311_ clknet_4_11_0_UserCLK_regs _0069_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[20\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ clknet_4_8_0_UserCLK_regs _0000_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[24\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2173_ net578 net607 _0953_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_4
X_1124_ Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_76_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1957_ net90 net690 net109 net653 Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_2
X_1888_ Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q net434 _0773_ Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q
+ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__a211oi_1
X_2509_ net769 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput107 S4END[1] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
Xinput118 W2END[0] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput129 W2MID[3] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_2
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_80 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _0325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2860_ net39 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_1
X_1811_ net683 _1073_ net402 _0706_ Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__mux4_2
X_2791_ clknet_4_3_0_UserCLK_regs _0127_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1742_ net648 net683 net431 net637 Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q
+ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__mux4_1
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1673_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q _0583_ VGND VGND VPWR VPWR _0584_
+ sky130_fd_sc_hd__or2_1
X_2225_ net629 net498 _0964_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__mux2_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2156_ _0942_ _0924_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__nor2_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__inv_1
XFILLER_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2087_ net556 net610 _0928_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_36_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2989_ SS4END[13] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2010_ _1031_ _0863_ Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q VGND VGND VPWR VPWR
+ _0864_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2912_ N4END[4] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2843_ net754 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
X_2774_ clknet_4_5_0_UserCLK_regs _0110_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1725_ net91 net107 net110 net119 Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__mux4_1
Xhold125 Inst_RegFile_32x4.mem\[1\]\[2\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 Inst_RegFile_32x4.mem\[30\]\[1\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 Inst_RegFile_32x4.mem\[20\]\[3\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 Inst_RegFile_32x4.mem\[17\]\[1\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 Inst_RegFile_32x4.mem\[27\]\[1\] VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 Inst_RegFile_32x4.mem\[27\]\[2\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ _0568_ _0569_ Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR VPWR
+ _0570_ sky130_fd_sc_hd__mux2_1
Xhold169 Inst_RegFile_32x4.mem\[21\]\[2\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ Inst_RegFile_32x4.mem\[18\]\[2\] Inst_RegFile_32x4.mem\[19\]\[2\] net627 VGND
+ VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux2_1
Xfanout605 _0900_ VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout649 net650 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__buf_8
Xfanout627 net628 VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__clkbuf_2
Xfanout638 net640 VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__buf_6
Xfanout616 A_ADR0 VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__buf_2
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2208_ net608 net525 _0961_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_84_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ net577 net632 _0946_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__mux2_4
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput208 net208 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput219 net219 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
X_2490_ net775 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1510_ Inst_RegFile_32x4.mem\[26\]\[1\] Inst_RegFile_32x4.mem\[27\]\[1\] net628 VGND
+ VGND VPWR VPWR _0434_ sky130_fd_sc_hd__mux2_1
XFILLER_57_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1441_ _0369_ _0344_ net688 VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux2_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1372_ Inst_RegFile_32x4.mem\[8\]\[3\] Inst_RegFile_32x4.mem\[9\]\[3\] net614 VGND
+ VGND VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
XFILLER_67_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2826_ EE4END[6] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_1
X_2757_ clknet_4_0_0_UserCLK_regs _0093_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2688_ net768 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1708_ net691 net670 net652 net646 Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__mux4_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1639_ _0553_ _0554_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q VGND VGND VPWR VPWR
+ _0555_ sky130_fd_sc_hd__mux2_4
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1990_ net70 net126 net98 Inst_RegFile_switch_matrix.JW2BEG4 Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_43_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2611_ net749 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
Xclkload12 clknet_4_14_0_UserCLK_regs VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinv_4
X_2542_ net48 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2473_ net758 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1424_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q _0205_ Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q
+ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__a21o_1
X_1355_ Inst_RegFile_32x4.AD_comb\[2\] Inst_RegFile_32x4.AD_reg\[2\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ VGND VGND VPWR VPWR AD2 sky130_fd_sc_hd__mux2_4
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3025_ W6END[10] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_2
X_1286_ _0182_ _0210_ _0209_ _0225_ VGND VGND VPWR VPWR Inst_RegFile_32x4.AD_comb\[0\]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_70_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload6 clknet_4_6_0_UserCLK_regs VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinv_2
X_2809_ net18 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1140_ net116 net674 net660 net413 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__mux4_1
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1973_ net680 net689 Inst_RegFile_switch_matrix.JW2BEG1 _0377_ Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N1BEG2
+ sky130_fd_sc_hd__mux4_2
X_2525_ net772 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2456_ net777 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1407_ _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__inv_2
X_2387_ net750 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1338_ _0266_ _0273_ net651 VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_4
XFILLER_83_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1269_ _0208_ _0193_ Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q VGND VGND VPWR VPWR
+ _0209_ sky130_fd_sc_hd__mux2_4
XFILLER_83_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3008_ Inst_RegFile_switch_matrix.JW2BEG7 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__buf_6
XFILLER_71_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput380 Inst_RegFile_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR WW4BEG[12] sky130_fd_sc_hd__buf_6
Xoutput391 net391 VGND VGND VPWR VPWR WW4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_86_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2310_ clknet_4_10_0_UserCLK_regs _0068_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[20\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2241_ net600 net496 _0967_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_68_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2172_ net537 net610 _0953_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_4
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1123_ Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__inv_2
XFILLER_65_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1956_ net91 net691 net106 net647 Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
X_1887_ Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q net684 VGND VGND VPWR VPWR _0773_
+ sky130_fd_sc_hd__nor2_1
X_2508_ net780 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput108 S4END[2] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
X_2439_ net760 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput119 W2END[1] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_2
XFILLER_56_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_70 NN4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 net359 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_92 _0697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1810_ net66 net94 net23 net122 Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q
+ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__mux4_2
X_2790_ clknet_4_1_0_UserCLK_regs _0126_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1741_ _0643_ _0640_ Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JS2BEG0 sky130_fd_sc_hd__mux2_4
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1672_ net690 net673 net658 net649 Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q
+ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__mux4_1
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2224_ net605 net520 _0964_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_4
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2155_ net554 net602 _0949_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__mux2_4
X_1106_ Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__inv_2
XFILLER_53_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2086_ _0927_ _0855_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__nor2_8
X_2988_ SS4END[12] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_2
X_1939_ _0683_ _1060_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q VGND VGND VPWR VPWR
+ _0819_ sky130_fd_sc_hd__mux2_2
Xinput90 S2END[0] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_5_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_5_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2911_ net77 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2842_ net757 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
X_2773_ clknet_4_5_0_UserCLK_regs _0109_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1724_ net61 net63 net6 net781 Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__mux4_1
Xhold104 Inst_RegFile_32x4.mem\[12\]\[3\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 Inst_RegFile_32x4.mem\[1\]\[1\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 Inst_RegFile_32x4.mem\[24\]\[1\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 Inst_RegFile_32x4.mem\[15\]\[3\] VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 Inst_RegFile_32x4.mem\[29\]\[2\] VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 Inst_RegFile_32x4.mem\[25\]\[1\] VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ net22 net93 net109 net121 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__mux4_1
X_1586_ Inst_RegFile_32x4.mem\[16\]\[2\] Inst_RegFile_32x4.mem\[17\]\[2\] net626 VGND
+ VGND VPWR VPWR _0506_ sky130_fd_sc_hd__mux2_1
Xfanout606 net607 VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_13_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout639 net640 VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_4
Xfanout617 A_ADR0 VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__clkbuf_4
Xfanout628 B_ADR0 VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__clkbuf_4
X_2207_ _0923_ net439 VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__nand2_8
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2138_ net511 net607 _0946_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__mux2_2
XFILLER_81_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2069_ _0865_ _0878_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__nand2b_1
XFILLER_41_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput209 net209 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
X_1440_ Inst_RegFile_32x4.mem\[24\]\[0\] Inst_RegFile_32x4.mem\[25\]\[0\] net628 VGND
+ VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux2_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1371_ Inst_RegFile_32x4.mem\[10\]\[3\] Inst_RegFile_32x4.mem\[11\]\[3\] net616 VGND
+ VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2825_ EE4END[5] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_1
X_2756_ clknet_4_0_0_UserCLK_regs _0092_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2687_ net770 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1707_ _1015_ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__or2_4
X_1638_ net681 net634 net665 net639 Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q
+ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__mux4_2
X_1569_ Inst_RegFile_32x4.mem\[0\]\[3\] Inst_RegFile_32x4.mem\[1\]\[3\] net625 VGND
+ VGND VPWR VPWR _0491_ sky130_fd_sc_hd__mux2_1
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2610_ net54 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
Xclkload13 clknet_4_15_0_UserCLK_regs VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinv_2
X_2541_ net769 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2472_ net46 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1423_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q _0352_ VGND VGND VPWR VPWR _0353_
+ sky130_fd_sc_hd__and2b_1
X_1354_ _0274_ _0289_ _0209_ VGND VGND VPWR VPWR Inst_RegFile_32x4.AD_comb\[2\] sky130_fd_sc_hd__mux2_4
XFILLER_83_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1285_ _0217_ _0224_ _0169_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__mux2_1
XFILLER_83_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3024_ W6END[9] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_2
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload7 clknet_4_8_0_UserCLK_regs VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinv_4
X_2808_ net17 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
X_2739_ clknet_4_8_0_UserCLK_regs Inst_RegFile_32x4.AD_comb\[3\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.AD_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1972_ net667 _0407_ Inst_RegFile_switch_matrix.JW2BEG2 _0827_ Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q
+ Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N1BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_81_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2524_ net34 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2455_ net778 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2386_ net54 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1406_ net80 net112 Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR
+ _0337_ sky130_fd_sc_hd__mux2_1
XFILLER_68_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1337_ _0269_ _0272_ net662 VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__mux2_4
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1268_ _0206_ _0207_ _1006_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1199_ Inst_RegFile_32x4.mem\[10\]\[0\] Inst_RegFile_32x4.mem\[11\]\[0\] net616 VGND
+ VGND VPWR VPWR _0143_ sky130_fd_sc_hd__mux2_1
X_3007_ Inst_RegFile_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__buf_1
XFILLER_36_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput370 net370 VGND VGND VPWR VPWR W6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput392 net392 VGND VGND VPWR VPWR WW4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput381 Inst_RegFile_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR WW4BEG[13] sky130_fd_sc_hd__buf_8
XFILLER_59_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2240_ net630 net454 _0967_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__mux2_2
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2171_ _0944_ _0921_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__nor2_8
XFILLER_76_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1122_ Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__inv_1
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1955_ net406 Inst_RegFile_switch_matrix.JS2BEG3 _0829_ _0828_ Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.W1BEG0
+ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_78_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1886_ net418 net2 net87 net674 Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q
+ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__mux4_1
X_2507_ net755 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput109 S4END[3] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
X_2438_ net762 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2369_ net767 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_13_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_13_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_71 NN4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_60 N4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_93 _0697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1740_ _0642_ _0641_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q VGND VGND VPWR VPWR
+ _0643_ sky130_fd_sc_hd__mux2_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1671_ _0582_ _0579_ Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.E2BEG2 sky130_fd_sc_hd__mux2_4
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2223_ net609 net476 _0964_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__mux2_4
XFILLER_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2154_ net474 net631 _0949_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__mux2_4
X_1105_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_64_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2085_ _0885_ _0919_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__or2_4
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2987_ SS4END[11] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_2
X_1938_ _0681_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q
+ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__a21oi_2
X_1869_ net684 net398 net668 net404 Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__mux4_1
Xinput91 S2END[1] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_4
Xinput80 N4END[2] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2910_ net76 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2841_ net38 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2772_ clknet_4_4_0_UserCLK_regs _0108_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1723_ _0626_ _0627_ Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q VGND VGND VPWR VPWR
+ _0628_ sky130_fd_sc_hd__mux2_4
Xhold105 Inst_RegFile_32x4.mem\[5\]\[2\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold116 Inst_RegFile_32x4.mem\[11\]\[2\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 Inst_RegFile_32x4.mem\[22\]\[0\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 Inst_RegFile_32x4.mem\[1\]\[3\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ net59 net65 net84 net8 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__mux4_1
Xhold149 Inst_RegFile_32x4.mem\[22\]\[3\] VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
X_1585_ _0501_ _0504_ net644 VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux2_1
Xfanout629 net630 VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_2
Xfanout618 net619 VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__clkbuf_2
Xfanout607 _0900_ VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2206_ net600 net505 _0960_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__mux2_4
XFILLER_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2137_ net573 net611 _0946_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux2_4
XFILLER_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2068_ net536 net602 _0888_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__mux2_4
XFILLER_81_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1370_ _0296_ _0303_ net651 VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_1
XFILLER_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3040_ WW4END[15] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__buf_2
XFILLER_84_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2824_ EE4END[4] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_1
X_2755_ clknet_4_6_0_UserCLK_regs _0091_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2686_ net771 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1706_ net680 net633 net665 net638 Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q
+ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__mux4_2
X_1637_ net691 net670 net657 net653 Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__mux4_2
XFILLER_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1568_ _0486_ _0489_ net643 VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux2_2
XFILLER_48_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1499_ Inst_RegFile_32x4.mem\[2\]\[0\] Inst_RegFile_32x4.mem\[3\]\[0\] net625 VGND
+ VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux2_1
XFILLER_58_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2540_ net27 net714 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2471_ net760 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1422_ net17 net102 net130 Inst_RegFile_switch_matrix.JS2BEG6 Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__mux4_2
XFILLER_68_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1353_ _0281_ _0288_ net393 VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__mux2_4
X_1284_ _0220_ _0223_ net664 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3023_ W6END[8] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload8 clknet_4_9_0_UserCLK_regs VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__clkinv_4
X_2807_ net16 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
X_2738_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.AD_comb\[2\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.AD_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_2669_ net769 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1971_ net64 net79 net781 net681 Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N4BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_60_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2523_ net33 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2454_ net28 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2385_ net53 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1405_ Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q net120 VGND VGND VPWR VPWR _0336_
+ sky130_fd_sc_hd__or2_1
XFILLER_68_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1336_ _0270_ _0271_ net675 VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_3_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 E1END[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_83_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1267_ net63 net91 Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q VGND VGND VPWR VPWR
+ _0207_ sky130_fd_sc_hd__mux2_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1198_ _0130_ _0141_ Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q VGND VGND VPWR VPWR
+ _0142_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_54_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput360 net360 VGND VGND VPWR VPWR W2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput371 net371 VGND VGND VPWR VPWR W6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput382 net382 VGND VGND VPWR VPWR WW4BEG[14] sky130_fd_sc_hd__buf_6
XFILLER_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2170_ net495 net603 _0952_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__mux2_4
X_1121_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_76_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1954_ net71 net14 net99 net127 Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q
+ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__mux4_2
X_1885_ _0765_ _0771_ Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.E6BEG0 sky130_fd_sc_hd__mux2_1
X_2506_ net756 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2437_ net763 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2368_ net768 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2299_ clknet_4_14_0_UserCLK_regs _0057_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[16\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1319_ _0255_ _0256_ net678 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_50 net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 NN4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 N4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 net693 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput190 net190 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__buf_2
XFILLER_47_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK VGND VGND VPWR VPWR clknet_1_0__leaf_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1670_ _0580_ _0581_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR VPWR
+ _0582_ sky130_fd_sc_hd__mux2_1
XFILLER_78_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2222_ _0933_ _0886_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__nand2_8
XFILLER_38_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2153_ net487 net606 _0949_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_64_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1104_ net74 VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__inv_2
X_2084_ _0885_ _0919_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__nor2_2
XFILLER_34_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2986_ SS4END[10] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_2
X_1937_ Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q net398 VGND VGND VPWR VPWR _0817_
+ sky130_fd_sc_hd__or2_1
X_1868_ _0682_ _0683_ _1073_ net402 Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__mux4_2
Xinput81 N4END[3] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
Xinput70 N2MID[0] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
Xinput92 S2END[2] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_4
X_1799_ _0693_ _0694_ _0695_ Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q VGND VGND
+ VPWR VPWR _0696_ sky130_fd_sc_hd__o22a_1
XFILLER_67_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2840_ net27 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_1
X_2771_ clknet_4_2_0_UserCLK_regs _0107_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1722_ net680 net633 net665 net638 Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__mux4_2
Xhold117 Inst_RegFile_32x4.mem\[7\]\[1\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 Inst_RegFile_32x4.mem\[0\]\[2\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
X_1653_ _0565_ _0566_ Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR VPWR
+ _0567_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold128 Inst_RegFile_32x4.mem\[0\]\[1\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 Inst_RegFile_32x4.mem\[31\]\[3\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
X_1584_ _0502_ _0503_ net687 VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__mux2_1
Xfanout608 net609 VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__buf_4
Xfanout619 A_ADR0 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__clkbuf_4
X_2205_ net630 net497 _0960_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux2_4
XFILLER_81_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2136_ _0927_ _0944_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__nor2_8
XFILLER_81_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2067_ _1024_ _0912_ _0917_ _0908_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__a31o_2
XFILLER_81_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2969_ S4END[9] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__buf_2
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone40 net625 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_1_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_1_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_48_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2754_ clknet_4_7_0_UserCLK_regs _0090_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1705_ _0609_ _0607_ _0612_ _1014_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG1
+ sky130_fd_sc_hd__a22o_4
X_2685_ net772 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1636_ _0542_ Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q _0546_ _0552_ VGND VGND
+ VPWR VPWR B_ADR0 sky130_fd_sc_hd__a22o_4
X_1567_ _0487_ _0488_ net686 VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__mux2_1
X_1498_ _0420_ _0423_ net417 VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
XFILLER_58_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2119_ net608 net568 _0940_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__mux2_4
XFILLER_39_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2470_ net761 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_55_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1421_ _0346_ _0348_ _0351_ _0982_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG6
+ sky130_fd_sc_hd__a22o_4
X_1352_ _0284_ _0287_ net664 VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_1
X_1283_ _0221_ _0222_ net678 VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__mux2_1
X_3022_ W6END[7] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_2
XFILLER_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload9 clknet_4_10_0_UserCLK_regs VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__bufinv_16
X_2806_ net15 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
X_2737_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.AD_comb\[1\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.AD_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_2668_ net780 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1619_ net418 net67 net85 net2 Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__mux4_1
X_2599_ net45 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_6_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout780 net27 VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__buf_4
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1970_ net65 net80 net782 net667 Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_60_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2522_ net32 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2453_ net747 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1404_ _0328_ _0330_ _0978_ _0333_ _0976_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__a221o_1
X_2384_ net52 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1335_ Inst_RegFile_32x4.mem\[4\]\[2\] Inst_RegFile_32x4.mem\[5\]\[2\] net612 VGND
+ VGND VPWR VPWR _0271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 E1END[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_6
XFILLER_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3005_ Inst_RegFile_switch_matrix.JW2BEG4 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_6
X_1266_ _0204_ _0205_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q VGND VGND VPWR VPWR
+ _0206_ sky130_fd_sc_hd__mux2_1
X_1197_ _0140_ _0139_ Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q VGND VGND VPWR VPWR
+ _0141_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_54_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput350 net350 VGND VGND VPWR VPWR W2BEG[1] sky130_fd_sc_hd__buf_8
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput361 net361 VGND VGND VPWR VPWR W2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput383 Inst_RegFile_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR WW4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput372 net372 VGND VGND VPWR VPWR W6BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1120_ Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__inv_1
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1953_ net80 net125 net7 Inst_RegFile_switch_matrix.E2BEG2 Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__mux4_2
X_1884_ _0768_ _0769_ _0770_ Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q VGND VGND
+ VPWR VPWR _0771_ sky130_fd_sc_hd__o22a_1
X_2505_ net47 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2436_ net764 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2367_ net770 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2298_ clknet_4_11_0_UserCLK_regs _0056_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[16\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1318_ Inst_RegFile_32x4.mem\[20\]\[1\] Inst_RegFile_32x4.mem\[21\]\[1\] net617 VGND
+ VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
X_1249_ _0190_ _0187_ Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JN2BEG5 sky130_fd_sc_hd__mux2_4
XFILLER_71_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_40 FrameStrobe[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 net259 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 NN4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_95 net693 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput191 net191 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput180 net180 VGND VGND VPWR VPWR EE4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_47_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2221_ net601 net481 _0963_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_4
XFILLER_78_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2152_ net480 net610 _0949_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__mux2_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1103_ Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__inv_2
X_2083_ net489 net602 _0925_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__mux2_4
X_2985_ SS4END[9] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_2
X_1936_ net61 net783 net692 net413 Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q
+ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__mux4_1
X_1867_ Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q _0754_ _0753_ _1022_ VGND VGND
+ VPWR VPWR _0755_ sky130_fd_sc_hd__a211o_1
Xinput82 NN4END[0] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_2
Xinput71 N2MID[1] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xinput60 N1END[2] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_4
X_1798_ net83 net4 net111 net692 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q
+ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__mux4_1
Xinput93 S2END[3] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2419_ net749 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2770_ clknet_4_0_0_UserCLK_regs _0106_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1721_ net690 net652 net657 net646 Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q
+ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__mux4_1
Xhold107 Inst_RegFile_32x4.mem\[20\]\[2\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ net683 net636 net667 net641 Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q
+ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__mux4_2
Xhold129 Inst_RegFile_32x4.mem\[4\]\[1\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 Inst_RegFile_32x4.mem\[11\]\[0\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
X_1583_ Inst_RegFile_32x4.mem\[30\]\[2\] Inst_RegFile_32x4.mem\[31\]\[2\] net624 VGND
+ VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux2_1
Xfanout609 net611 VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__buf_6
XFILLER_78_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2204_ net604 net533 _0960_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__mux2_4
X_2135_ net541 net603 _0945_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux2_4
XFILLER_81_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2066_ Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q _0915_ _0916_ VGND VGND VPWR VPWR
+ _0917_ sky130_fd_sc_hd__a21o_1
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2968_ S4END[8] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_2
X_1919_ net418 net2 net115 net673 Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q
+ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__mux4_1
X_2899_ Inst_RegFile_switch_matrix.JN2BEG3 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone52 net677 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__buf_8
XFILLER_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2822_ Inst_RegFile_switch_matrix.E6BEG0 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
X_2753_ clknet_4_7_0_UserCLK_regs _0089_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1704_ _0610_ _0611_ _1013_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__mux2_1
X_2684_ net773 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1635_ Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q _0551_ VGND VGND VPWR VPWR _0552_
+ sky130_fd_sc_hd__nor2_1
X_1566_ Inst_RegFile_32x4.mem\[14\]\[3\] Inst_RegFile_32x4.mem\[15\]\[3\] net621 VGND
+ VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux2_1
XFILLER_86_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1497_ _0421_ _0422_ net685 VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2118_ _0920_ _0939_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__nand2_8
X_2049_ net79 net690 net781 Inst_RegFile_switch_matrix.JS2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_80_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1420_ _0349_ _0350_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR VPWR
+ _0351_ sky130_fd_sc_hd__mux2_1
X_1351_ _0285_ _0286_ net679 VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
XFILLER_83_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1282_ Inst_RegFile_32x4.mem\[20\]\[0\] Inst_RegFile_32x4.mem\[21\]\[0\] net617 VGND
+ VGND VPWR VPWR _0222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3021_ W6END[6] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2805_ net14 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_1
X_2736_ clknet_4_2_0_UserCLK_regs Inst_RegFile_32x4.AD_comb\[0\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.AD_reg\[0\] sky130_fd_sc_hd__dfxtp_1
X_2667_ net755 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1618_ _0968_ _0535_ Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q VGND VGND VPWR VPWR
+ _0536_ sky130_fd_sc_hd__o21a_1
XFILLER_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2598_ net761 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1549_ _0470_ _0469_ net688 VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_1
XFILLER_59_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_regs_0_UserCLK UserCLK VGND VGND VPWR VPWR UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout770 net37 VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__clkbuf_4
Xfanout781 net22 VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__buf_2
XFILLER_18_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_130 net139 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2521_ net31 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2452_ net748 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1403_ _0334_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG4 sky130_fd_sc_hd__inv_4
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2383_ net51 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1334_ Inst_RegFile_32x4.mem\[6\]\[2\] Inst_RegFile_32x4.mem\[7\]\[2\] net612 VGND
+ VGND VPWR VPWR _0270_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1265_ net75 net18 net103 net131 Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q
+ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__mux4_1
X_3004_ Inst_RegFile_switch_matrix.JW2BEG3 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__buf_1
Xinput3 E1END[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
X_1196_ net67 net10 net111 net123 Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q
+ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_19_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2719_ net37 net744 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput340 net340 VGND VGND VPWR VPWR SS4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput351 net351 VGND VGND VPWR VPWR W2BEG[2] sky130_fd_sc_hd__buf_8
Xoutput362 net362 VGND VGND VPWR VPWR W2BEGb[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput384 net384 VGND VGND VPWR VPWR WW4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput373 net373 VGND VGND VPWR VPWR W6BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1952_ net427 _0563_ Inst_RegFile_switch_matrix.JS2BEG0 net396 Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__mux4_2
X_1883_ net684 net398 net668 net642 Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q
+ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2504_ net46 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2435_ net765 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2366_ net771 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2297_ clknet_4_6_0_UserCLK_regs _0055_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1317_ Inst_RegFile_32x4.mem\[22\]\[1\] Inst_RegFile_32x4.mem\[23\]\[1\] net617 VGND
+ VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
X_1248_ _0189_ _0188_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q VGND VGND VPWR VPWR
+ _0190_ sky130_fd_sc_hd__mux2_1
XFILLER_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _1067_ _1065_ _1070_ _1000_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__a22oi_4
XFILLER_64_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_30 net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 FrameStrobe[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 NN4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 N4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 net693 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput170 net170 VGND VGND VPWR VPWR E6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput192 net192 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput181 net181 VGND VGND VPWR VPWR EE4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2220_ net629 net467 _0963_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_4
XFILLER_78_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2151_ _0942_ _0887_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__nor2_8
X_1102_ Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__inv_2
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2082_ net472 net631 _0925_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__mux2_4
XFILLER_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2984_ SS4END[8] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_2
XFILLER_61_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1935_ Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q _0809_ _0811_ _0813_ _0815_ VGND
+ VGND VPWR VPWR Inst_RegFile_switch_matrix.NN4BEG2 sky130_fd_sc_hd__a32oi_1
X_1866_ net413 net405 Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q VGND VGND VPWR VPWR
+ _0754_ sky130_fd_sc_hd__mux2_1
Xinput50 FrameData[31] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
Xinput72 N2MID[2] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
Xinput61 N1END[3] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_4
X_1797_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0691_ Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__a21bo_1
Xinput94 S2END[4] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_2
Xinput83 NN4END[1] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_2
XFILLER_69_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2418_ net751 net696 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2349_ net769 net57 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1720_ _0625_ _0622_ Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JW2BEG7 sky130_fd_sc_hd__mux2_4
XFILLER_78_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold108 Inst_RegFile_32x4.mem\[6\]\[3\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ net135 net672 net658 net648 Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__mux4_1
Xhold119 Inst_RegFile_32x4.mem\[23\]\[1\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1582_ Inst_RegFile_32x4.mem\[28\]\[2\] Inst_RegFile_32x4.mem\[29\]\[2\] net624 VGND
+ VGND VPWR VPWR _0502_ sky130_fd_sc_hd__mux2_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2203_ net608 net504 _0960_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__mux2_4
X_2134_ net542 net632 _0945_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__mux2_4
XFILLER_81_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2065_ Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q _0914_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__o21ai_1
XFILLER_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2967_ S4END[7] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_2
X_1918_ _0798_ _0800_ _0796_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.EE4BEG0
+ sky130_fd_sc_hd__a21oi_1
X_2898_ Inst_RegFile_switch_matrix.JN2BEG2 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__buf_6
X_1849_ _0681_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q
+ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__a21oi_2
XFILLER_78_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone53 net677 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2821_ E6END[11] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2752_ clknet_4_3_0_UserCLK_regs _0088_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1703_ net58 net64 net80 net83 Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q
+ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__mux4_1
X_2683_ net774 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1634_ Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q _0548_ _0550_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q
+ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__o211a_1
X_1565_ Inst_RegFile_32x4.mem\[12\]\[3\] Inst_RegFile_32x4.mem\[13\]\[3\] net621 VGND
+ VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux2_1
X_1496_ Inst_RegFile_32x4.mem\[14\]\[0\] Inst_RegFile_32x4.mem\[15\]\[0\] net432 VGND
+ VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux2_1
XFILLER_66_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2117_ _0936_ net437 VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__nor2_8
XFILLER_81_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2048_ net507 net606 _0888_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__mux2_4
XFILLER_54_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1350_ Inst_RegFile_32x4.mem\[20\]\[2\] Inst_RegFile_32x4.mem\[21\]\[2\] net617 VGND
+ VGND VPWR VPWR _0286_ sky130_fd_sc_hd__mux2_1
X_1281_ Inst_RegFile_32x4.mem\[22\]\[0\] Inst_RegFile_32x4.mem\[23\]\[0\] net617 VGND
+ VGND VPWR VPWR _0221_ sky130_fd_sc_hd__mux2_1
XFILLER_76_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3020_ W6END[5] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2804_ net13 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2735_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.BD_comb\[3\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.BD_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_2666_ net756 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1617_ net648 net428 net667 net641 Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__mux4_2
X_2597_ net763 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1548_ Inst_RegFile_32x4.mem\[24\]\[3\] Inst_RegFile_32x4.mem\[25\]\[3\] net628 VGND
+ VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux2_1
X_1479_ _0153_ Inst_RegFile_switch_matrix.JS2BEG6 Inst_RegFile_switch_matrix.JN2BEG6
+ Inst_RegFile_switch_matrix.JW2BEG6 Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q
+ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux4_1
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_UserCLK_regs UserCLK_regs VGND VGND VPWR VPWR clknet_0_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout760 net45 VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__buf_4
Xfanout782 net21 VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__clkbuf_4
Xfanout771 net36 VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_120 net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_131 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2520_ net30 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2451_ net750 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1402_ _0330_ _0328_ _0333_ _0978_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a22oi_4
X_2382_ net48 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1333_ _0267_ _0268_ net676 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_3_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1264_ _0201_ _0202_ _0203_ _0975_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__a22o_1
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3003_ Inst_RegFile_switch_matrix.JW2BEG2 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__buf_6
Xinput4 E1END[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_1195_ net79 net122 net111 Inst_RegFile_switch_matrix.JS2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_19_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2718_ net36 net744 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput352 net352 VGND VGND VPWR VPWR W2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput341 net341 VGND VGND VPWR VPWR SS4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput330 net330 VGND VGND VPWR VPWR SS4BEG[11] sky130_fd_sc_hd__buf_2
X_2649_ net776 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput363 net363 VGND VGND VPWR VPWR W2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput385 net385 VGND VGND VPWR VPWR WW4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput374 net374 VGND VGND VPWR VPWR W6BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1951_ net638 net689 Inst_RegFile_switch_matrix.JS2BEG1 _0377_ Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.W1BEG2
+ sky130_fd_sc_hd__mux4_2
X_1882_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q _0766_ Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q
+ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__a21bo_1
X_2503_ net760 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2434_ net766 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2365_ net772 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1316_ _0253_ _0252_ net678 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2296_ clknet_4_4_0_UserCLK_regs _0054_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1247_ net60 net84 net68 net784 Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q
+ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux4_1
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1178_ _1068_ _1069_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR VPWR
+ _1070_ sky130_fd_sc_hd__mux2_1
XFILLER_64_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_31 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 FrameData[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_53 N4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 NN4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 NN4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 FrameStrobe[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 W2END[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 net693 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput160 net160 VGND VGND VPWR VPWR E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput171 net171 VGND VGND VPWR VPWR E6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput193 net193 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput182 net182 VGND VGND VPWR VPWR EE4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2150_ net600 net529 _0948_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux2_4
X_1101_ Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__inv_2
X_2081_ net484 net606 _0925_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__mux2_4
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2983_ SS4END[7] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_2
X_1934_ Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q _0814_ Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q
+ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__a21oi_1
Xinput40 FrameData[21] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
X_1865_ Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q _0752_ VGND VGND VPWR VPWR _0753_
+ sky130_fd_sc_hd__and2b_1
Xinput62 N2END[0] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
Xinput73 N2MID[3] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
X_1796_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0692_ VGND VGND VPWR VPWR _0693_
+ sky130_fd_sc_hd__and2b_1
Xinput51 FrameData[3] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
Xinput95 S2END[5] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_6
Xinput84 NN4END[2] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_4
X_2417_ net752 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2348_ net780 net57 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2279_ clknet_4_14_0_UserCLK_regs _0037_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[17\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1650_ _0564_ _0561_ Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q VGND VGND VPWR VPWR
+ A_ADR0 sky130_fd_sc_hd__mux2_4
Xhold109 Inst_RegFile_32x4.mem\[31\]\[2\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
X_1581_ _0500_ _0499_ net688 VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux2_1
X_2202_ _0920_ _0958_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__nand2_8
X_2133_ net458 net607 _0945_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__mux2_4
XFILLER_81_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2064_ net99 net127 Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q VGND VGND VPWR VPWR
+ _0915_ sky130_fd_sc_hd__mux2_1
XFILLER_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2966_ S4END[6] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_32_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1917_ _0799_ Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q
+ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a21oi_2
X_2897_ Inst_RegFile_switch_matrix.JN2BEG1 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_8
X_1848_ Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q net635 VGND VGND VPWR VPWR _0738_
+ sky130_fd_sc_hd__or2_1
X_1779_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__inv_1
XFILLER_72_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone21 net656 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkbuf_1
Xclone54 net679 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2820_ E6END[10] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_1
X_2751_ clknet_4_12_0_UserCLK_regs _0087_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[31\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1702_ net7 net92 net782 net120 Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q
+ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__mux4_1
X_2682_ net775 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1633_ Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q _0549_ VGND VGND VPWR VPWR _0550_
+ sky130_fd_sc_hd__nand2_1
X_1564_ _0485_ _0484_ net685 VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
X_1495_ Inst_RegFile_32x4.mem\[12\]\[0\] Inst_RegFile_32x4.mem\[13\]\[0\] net432 VGND
+ VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux2_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2116_ net601 net526 _0938_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__mux2_4
XFILLER_81_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2047_ _0897_ _0899_ Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q VGND VGND VPWR VPWR
+ _0900_ sky130_fd_sc_hd__mux2_2
XFILLER_54_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2949_ Inst_RegFile_switch_matrix.JS2BEG1 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_9_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1280_ _0219_ _0218_ net679 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2803_ Inst_RegFile_switch_matrix.E2BEG7 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_14_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2734_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.BD_comb\[2\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.BD_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2665_ net758 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2596_ net764 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1616_ Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q _0533_ VGND VGND VPWR VPWR _0534_
+ sky130_fd_sc_hd__or2_1
X_1547_ Inst_RegFile_32x4.mem\[26\]\[3\] Inst_RegFile_32x4.mem\[27\]\[3\] net628 VGND
+ VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux2_1
XFILLER_86_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1478_ _0404_ _0401_ Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JN2BEG6 sky130_fd_sc_hd__mux2_4
XFILLER_86_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout750 FrameData[7] VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout761 net762 VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__clkbuf_4
Xfanout772 net35 VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__clkbuf_4
Xfanout783 net4 VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__clkbuf_4
XFILLER_73_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_121 W2MID[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_110 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2450_ net751 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_53_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1401_ _0331_ _0332_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q VGND VGND VPWR VPWR
+ _0333_ sky130_fd_sc_hd__mux2_4
XFILLER_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2381_ net38 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1332_ Inst_RegFile_32x4.mem\[0\]\[2\] Inst_RegFile_32x4.mem\[1\]\[2\] net614 VGND
+ VGND VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_1
X_1263_ net72 net100 Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q VGND VGND VPWR VPWR
+ _0203_ sky130_fd_sc_hd__mux2_1
X_3002_ Inst_RegFile_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_6
Xinput5 E2END[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1194_ Inst_RegFile_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__inv_1
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2717_ net35 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput353 net353 VGND VGND VPWR VPWR W2BEG[4] sky130_fd_sc_hd__buf_8
Xoutput320 net320 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput331 Inst_RegFile_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR SS4BEG[12] sky130_fd_sc_hd__buf_6
Xoutput342 net342 VGND VGND VPWR VPWR SS4BEG[8] sky130_fd_sc_hd__buf_2
X_2648_ net777 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2579_ net749 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput386 net386 VGND VGND VPWR VPWR WW4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput364 net364 VGND VGND VPWR VPWR W2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput375 net375 VGND VGND VPWR VPWR W6BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1950_ net414 _0407_ Inst_RegFile_switch_matrix.JS2BEG2 _0827_ Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__mux4_2
X_1881_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q _0767_ VGND VGND VPWR VPWR _0768_
+ sky130_fd_sc_hd__and2b_1
X_2502_ net761 net705 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2433_ net767 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2364_ net773 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1315_ Inst_RegFile_32x4.mem\[18\]\[1\] Inst_RegFile_32x4.mem\[19\]\[1\] net618 VGND
+ VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2295_ clknet_4_4_0_UserCLK_regs _0053_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1246_ net11 net88 net96 net114 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux4_1
X_1177_ net88 net96 net112 net114 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__mux4_1
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_10 EE4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 FrameStrobe[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 NN4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 N4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_43 FrameStrobe[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 net722 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 net307 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_87 net365 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput150 Inst_RegFile_switch_matrix.E2BEG6 VGND VGND VPWR VPWR E2BEG[6] sky130_fd_sc_hd__buf_8
Xoutput161 net161 VGND VGND VPWR VPWR E6BEG[10] sky130_fd_sc_hd__buf_6
Xoutput194 net194 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput172 net172 VGND VGND VPWR VPWR EE4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput183 net183 VGND VGND VPWR VPWR EE4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_47_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1100_ Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__inv_2
X_2080_ net469 net610 _0925_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__mux2_4
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2982_ SS4END[6] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_72_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1933_ net114 net648 Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR
+ _0814_ sky130_fd_sc_hd__mux2_1
Xinput30 FrameData[12] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
X_1864_ net674 net660 Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q VGND VGND VPWR VPWR
+ _0752_ sky130_fd_sc_hd__mux2_1
Xinput41 FrameData[22] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xinput52 FrameData[4] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
Xinput63 N2END[1] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
X_1795_ net672 net658 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q VGND VGND VPWR VPWR
+ _0692_ sky130_fd_sc_hd__mux2_1
Xinput96 S2END[6] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 NN4END[3] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xinput74 N2MID[4] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
XFILLER_69_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2416_ net753 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2347_ net50 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2278_ clknet_4_14_0_UserCLK_regs _0036_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[17\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1229_ Inst_RegFile_32x4.mem\[14\]\[0\] Inst_RegFile_32x4.mem\[15\]\[0\] net395 VGND
+ VGND VPWR VPWR _0171_ sky130_fd_sc_hd__mux2_1
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1580_ Inst_RegFile_32x4.mem\[24\]\[2\] Inst_RegFile_32x4.mem\[25\]\[2\] net628 VGND
+ VGND VPWR VPWR _0500_ sky130_fd_sc_hd__mux2_1
X_2201_ net600 net456 _0959_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__mux2_4
X_2132_ net519 net611 _0945_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__mux2_4
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2063_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_49_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2965_ S4END[5] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_32_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1916_ net88 net660 Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q VGND VGND VPWR VPWR
+ _0799_ sky130_fd_sc_hd__mux2_2
X_2896_ Inst_RegFile_switch_matrix.JN2BEG0 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_8
XFILLER_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1847_ net61 net783 net692 net653 Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q
+ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__mux4_1
X_1778_ net672 net659 Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q VGND VGND VPWR VPWR
+ _0676_ sky130_fd_sc_hd__mux2_1
XFILLER_1_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone22 net671 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__buf_8
Xclone55 net642 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2750_ clknet_4_12_0_UserCLK_regs _0086_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[31\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1701_ _0608_ _1013_ Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q VGND VGND VPWR VPWR
+ _0609_ sky130_fd_sc_hd__o21a_1
X_2681_ net776 net730 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1632_ net105 net133 Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q VGND VGND VPWR VPWR
+ _0549_ sky130_fd_sc_hd__mux2_1
X_1563_ Inst_RegFile_32x4.mem\[8\]\[3\] Inst_RegFile_32x4.mem\[9\]\[3\] net623 VGND
+ VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux2_1
X_1494_ _0418_ _0419_ net685 VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux2_1
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2115_ net629 net494 _0938_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__mux2_4
XFILLER_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2046_ _0804_ _0898_ Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q VGND VGND VPWR VPWR
+ _0899_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2948_ Inst_RegFile_switch_matrix.JS2BEG0 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__buf_6
XFILLER_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2879_ net705 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2733_ clknet_4_9_0_UserCLK_regs Inst_RegFile_32x4.BD_comb\[1\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.BD_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2664_ net759 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2595_ net42 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1615_ net692 net673 net659 net655 Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__mux4_1
XFILLER_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1546_ Inst_RegFile_32x4.BD_comb\[1\] Inst_RegFile_32x4.BD_reg\[1\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR BD1 sky130_fd_sc_hd__mux2_4
X_1477_ _0402_ _0403_ Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q VGND VGND VPWR VPWR
+ _0404_ sky130_fd_sc_hd__mux2_1
XFILLER_82_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2029_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q _0807_ VGND VGND VPWR VPWR _0883_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_40_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout751 net54 VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__buf_2
Xfanout740 FrameStrobe[10] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout762 FrameData[26] VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__buf_2
Xfanout784 net3 VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout773 net34 VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__clkbuf_4
XFILLER_85_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_100 net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _0827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_111 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1400_ net26 net87 net89 net95 Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux4_2
XFILLER_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2380_ net780 net740 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1331_ Inst_RegFile_32x4.mem\[2\]\[2\] Inst_RegFile_32x4.mem\[3\]\[2\] net614 VGND
+ VGND VPWR VPWR _0267_ sky130_fd_sc_hd__mux2_1
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1262_ Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q net128 Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q
+ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__o21a_1
X_3001_ Inst_RegFile_switch_matrix.JW2BEG0 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__buf_6
Xinput6 E2END[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
X_1193_ _0132_ _0134_ _0137_ _1002_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JS2BEG3
+ sky130_fd_sc_hd__a22o_4
XFILLER_51_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2716_ net34 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput310 net310 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__buf_2
X_2647_ net778 net726 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput321 net321 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput332 net332 VGND VGND VPWR VPWR SS4BEG[13] sky130_fd_sc_hd__buf_8
Xoutput343 net343 VGND VGND VPWR VPWR SS4BEG[9] sky130_fd_sc_hd__buf_2
X_2578_ net751 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput354 Inst_RegFile_switch_matrix.JW2BEG5 VGND VGND VPWR VPWR W2BEG[5] sky130_fd_sc_hd__buf_6
Xoutput387 net387 VGND VGND VPWR VPWR WW4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput365 net365 VGND VGND VPWR VPWR W6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput376 net376 VGND VGND VPWR VPWR W6BEG[9] sky130_fd_sc_hd__buf_2
X_1529_ Inst_RegFile_32x4.mem\[14\]\[1\] Inst_RegFile_32x4.mem\[15\]\[1\] net621 VGND
+ VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux2_1
XFILLER_59_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _0697_ _0698_ Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _0767_ sky130_fd_sc_hd__mux2_1
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2501_ net763 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2432_ net768 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2363_ net33 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1314_ Inst_RegFile_32x4.mem\[16\]\[1\] Inst_RegFile_32x4.mem\[17\]\[1\] net618 VGND
+ VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_16_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2294_ clknet_4_4_0_UserCLK_regs _0052_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1245_ _0185_ _0186_ Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q VGND VGND VPWR VPWR
+ _0187_ sky130_fd_sc_hd__mux2_4
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1176_ net60 net68 net784 net11 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__mux4_1
XFILLER_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_11 EE4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net193 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 FrameStrobe[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 NN4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 N4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 net318 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_88 net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 net732 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput140 Inst_RegFile_switch_matrix.E1BEG0 VGND VGND VPWR VPWR E1BEG[0] sky130_fd_sc_hd__buf_6
Xoutput151 net151 VGND VGND VPWR VPWR E2BEG[7] sky130_fd_sc_hd__buf_4
Xoutput195 net195 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput162 Inst_RegFile_switch_matrix.E6BEG1 VGND VGND VPWR VPWR E6BEG[11] sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_34_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput173 net173 VGND VGND VPWR VPWR EE4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput184 net184 VGND VGND VPWR VPWR EE4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2981_ SS4END[5] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_72_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1932_ _1010_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q
+ _0812_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__a211o_1
X_1863_ _0748_ _0749_ _0750_ Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__a221o_1
Xinput31 FrameData[13] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xinput20 E2MID[7] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
Xinput42 FrameData[23] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
Xinput64 N2END[2] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
X_1794_ net419 net648 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q VGND VGND VPWR VPWR
+ _0691_ sky130_fd_sc_hd__mux2_1
Xinput53 FrameData[5] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
Xinput97 S2END[7] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_2
Xinput86 S1END[0] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
Xinput75 N2MID[5] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
X_2415_ net754 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2346_ net756 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2277_ clknet_4_2_0_UserCLK_regs _0035_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1228_ Inst_RegFile_32x4.mem\[12\]\[0\] Inst_RegFile_32x4.mem\[13\]\[0\] net394 VGND
+ VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_1
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1159_ net782 net94 net113 net122 Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__mux4_1
XFILLER_52_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2200_ net630 net453 _0959_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__mux2_4
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2131_ _0944_ _0924_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__nor2_8
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2062_ net71 net14 Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q VGND VGND VPWR VPWR
+ _0913_ sky130_fd_sc_hd__mux2_1
XFILLER_19_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2964_ S4END[4] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1915_ Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q _0797_ VGND VGND VPWR VPWR _0798_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_32_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1846_ Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q _0730_ _0732_ _0734_ _0736_ VGND
+ VGND VPWR VPWR Inst_RegFile_switch_matrix.SS4BEG2 sky130_fd_sc_hd__a32oi_1
X_1777_ _0672_ _0673_ _0674_ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2329_ net776 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone23 net661 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone12 net412 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__buf_8
XFILLER_4_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2680_ net777 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1700_ net682 net635 net666 net640 Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q
+ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__mux4_2
X_1631_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__inv_1
X_1562_ Inst_RegFile_32x4.mem\[10\]\[3\] Inst_RegFile_32x4.mem\[11\]\[3\] net623 VGND
+ VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux2_1
X_1493_ Inst_RegFile_32x4.mem\[10\]\[0\] Inst_RegFile_32x4.mem\[11\]\[0\] net623 VGND
+ VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
X_2114_ net605 net549 _0938_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__mux2_4
XFILLER_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2045_ net25 net125 net108 Inst_RegFile_switch_matrix.E2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_80_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2878_ net710 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_1
X_1829_ net60 net88 net693 net658 Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q
+ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__mux4_1
XFILLER_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_8_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_8_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2801_ Inst_RegFile_switch_matrix.E2BEG5 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_14_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2732_ clknet_4_8_0_UserCLK_regs Inst_RegFile_32x4.BD_comb\[0\] VGND VGND VPWR VPWR
+ Inst_RegFile_32x4.BD_reg\[0\] sky130_fd_sc_hd__dfxtp_1
X_2663_ net45 net726 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2594_ net41 net718 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1614_ Inst_RegFile_32x4.BD_comb\[2\] Inst_RegFile_32x4.BD_reg\[2\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR BD2 sky130_fd_sc_hd__mux2_4
XFILLER_5_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1545_ _0468_ _0448_ _0409_ VGND VGND VPWR VPWR Inst_RegFile_32x4.BD_comb\[1\] sky130_fd_sc_hd__mux2_4
X_1476_ net12 net89 net97 net115 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__mux4_1
XFILLER_79_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2028_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q _0828_ VGND VGND VPWR VPWR _0882_
+ sky130_fd_sc_hd__nand2_1
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout730 FrameStrobe[1] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkbuf_2
Xfanout741 net742 VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__clkbuf_2
Xfanout763 net44 VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__buf_4
Xfanout774 net33 VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__clkbuf_4
Xfanout752 net53 VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__clkbuf_4
XFILLER_73_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_123 net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_101 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1330_ _0262_ _0265_ net663 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_4
X_1261_ _0195_ _0197_ _0200_ _0973_ _0971_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a221o_1
X_1192_ _0135_ _0136_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q VGND VGND VPWR VPWR
+ _0137_ sky130_fd_sc_hd__mux2_1
Xinput7 E2END[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
X_3000_ Inst_RegFile_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__buf_6
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2715_ net774 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput300 net300 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__buf_8
X_2646_ net779 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput344 net344 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
Xoutput311 net311 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput322 net322 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput333 net333 VGND VGND VPWR VPWR SS4BEG[14] sky130_fd_sc_hd__buf_4
X_2577_ net752 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput355 net355 VGND VGND VPWR VPWR W2BEG[6] sky130_fd_sc_hd__buf_4
Xoutput377 net377 VGND VGND VPWR VPWR WW4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput366 Inst_RegFile_switch_matrix.W6BEG0 VGND VGND VPWR VPWR W6BEG[10] sky130_fd_sc_hd__buf_8
X_1528_ _0993_ net622 net685 _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__o211a_1
Xoutput388 net388 VGND VGND VPWR VPWR WW4BEG[5] sky130_fd_sc_hd__buf_2
X_1459_ _0383_ _0381_ _0386_ Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG6 sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_2_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2500_ net764 net704 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2431_ net770 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2362_ net32 net738 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2293_ clknet_4_6_0_UserCLK_regs _0051_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1313_ _0247_ _0250_ net664 VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__mux2_1
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1244_ net405 BD0 BD2 net412 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux4_2
X_1175_ _1066_ _0999_ Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q VGND VGND VPWR VPWR
+ _1067_ sky130_fd_sc_hd__o21a_1
XFILLER_64_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 EE4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 net193 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 FrameStrobe[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 N4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 NN4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 net319 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_89 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2629_ net763 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput152 net152 VGND VGND VPWR VPWR E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput141 net141 VGND VGND VPWR VPWR E1BEG[1] sky130_fd_sc_hd__buf_8
Xoutput185 net185 VGND VGND VPWR VPWR EE4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput174 net174 VGND VGND VPWR VPWR EE4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput163 net163 VGND VGND VPWR VPWR E6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput196 net196 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__buf_2
XFILLER_46_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2980_ SS4END[4] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_72_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1931_ net58 Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR _0812_
+ sky130_fd_sc_hd__nor2_1
X_1862_ net113 net693 Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q VGND VGND VPWR VPWR
+ _0750_ sky130_fd_sc_hd__mux2_1
Xinput10 E2END[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_6
Xinput21 E6END[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
X_1793_ _1021_ _0675_ _0680_ _0690_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.W6BEG1
+ sky130_fd_sc_hd__a31o_4
Xinput43 FrameData[24] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 FrameData[14] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput54 FrameData[6] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
Xinput98 S2MID[0] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
Xinput87 S1END[1] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_4
Xinput65 N2END[3] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xinput76 N2MID[6] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
X_2414_ net757 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2345_ net758 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2276_ clknet_4_1_0_UserCLK_regs _0034_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1227_ _1005_ _0154_ _0167_ _0168_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__a2bb2o_4
X_1158_ net60 net66 net78 net9 Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__mux4_1
XFILLER_37_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1089_ net130 VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__inv_2
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2130_ _0941_ _0854_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__nand2_8
XFILLER_66_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2061_ Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q _0909_ _0910_ _0911_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__a221o_1
XFILLER_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2963_ net105 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_2
X_1914_ net60 net784 Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q VGND VGND VPWR VPWR
+ _0797_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2894_ Inst_RegFile_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_6
X_1845_ Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q _0735_ Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q
+ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_62_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1776_ net112 net693 Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q VGND VGND VPWR VPWR
+ _0674_ sky130_fd_sc_hd__mux2_1
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2328_ net777 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2259_ clknet_4_3_0_UserCLK_regs _0017_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[28\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone35 net635 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__buf_6
Xclone24 net663 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkbuf_1
Xclone13 AD3 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1630_ net77 net20 Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q VGND VGND VPWR VPWR
+ _0547_ sky130_fd_sc_hd__mux2_1
X_1561_ _0475_ _0482_ _0394_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__mux2_1
X_1492_ Inst_RegFile_32x4.mem\[8\]\[0\] Inst_RegFile_32x4.mem\[9\]\[0\] net623 VGND
+ VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2113_ net609 net562 _0938_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux2_4
XFILLER_66_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2044_ _0406_ _0697_ Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q VGND VGND VPWR VPWR
+ _0897_ sky130_fd_sc_hd__mux2_1
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2877_ net714 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
X_1828_ Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q _0720_ Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q
+ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__o21ai_1
X_1759_ net649 net684 net668 net637 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__mux4_1
XFILLER_57_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2731_ net755 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2662_ net761 net726 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2593_ net40 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1613_ _0532_ _0513_ _0409_ VGND VGND VPWR VPWR Inst_RegFile_32x4.BD_comb\[2\] sky130_fd_sc_hd__mux2_4
X_1544_ _0456_ _0457_ _0461_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__o2bb2a_1
X_1475_ net61 net69 net83 net783 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux4_1
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2027_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q _0698_ Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q
+ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__a21oi_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2929_ NN4END[5] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__buf_1
XFILLER_49_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout731 net732 VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__buf_2
Xfanout720 FrameStrobe[3] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout742 FrameStrobe[10] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__buf_2
Xfanout764 net43 VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__clkbuf_4
Xfanout775 net32 VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__clkbuf_4
Xfanout753 net52 VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__clkbuf_4
XFILLER_85_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_124 net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_113 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1260_ _0195_ _0197_ _0200_ _0973_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG6
+ sky130_fd_sc_hd__a22o_4
XFILLER_49_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1191_ net21 net94 net106 net122 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__mux4_1
Xinput8 E2END[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_19_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2714_ net775 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput301 Inst_RegFile_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__buf_8
X_2645_ net747 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput312 net312 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput323 net323 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput334 net334 VGND VGND VPWR VPWR SS4BEG[15] sky130_fd_sc_hd__buf_6
Xoutput345 net345 VGND VGND VPWR VPWR W1BEG[0] sky130_fd_sc_hd__buf_6
X_2576_ net753 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput356 net356 VGND VGND VPWR VPWR W2BEG[7] sky130_fd_sc_hd__buf_6
Xoutput378 net378 VGND VGND VPWR VPWR WW4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput367 Inst_RegFile_switch_matrix.W6BEG1 VGND VGND VPWR VPWR W6BEG[11] sky130_fd_sc_hd__buf_8
X_1527_ Inst_RegFile_32x4.mem\[11\]\[1\] net622 VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__nand2_1
Xoutput389 net389 VGND VGND VPWR VPWR WW4BEG[6] sky130_fd_sc_hd__buf_2
X_1458_ _0384_ _0385_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q VGND VGND VPWR VPWR
+ _0386_ sky130_fd_sc_hd__mux2_1
XFILLER_59_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1389_ _0209_ _0304_ _0322_ _0313_ VGND VGND VPWR VPWR Inst_RegFile_32x4.AD_comb\[3\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2430_ net771 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_51_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2361_ net31 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2292_ clknet_4_4_0_UserCLK_regs _0050_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1312_ _0248_ _0249_ net446 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
X_1243_ net693 net674 net660 net656 Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__mux4_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1174_ net649 net683 net428 net641 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_75_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_13 EE4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_46 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 FrameStrobe[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 N4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 NN4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 net333 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2628_ net43 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput142 Inst_RegFile_switch_matrix.E1BEG2 VGND VGND VPWR VPWR E1BEG[2] sky130_fd_sc_hd__buf_8
X_2559_ net37 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput153 net153 VGND VGND VPWR VPWR E2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput164 net164 VGND VGND VPWR VPWR E6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput175 net175 VGND VGND VPWR VPWR EE4BEG[12] sky130_fd_sc_hd__buf_6
Xoutput186 net186 VGND VGND VPWR VPWR EE4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput197 net197 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
XFILLER_47_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1930_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q _1045_ _0810_ Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q
+ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__a211o_1
X_1861_ net85 Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__o21ba_1
Xinput11 E2END[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 E6END[1] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
X_1792_ Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q _0689_ Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q
+ _0688_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__o211a_1
Xinput44 FrameData[25] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xinput33 FrameData[15] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_2
Xinput55 FrameData[8] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xinput88 S1END[2] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xinput66 N2END[4] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
Xinput77 N2MID[7] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput99 S2MID[1] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
X_2413_ net769 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2344_ net759 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2275_ clknet_4_1_0_UserCLK_regs _0033_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1226_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q _0163_ _1005_ VGND VGND VPWR VPWR
+ _0168_ sky130_fd_sc_hd__o21a_1
XFILLER_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1157_ _0990_ _1049_ Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q VGND VGND VPWR VPWR
+ _1050_ sky130_fd_sc_hd__o21a_1
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1088_ Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_35_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2060_ net70 Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q
+ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__o21ba_1
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2962_ net104 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_1
X_1913_ Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q _0795_ _0793_ Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q
+ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__o211a_1
X_2893_ Inst_RegFile_switch_matrix.N1BEG1 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__buf_6
X_1844_ net114 net647 Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q VGND VGND VPWR VPWR
+ _0735_ sky130_fd_sc_hd__mux2_1
X_1775_ net84 Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__o21ba_1
XFILLER_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2327_ net778 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2258_ clknet_4_6_0_UserCLK_regs _0016_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[28\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1209_ net26 net137 net106 Inst_RegFile_switch_matrix.JW2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_83_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2189_ net501 net632 _0956_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__mux2_2
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone25 net644 VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_6
Xclone14 net669 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__buf_8
Xclone36 net637 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__buf_8
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1560_ _0478_ _0481_ net645 VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux2_1
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1491_ _0398_ _0416_ _0394_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
XFILLER_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2112_ _0920_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__nand2_8
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2043_ net471 net610 _0888_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_80_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2876_ net718 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
X_1827_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__inv_1
X_1758_ net693 net673 net659 net654 Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux4_1
X_1689_ _0598_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG1 sky130_fd_sc_hd__inv_2
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2730_ net756 net743 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2661_ net44 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1612_ net397 _0517_ _0521_ _0531_ _0525_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__o32a_4
X_2592_ net39 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1543_ net643 _0463_ _0466_ _0393_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__a31o_1
X_1474_ _0399_ _0400_ Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q VGND VGND VPWR VPWR
+ _0401_ sky130_fd_sc_hd__mux2_2
XFILLER_79_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2026_ Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q _0860_ VGND VGND VPWR VPWR _0880_
+ sky130_fd_sc_hd__or2_1
XFILLER_35_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2928_ NN4END[4] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_1
X_2859_ net770 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout721 net722 VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__buf_2
Xfanout732 net734 VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__buf_2
Xfanout710 FrameStrobe[6] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__clkbuf_2
Xfanout765 net42 VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout743 net744 VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__clkbuf_2
Xfanout754 net51 VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__buf_4
Xfanout776 net31 VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__clkbuf_4
XFILLER_73_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_103 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 net139 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_4_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_4_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1190_ net66 net9 net784 net26 Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q
+ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__mux4_1
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 E2END[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_19_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2713_ net31 net744 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2644_ net748 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2575_ net754 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput324 net324 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput313 net313 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput335 net335 VGND VGND VPWR VPWR SS4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput302 net302 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput346 Inst_RegFile_switch_matrix.W1BEG1 VGND VGND VPWR VPWR W1BEG[1] sky130_fd_sc_hd__buf_6
Xoutput357 net357 VGND VGND VPWR VPWR W2BEGb[0] sky130_fd_sc_hd__buf_2
X_1526_ net685 _0449_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__nor2_1
Xoutput368 net368 VGND VGND VPWR VPWR W6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput379 net379 VGND VGND VPWR VPWR WW4BEG[11] sky130_fd_sc_hd__buf_2
X_1457_ net87 net97 net89 net692 Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__mux4_1
XFILLER_67_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1388_ _0321_ _0317_ net651 _0209_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__a31oi_1
XFILLER_67_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2009_ net65 net93 Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q VGND VGND VPWR VPWR
+ _0863_ sky130_fd_sc_hd__mux2_1
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2360_ net30 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2291_ clknet_4_1_0_UserCLK_regs _0049_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1311_ Inst_RegFile_32x4.mem\[28\]\[1\] Inst_RegFile_32x4.mem\[29\]\[1\] net615 VGND
+ VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1242_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q Inst_RegFile_switch_matrix.JS2BEG5
+ Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__o21a_1
XFILLER_49_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q _1064_ VGND VGND VPWR VPWR _1065_
+ sky130_fd_sc_hd__or2_1
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_14 EE4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_47 net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 FrameStrobe[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_58 N4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 NN4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2627_ net765 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput143 Inst_RegFile_switch_matrix.E1BEG3 VGND VGND VPWR VPWR E1BEG[3] sky130_fd_sc_hd__buf_8
Xoutput165 net165 VGND VGND VPWR VPWR E6BEG[3] sky130_fd_sc_hd__buf_2
X_2558_ net36 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput154 net154 VGND VGND VPWR VPWR E2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput176 Inst_RegFile_switch_matrix.EE4BEG1 VGND VGND VPWR VPWR EE4BEG[13] sky130_fd_sc_hd__buf_6
Xoutput198 net198 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
X_1509_ Inst_RegFile_32x4.BD_comb\[0\] Inst_RegFile_32x4.BD_reg\[0\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR BD0 sky130_fd_sc_hd__mux2_4
Xoutput187 net187 VGND VGND VPWR VPWR EE4BEG[9] sky130_fd_sc_hd__buf_2
X_2489_ net776 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1860_ net784 Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q VGND VGND VPWR VPWR _0748_
+ sky130_fd_sc_hd__nand2b_1
X_1791_ net683 net428 net667 net447 Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q
+ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__mux4_1
Xinput12 E2END[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
Xinput45 FrameData[27] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
Xinput34 FrameData[16] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput23 EE4END[0] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
Xinput89 S1END[3] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_6
Xinput56 FrameData[9] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
Xinput78 N4END[0] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
Xinput67 N2END[5] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_6
X_2412_ net780 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2343_ net760 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2274_ clknet_4_1_0_UserCLK_regs _0032_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1225_ _1004_ _0165_ _0166_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__o21ai_1
X_1156_ net681 net634 net406 net639 Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q
+ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__mux4_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1087_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_35_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1989_ _1027_ _0191_ _0840_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__a22o_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2961_ net103 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__buf_1
X_1912_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__inv_1
XFILLER_63_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2892_ Inst_RegFile_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__buf_6
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1843_ _1010_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__a211o_1
X_1774_ net784 Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q VGND VGND VPWR VPWR _0672_
+ sky130_fd_sc_hd__nand2b_1
X_2326_ net779 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2257_ clknet_4_15_0_UserCLK_regs _0015_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[27\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1208_ _0151_ _0148_ Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JW2BEG3 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_83_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2188_ net544 net606 _0956_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__mux2_4
XFILLER_80_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1139_ _1032_ _0995_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__or2_4
XFILLER_80_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone15 net653 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__buf_8
Xclone26 N1END[1] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1490_ _0412_ _0415_ net645 VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
XFILLER_79_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2111_ _0936_ _0854_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__nor2_8
XFILLER_66_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2042_ _0895_ _0889_ Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q VGND VGND VPWR VPWR
+ _0896_ sky130_fd_sc_hd__mux2_2
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2944_ Inst_RegFile_switch_matrix.S1BEG0 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_6
X_2875_ net722 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
X_1826_ net667 _0697_ Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q VGND VGND VPWR VPWR
+ _0719_ sky130_fd_sc_hd__mux2_1
X_1757_ _0654_ _0652_ _0657_ _1020_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E2BEG0
+ sky130_fd_sc_hd__a22o_1
X_1688_ Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q _0595_ _0597_ _0593_ _0591_ VGND
+ VGND VPWR VPWR _0598_ sky130_fd_sc_hd__o32a_4
XFILLER_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2309_ clknet_4_6_0_UserCLK_regs _0067_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_12_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_12_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_79_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2660_ net43 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1611_ _0527_ net643 _0530_ _0393_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a31o_1
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2591_ net770 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1542_ net686 _0465_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__nand2_1
X_1473_ net648 net683 net667 net642 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux4_1
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2025_ _0878_ _0865_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__or2_4
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2927_ Inst_RegFile_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__buf_4
X_2858_ net771 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
X_2789_ clknet_4_1_0_UserCLK_regs _0125_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1809_ net418 net87 net115 net672 Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q
+ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_68_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout700 net701 VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout722 FrameStrobe[3] VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__clkbuf_4
Xfanout711 FrameStrobe[5] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__buf_2
Xfanout733 net734 VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__clkbuf_4
Xfanout766 net41 VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout744 net746 VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout755 net50 VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__buf_4
XFILLER_85_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout777 net30 VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__clkbuf_4
XFILLER_73_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_115 EE4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_104 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2712_ net30 net746 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2643_ net749 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2574_ net757 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput303 net303 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__buf_8
Xoutput325 net325 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput314 net314 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__buf_2
X_1525_ Inst_RegFile_32x4.mem\[8\]\[1\] Inst_RegFile_32x4.mem\[9\]\[1\] net622 VGND
+ VGND VPWR VPWR _0449_ sky130_fd_sc_hd__mux2_1
Xoutput347 Inst_RegFile_switch_matrix.W1BEG2 VGND VGND VPWR VPWR W1BEG[2] sky130_fd_sc_hd__buf_6
Xoutput336 net336 VGND VGND VPWR VPWR SS4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput358 net358 VGND VGND VPWR VPWR W2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput369 net369 VGND VGND VPWR VPWR W6BEG[2] sky130_fd_sc_hd__buf_2
X_1456_ net61 net69 net783 net12 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_2_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1387_ net675 _0320_ _0319_ net662 VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__o211ai_1
XFILLER_82_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2008_ _1030_ _0860_ _0861_ _1031_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__a211o_1
XFILLER_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2290_ clknet_4_4_0_UserCLK_regs _0048_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1310_ Inst_RegFile_32x4.mem\[30\]\[1\] Inst_RegFile_32x4.mem\[31\]\[1\] net615 VGND
+ VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1241_ Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q _0162_ VGND VGND VPWR VPWR _0183_
+ sky130_fd_sc_hd__nand2_1
X_1172_ net693 net672 net658 net419 Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_67_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_48 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 EE4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 N4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2626_ net766 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput144 net144 VGND VGND VPWR VPWR E2BEG[0] sky130_fd_sc_hd__buf_8
Xoutput155 net155 VGND VGND VPWR VPWR E2BEGb[3] sky130_fd_sc_hd__buf_2
X_2557_ net35 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput166 net166 VGND VGND VPWR VPWR E6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput177 net177 VGND VGND VPWR VPWR EE4BEG[14] sky130_fd_sc_hd__buf_8
Xoutput199 net199 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput188 net188 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
X_1508_ _0433_ _0417_ _0409_ VGND VGND VPWR VPWR Inst_RegFile_32x4.BD_comb\[0\] sky130_fd_sc_hd__mux2_4
X_2488_ net777 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1439_ _0354_ _0353_ _0364_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__o22a_1
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1790_ _0687_ _0685_ Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q VGND VGND VPWR VPWR
+ _0688_ sky130_fd_sc_hd__o21ai_2
Xinput13 E2MID[0] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
Xinput46 FrameData[28] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput35 FrameData[17] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput24 EE4END[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput79 N4END[1] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
Xinput68 N2END[6] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
Xinput57 FrameStrobe[11] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
X_2411_ net755 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2342_ net761 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2273_ clknet_4_5_0_UserCLK_regs _0031_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1224_ Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q _0164_ Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__o21a_1
XFILLER_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1155_ Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q _1047_ VGND VGND VPWR VPWR _1048_
+ sky130_fd_sc_hd__or2_4
XFILLER_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1086_ net102 VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__inv_1
XFILLER_52_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1988_ Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q _0841_ Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q
+ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__o21a_1
X_2609_ net752 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_75_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2960_ net102 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_2
X_2891_ FrameStrobe[19] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_1
X_1911_ net668 _0697_ Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q VGND VGND VPWR VPWR
+ _0794_ sky130_fd_sc_hd__mux2_1
X_1842_ net58 Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q VGND VGND VPWR VPWR _0733_
+ sky130_fd_sc_hd__nor2_1
X_1773_ _0671_ _0668_ Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JN2BEG0 sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_31_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2325_ net747 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2256_ clknet_4_13_0_UserCLK_regs _0014_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[27\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1207_ _0149_ _0150_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q VGND VGND VPWR VPWR
+ _0151_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2187_ net523 net609 _0956_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_40_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1138_ net650 net684 net398 net404 Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__mux4_2
XFILLER_80_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone27 net655 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2110_ _0838_ _0846_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__nand2_4
X_2041_ _1026_ _0890_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__a21o_1
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2943_ Inst_RegFile_switch_matrix.NN4BEG3 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_2
X_2874_ net726 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1825_ Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q _0366_ _0717_ VGND VGND VPWR VPWR
+ _0718_ sky130_fd_sc_hd__a21oi_1
X_1756_ _0655_ _0656_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q VGND VGND VPWR VPWR
+ _0657_ sky130_fd_sc_hd__mux2_1
X_1687_ _1009_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__nor2_1
XFILLER_85_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2308_ clknet_4_7_0_UserCLK_regs _0066_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2239_ net604 net543 _0967_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_4
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1610_ net686 _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__nand2_1
X_2590_ net771 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1541_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__inv_1
X_1472_ net692 net673 net659 net655 Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__mux4_1
XFILLER_67_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2024_ _0867_ Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q _0871_ _0877_ VGND VGND
+ VPWR VPWR _0878_ sky130_fd_sc_hd__a22o_4
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2857_ net772 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_1
X_1808_ _0696_ _0704_ Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.W6BEG0 sky130_fd_sc_hd__mux2_4
X_2788_ clknet_4_1_0_UserCLK_regs _0124_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1739_ net63 net6 net783 net781 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__mux4_1
Xfanout723 net724 VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__clkbuf_2
Xfanout712 FrameStrobe[5] VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout701 FrameStrobe[8] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__buf_2
XFILLER_49_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout767 net40 VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__clkbuf_4
Xfanout756 net49 VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout734 FrameStrobe[12] VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__buf_1
Xfanout745 net746 VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__clkbuf_2
Xfanout778 net29 VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__clkbuf_4
XFILLER_73_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_116 EE4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_105 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2711_ net29 net744 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2642_ net751 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2573_ net769 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput304 net304 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput326 net326 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput315 net315 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__buf_4
Xoutput348 net348 VGND VGND VPWR VPWR W1BEG[3] sky130_fd_sc_hd__buf_6
Xoutput337 net337 VGND VGND VPWR VPWR SS4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput359 net359 VGND VGND VPWR VPWR W2BEGb[2] sky130_fd_sc_hd__buf_2
X_1524_ _0440_ _0447_ _0394_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__mux2_4
X_1455_ _0382_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__a21bo_1
X_1386_ Inst_RegFile_32x4.mem\[6\]\[3\] Inst_RegFile_32x4.mem\[7\]\[3\] net612 VGND
+ VGND VPWR VPWR _0320_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2007_ _1030_ _0848_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__nor2_1
XFILLER_82_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2909_ net75 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1240_ net416 _0175_ _0177_ _0181_ net393 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__o311a_1
XFILLER_49_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1171_ Inst_RegFile_32x4.mem\[8\]\[0\] Inst_RegFile_32x4.mem\[9\]\[0\] net616 VGND
+ VGND VPWR VPWR _1063_ sky130_fd_sc_hd__mux2_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_0_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_0_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_64_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_16 EE4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 FrameStrobe[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2625_ net40 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput167 net167 VGND VGND VPWR VPWR E6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput145 net145 VGND VGND VPWR VPWR E2BEG[1] sky130_fd_sc_hd__buf_8
Xoutput156 net156 VGND VGND VPWR VPWR E2BEGb[4] sky130_fd_sc_hd__buf_2
X_2556_ net34 net713 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput189 net189 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
X_1507_ net397 _0424_ _0432_ _0428_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__o22a_1
X_2487_ net29 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput178 net178 VGND VGND VPWR VPWR EE4BEG[15] sky130_fd_sc_hd__buf_6
X_1438_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q _0366_ Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q
+ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__o21ai_1
X_1369_ _0299_ _0302_ net664 VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_1
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3039_ WW4END[14] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_38_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 FrameData[18] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xinput14 E2MID[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
Xinput25 EE4END[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
Xinput47 FrameData[29] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
Xinput69 N2END[7] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
Xinput58 N1END[0] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_4
X_2410_ net756 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2341_ net44 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2272_ clknet_4_5_0_UserCLK_regs _0030_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1223_ net99 net127 Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q VGND VGND VPWR VPWR
+ _0165_ sky130_fd_sc_hd__mux2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1154_ net691 net671 net657 net652 Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q
+ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__mux4_2
XFILLER_37_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1085_ net17 VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__inv_1
XFILLER_52_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1987_ net78 net110 Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q VGND VGND VPWR VPWR
+ _0841_ sky130_fd_sc_hd__mux2_1
X_2608_ net753 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2539_ net755 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2890_ FrameStrobe[18] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_1
X_1910_ Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q _0792_ VGND VGND VPWR VPWR _0793_
+ sky130_fd_sc_hd__nand2_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1841_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q _1045_ _0731_ Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__a211o_1
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1772_ _0669_ _0670_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q VGND VGND VPWR VPWR
+ _0671_ sky130_fd_sc_hd__mux2_1
X_2324_ net748 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2255_ clknet_4_13_0_UserCLK_regs _0013_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[27\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1206_ net21 net94 net106 net122 Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__mux4_1
X_2186_ _0927_ _0930_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__nor2_8
X_1137_ Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2040_ _1025_ _0893_ _0892_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q VGND VGND
+ VPWR VPWR _0894_ sky130_fd_sc_hd__o211a_1
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2942_ Inst_RegFile_switch_matrix.NN4BEG2 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__buf_4
X_2873_ net730 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_2
X_1824_ Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q _0698_ Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q
+ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__o21ai_1
X_1755_ net6 net91 net781 net119 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__mux4_1
X_1686_ net92 net108 net111 net120 Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q
+ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__mux4_1
XFILLER_85_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2307_ clknet_4_7_0_UserCLK_regs _0065_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2238_ net608 net479 _0967_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_2
XFILLER_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2169_ net499 net631 _0952_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_0_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1540_ Inst_RegFile_32x4.mem\[6\]\[1\] Inst_RegFile_32x4.mem\[7\]\[1\] net620 VGND
+ VGND VPWR VPWR _0464_ sky130_fd_sc_hd__mux2_1
XFILLER_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1471_ _0370_ _0397_ net644 VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux2_1
XFILLER_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2023_ Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q _0876_ VGND VGND VPWR VPWR _0877_
+ sky130_fd_sc_hd__nor2_1
XFILLER_62_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2925_ Inst_RegFile_switch_matrix.N4BEG1 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__buf_1
X_2856_ net773 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_13_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1807_ _0701_ _0702_ Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q _0703_ VGND VGND
+ VPWR VPWR _0704_ sky130_fd_sc_hd__o22a_1
X_2787_ clknet_4_5_0_UserCLK_regs _0123_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1738_ net91 net119 net107 net136 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux4_1
X_1669_ net781 net93 net112 net121 Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__mux4_1
Xfanout702 net706 VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__clkbuf_2
Xfanout713 net714 VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__clkbuf_2
Xfanout724 net726 VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout757 net48 VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__buf_4
Xfanout735 net57 VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__buf_2
Xfanout746 FrameStrobe[0] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__buf_1
XFILLER_85_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout768 net39 VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__clkbuf_4
Xfanout779 net28 VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__buf_4
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2710_ net28 net744 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2641_ net752 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2572_ net780 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput305 net305 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput316 net316 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__buf_6
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput349 net349 VGND VGND VPWR VPWR W2BEG[0] sky130_fd_sc_hd__buf_8
Xoutput327 net327 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput338 net338 VGND VGND VPWR VPWR SS4BEG[4] sky130_fd_sc_hd__buf_2
X_1523_ _0443_ _0446_ net645 VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__mux2_4
XFILLER_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1454_ net648 net683 net667 net447 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux4_2
X_1385_ _0318_ net675 VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__nand2b_1
XFILLER_82_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2006_ _0970_ _0974_ _0989_ net435 Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q
+ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_53_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2908_ net74 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_1
X_2839_ Inst_RegFile_switch_matrix.EE4BEG3 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1170_ _1043_ _1046_ _1059_ _1061_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__a22oi_2
XFILLER_64_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_17 EE4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 FrameStrobe[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2624_ net39 net722 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput168 net168 VGND VGND VPWR VPWR E6BEG[6] sky130_fd_sc_hd__buf_2
X_2555_ net774 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput157 net157 VGND VGND VPWR VPWR E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput146 net146 VGND VGND VPWR VPWR E2BEG[2] sky130_fd_sc_hd__buf_8
X_1506_ net417 _0431_ _0393_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__a21o_1
X_2486_ net28 net706 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput179 net179 VGND VGND VPWR VPWR EE4BEG[1] sky130_fd_sc_hd__buf_2
X_1437_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__inv_2
X_1368_ _0300_ _0301_ net679 VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__mux2_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1299_ Inst_RegFile_32x4.mem\[2\]\[1\] Inst_RegFile_32x4.mem\[3\]\[1\] net614 VGND
+ VGND VPWR VPWR _0237_ sky130_fd_sc_hd__mux2_1
XFILLER_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3038_ WW4END[13] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_38_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput37 FrameData[19] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 E2MID[2] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
Xinput26 EE4END[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_6
Xinput59 N1END[1] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_12
Xinput48 FrameData[2] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
X_2340_ net43 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2271_ clknet_4_7_0_UserCLK_regs _0029_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1222_ net71 net14 Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q VGND VGND VPWR VPWR
+ _0164_ sky130_fd_sc_hd__mux2_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1153_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q _1045_ Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q
+ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__a21oi_1
X_1084_ Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__inv_2
XFILLER_52_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1986_ Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q Inst_RegFile_switch_matrix.JW2BEG2
+ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__a21o_1
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2607_ net754 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2538_ net756 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_75_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2469_ net763 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1840_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q net640 VGND VGND VPWR VPWR _0731_
+ sky130_fd_sc_hd__nor2_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1771_ net23 net781 net91 net119 Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q
+ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__mux4_1
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2323_ net749 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2254_ clknet_4_14_0_UserCLK_regs _0012_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[27\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1205_ net60 net66 net85 net9 Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__mux4_1
X_2185_ net600 net563 _0955_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__mux2_4
X_1136_ Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__inv_2
XFILLER_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1969_ net62 net690 net81 net428 Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N4BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_68_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2872_ net746 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_2
X_1823_ _0715_ _0716_ Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.WW4BEG1 sky130_fd_sc_hd__mux2_4
X_1754_ net61 net63 net79 net82 Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q
+ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux4_1
XFILLER_7_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1685_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q _0594_ VGND VGND VPWR VPWR _0595_
+ sky130_fd_sc_hd__nor2_1
X_2306_ clknet_4_6_0_UserCLK_regs _0064_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2237_ _0939_ _0886_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__nand2_4
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2168_ net473 net607 _0952_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_0_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__inv_2
X_2099_ _0932_ _0854_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__nor2_8
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1470_ _0395_ _0396_ net687 VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2022_ Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q _0873_ _0875_ Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q
+ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__o211a_1
XFILLER_35_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2924_ Inst_RegFile_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_6
X_2855_ net33 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_28_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1806_ net683 net636 net667 net447 Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__mux4_2
X_2786_ clknet_4_5_0_UserCLK_regs _0122_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1737_ _0638_ _0639_ Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q VGND VGND VPWR VPWR
+ _0640_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1668_ net59 net65 net81 net8 Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__mux4_1
Xfanout714 FrameStrobe[5] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__buf_2
Xfanout703 net704 VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__buf_2
Xfanout725 net726 VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__clkbuf_2
Xfanout736 net737 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__clkbuf_2
X_1599_ Inst_RegFile_32x4.mem\[15\]\[2\] net622 net685 VGND VGND VPWR VPWR _0519_
+ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_5_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout758 net47 VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__buf_4
Xfanout747 net56 VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__buf_4
XFILLER_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout769 net38 VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__buf_4
XFILLER_73_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_107 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 Inst_RegFile_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_129 net139 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2640_ net753 net723 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput306 net306 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput317 net317 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__buf_8
X_2571_ net755 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_73_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput328 net328 VGND VGND VPWR VPWR SS4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput339 net339 VGND VGND VPWR VPWR SS4BEG[5] sky130_fd_sc_hd__buf_2
X_1522_ _0444_ _0445_ _0343_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux2_4
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1453_ Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q _0380_ VGND VGND VPWR VPWR _0381_
+ sky130_fd_sc_hd__and2b_1
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1384_ Inst_RegFile_32x4.mem\[4\]\[3\] Inst_RegFile_32x4.mem\[5\]\[3\] net612 VGND
+ VGND VPWR VPWR _0318_ sky130_fd_sc_hd__mux2_1
XFILLER_82_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2005_ _1031_ _0856_ _0858_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2907_ net73 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_61_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2838_ Inst_RegFile_switch_matrix.EE4BEG2 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_4
X_2769_ clknet_4_2_0_UserCLK_regs _0105_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_18 EE4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2623_ net770 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2554_ net775 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1505_ _0430_ _0429_ net686 VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
Xoutput147 net147 VGND VGND VPWR VPWR E2BEG[3] sky130_fd_sc_hd__buf_6
Xoutput158 net158 VGND VGND VPWR VPWR E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput169 net169 VGND VGND VPWR VPWR E6BEG[7] sky130_fd_sc_hd__buf_2
X_2485_ net747 net705 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1436_ net83 net10 net95 net123 Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q
+ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux4_1
X_1367_ Inst_RegFile_32x4.mem\[20\]\[3\] Inst_RegFile_32x4.mem\[21\]\[3\] net617 VGND
+ VGND VPWR VPWR _0301_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1298_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__inv_2
X_3037_ WW4END[12] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__buf_2
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput16 E2MID[3] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 FrameData[0] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput49 FrameData[30] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
Xinput38 FrameData[1] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2270_ clknet_4_4_0_UserCLK_regs _0028_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1221_ _0986_ _0987_ _1003_ _0162_ Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q
+ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__mux4_1
XFILLER_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1152_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__clkinv_2
X_1083_ Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__inv_1
XFILLER_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1985_ _0991_ Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q
+ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__o21ai_1
X_2606_ net757 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2537_ net758 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2468_ net764 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1419_ net89 net97 net111 net115 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__mux4_1
X_2399_ net37 net742 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1770_ net63 net79 net783 net6 Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q
+ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__mux4_1
XFILLER_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2322_ net751 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2253_ clknet_4_15_0_UserCLK_regs _0011_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[26\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1204_ _0146_ _0147_ Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q VGND VGND VPWR VPWR
+ _0148_ sky130_fd_sc_hd__mux2_4
X_2184_ net630 net540 _0955_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__mux2_4
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1135_ Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__inv_2
XFILLER_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1968_ net63 net78 net691 net639 Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q
+ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.N4BEG3 sky130_fd_sc_hd__mux4_1
X_1899_ _1010_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__a211o_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone1 _0169_ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__buf_6
XFILLER_56_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2871_ net755 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1822_ net634 _0682_ _0683_ _0140_ Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q
+ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__mux4_2
X_1753_ _0653_ _1019_ Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR VPWR
+ _0654_ sky130_fd_sc_hd__o21a_1
X_1684_ net58 net7 net64 net782 Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q
+ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__mux4_1
XFILLER_85_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2305_ clknet_4_15_0_UserCLK_regs _0063_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[18\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2236_ net601 net570 _0966_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_4
X_2167_ net452 net610 _0952_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_4
X_1118_ Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_0_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ _0846_ _0838_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__nand2b_4
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2021_ Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q _0874_ VGND VGND VPWR VPWR _0875_
+ sky130_fd_sc_hd__nand2_1
XFILLER_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2923_ N4END[15] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_1
X_2854_ net32 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_13_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2785_ clknet_4_7_0_UserCLK_regs _0121_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1805_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0699_ Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q
+ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__a21bo_1
X_1736_ net680 net633 net665 net638 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__mux4_2
XFILLER_7_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1667_ _0577_ _0578_ Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR VPWR
+ _0579_ sky130_fd_sc_hd__mux2_4
X_1598_ net622 Inst_RegFile_32x4.mem\[14\]\[2\] VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__and2b_1
Xfanout715 net718 VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__buf_2
Xfanout704 net705 VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__clkbuf_2
Xfanout726 FrameStrobe[2] VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout737 net738 VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__buf_2
Xfanout748 net55 VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__buf_4
Xfanout759 net46 VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__buf_4
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2219_ net605 net512 _0963_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_4
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_108 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 Inst_RegFile_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput307 net307 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__buf_2
X_2570_ net756 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput318 net318 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__buf_4
Xoutput329 net329 VGND VGND VPWR VPWR SS4BEG[10] sky130_fd_sc_hd__buf_2
X_1521_ Inst_RegFile_32x4.mem\[22\]\[1\] Inst_RegFile_32x4.mem\[23\]\[1\] net626 VGND
+ VGND VPWR VPWR _0445_ sky130_fd_sc_hd__mux2_1
XFILLER_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1452_ net137 net672 net658 net654 Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux4_2
X_1383_ net663 _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__nand2b_1
XFILLER_67_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2004_ Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q Inst_RegFile_switch_matrix.JN2BEG0
+ _0857_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__a21o_1
XFILLER_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2906_ net72 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_61_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2768_ clknet_4_0_0_UserCLK_regs _0104_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1719_ _0624_ _0623_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q VGND VGND VPWR VPWR
+ _0625_ sky130_fd_sc_hd__mux2_1
X_2699_ net50 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_19 EE4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2622_ net771 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2553_ net776 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1504_ Inst_RegFile_32x4.mem\[4\]\[0\] Inst_RegFile_32x4.mem\[5\]\[0\] net432 VGND
+ VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux2_1
Xoutput148 Inst_RegFile_switch_matrix.E2BEG4 VGND VGND VPWR VPWR E2BEG[4] sky130_fd_sc_hd__buf_8
Xoutput159 net159 VGND VGND VPWR VPWR E2BEGb[7] sky130_fd_sc_hd__buf_2
X_2484_ net748 net705 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1435_ Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q _0363_ _0362_ Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q
+ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__o211a_1
X_1366_ Inst_RegFile_32x4.mem\[22\]\[3\] Inst_RegFile_32x4.mem\[23\]\[3\] net617 VGND
+ VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3036_ WW4END[11] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__buf_4
X_1297_ Inst_RegFile_32x4.mem\[0\]\[1\] Inst_RegFile_32x4.mem\[1\]\[1\] net616 VGND
+ VGND VPWR VPWR _0235_ sky130_fd_sc_hd__mux2_1
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput28 FrameData[10] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
Xinput17 E2MID[4] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
Xinput39 FrameData[20] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1220_ _0162_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JW2BEG5 sky130_fd_sc_hd__inv_2
XFILLER_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1151_ net73 net16 net101 net129 Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q
+ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__mux4_2
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1082_ Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__inv_2
XFILLER_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1984_ _0835_ _0837_ Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q _0833_ VGND VGND VPWR
+ VPWR _0838_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2605_ net769 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2536_ net759 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2467_ net765 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1418_ net61 net69 net783 net12 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__mux4_1
XFILLER_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2398_ net36 net742 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1349_ Inst_RegFile_32x4.mem\[22\]\[2\] Inst_RegFile_32x4.mem\[23\]\[2\] net617 VGND
+ VGND VPWR VPWR _0285_ sky130_fd_sc_hd__mux2_1
XFILLER_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3019_ W6END[4] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_34_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2321_ net752 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2252_ clknet_4_12_0_UserCLK_regs _0010_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[26\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1203_ net681 net634 net406 net639 Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q
+ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__mux4_2
XFILLER_65_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2183_ net604 net553 _0955_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__mux2_4
X_1134_ Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__inv_2
XFILLER_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1967_ net647 Inst_RegFile_switch_matrix.JN2BEG3 _0829_ _0828_ Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E1BEG0
+ sky130_fd_sc_hd__mux4_2
X_1898_ net58 Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR _0783_
+ sky130_fd_sc_hd__nor2_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2519_ net778 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
Xclone2 net395 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__buf_6
XFILLER_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2870_ net49 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_4_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1821_ net61 net89 net692 net419 Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q
+ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__mux4_1
X_1752_ net680 net427 net665 net638 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__mux4_2
X_1683_ _0592_ _1009_ Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q VGND VGND VPWR VPWR
+ _0593_ sky130_fd_sc_hd__o21ai_2
XFILLER_85_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2304_ clknet_4_15_0_UserCLK_regs _0062_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[18\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2235_ net629 net508 _0966_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__mux2_4
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2166_ _0944_ _0887_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__nor2_8
X_1117_ Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__inv_1
XFILLER_80_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2097_ net600 net522 _0931_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__mux2_4
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2020_ net105 net133 Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q VGND VGND VPWR VPWR
+ _0874_ sky130_fd_sc_hd__mux2_1
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2922_ N4END[14] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2853_ net776 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_4
X_2784_ clknet_4_4_0_UserCLK_regs _0120_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1804_ Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q _0700_ VGND VGND VPWR VPWR _0701_
+ sky130_fd_sc_hd__and2b_1
X_1735_ net690 net652 net415 net646 Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q
+ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__mux4_1
X_1666_ net680 net633 net666 net638 Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q
+ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__mux4_2
X_1597_ net643 _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__and2b_1
Xfanout705 net706 VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__clkbuf_2
Xfanout716 net717 VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__clkbuf_2
Xfanout749 net750 VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 net57 VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkbuf_2
Xfanout727 net730 VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__buf_2
XFILLER_73_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2218_ net609 net477 _0963_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_4
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_109 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2149_ net629 net579 _0948_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__mux2_4
XFILLER_81_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput308 net308 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput319 net319 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_58_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1520_ Inst_RegFile_32x4.mem\[20\]\[1\] Inst_RegFile_32x4.mem\[21\]\[1\] net627 VGND
+ VGND VPWR VPWR _0444_ sky130_fd_sc_hd__mux2_1
XFILLER_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1451_ _0377_ _0378_ _0985_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux2_2
X_1382_ _0314_ _0315_ net676 VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
X_2003_ _1030_ _0378_ Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q VGND VGND VPWR VPWR
+ _0857_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_18_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2905_ net71 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_61_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2836_ Inst_RegFile_switch_matrix.EE4BEG0 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_4
X_2767_ clknet_4_2_0_UserCLK_regs _0103_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2698_ net49 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1718_ net58 net1 net62 net5 Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q
+ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__mux4_1
X_1649_ _0562_ _0563_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q VGND VGND VPWR VPWR
+ _0564_ sky130_fd_sc_hd__mux2_1
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2621_ net772 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2552_ net777 net712 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1503_ Inst_RegFile_32x4.mem\[6\]\[0\] Inst_RegFile_32x4.mem\[7\]\[0\] net432 VGND
+ VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
Xoutput149 net149 VGND VGND VPWR VPWR E2BEG[5] sky130_fd_sc_hd__clkbuf_4
X_2483_ net749 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1434_ net22 net107 Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q VGND VGND VPWR VPWR
+ _0363_ sky130_fd_sc_hd__mux2_1
X_1365_ _0298_ _0297_ net678 VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3035_ WW4END[10] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__buf_4
X_1296_ _0233_ _0229_ net651 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__nor3_2
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2819_ E6END[9] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 E2MID[5] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
Xinput29 FrameData[11] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1150_ _1039_ _1040_ _1042_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q VGND VGND
+ VPWR VPWR _1043_ sky130_fd_sc_hd__a211o_1
XFILLER_77_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1081_ Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__inv_2
XFILLER_60_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1983_ _1029_ _0836_ Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q VGND VGND VPWR VPWR
+ _0837_ sky130_fd_sc_hd__a21o_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2604_ net780 net719 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2535_ net760 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2466_ net766 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1417_ _0347_ _0981_ Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q VGND VGND VPWR VPWR
+ _0348_ sky130_fd_sc_hd__o21a_1
XFILLER_68_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2397_ net35 net742 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1348_ _0283_ _0282_ net678 VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_1
XFILLER_28_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1279_ Inst_RegFile_32x4.mem\[18\]\[0\] Inst_RegFile_32x4.mem\[19\]\[0\] net618 VGND
+ VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_1
XFILLER_83_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3018_ W6END[3] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_34_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2320_ net753 net733 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2251_ clknet_4_13_0_UserCLK_regs _0009_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[26\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1202_ net691 net414 net415 net653 Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q
+ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux4_2
X_2182_ net609 net557 _0955_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__mux2_4
X_1133_ Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__inv_2
XFILLER_80_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1966_ net682 _0563_ Inst_RegFile_switch_matrix.JN2BEG0 net396 Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E1BEG1
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_31_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1897_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q _1045_ Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q
+ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__a211o_1
X_2518_ net779 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2449_ net53 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone3 _0564_ _0561_ Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q VGND VGND VPWR VPWR
+ net395 sky130_fd_sc_hd__mux2_4
XFILLER_56_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1820_ Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q _0714_ _0713_ VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.WW4BEG2 sky130_fd_sc_hd__o21ba_1
X_1751_ Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q _0651_ VGND VGND VPWR VPWR _0652_
+ sky130_fd_sc_hd__or2_1
X_1682_ net680 net427 net665 net638 Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q
+ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__mux4_2
X_2303_ clknet_4_15_0_UserCLK_regs _0061_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[18\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2234_ net605 net547 _0966_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__mux2_4
X_2165_ net601 net530 _0951_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux2_2
XFILLER_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1116_ net1 VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__inv_2
XFILLER_53_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2096_ net630 net475 _0931_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__mux2_4
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1949_ net85 net109 net136 Inst_RegFile_switch_matrix.JN2BEG1 Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_8_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2921_ N4END[13] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_1
XFILLER_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2852_ net777 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_4
X_2783_ clknet_4_5_0_UserCLK_regs _0119_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1803_ _0697_ _0698_ Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q VGND VGND VPWR VPWR
+ _0700_ sky130_fd_sc_hd__mux2_1
X_1734_ _0637_ _0634_ Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JS2BEG7 sky130_fd_sc_hd__mux2_4
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1665_ net690 net670 net657 net646 Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__mux4_1
X_1596_ _0514_ _0515_ net685 VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__mux2_1
Xfanout706 FrameStrobe[7] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__clkbuf_2
Xfanout717 net718 VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__buf_2
Xfanout728 net729 VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__clkbuf_2
Xfanout739 FrameStrobe[10] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__buf_2
XFILLER_85_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2217_ _0886_ _0937_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__nand2_8
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2148_ net604 net558 _0948_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux2_4
XFILLER_53_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2079_ _0924_ _0855_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__nor2_8
XFILLER_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput309 net309 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__buf_2
XFILLER_4_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1450_ net63 net91 net26 net119 Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q
+ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__mux4_2
XFILLER_4_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1381_ Inst_RegFile_32x4.mem\[0\]\[3\] Inst_RegFile_32x4.mem\[1\]\[3\] net615 VGND
+ VGND VPWR VPWR _0315_ sky130_fd_sc_hd__mux2_1
XFILLER_67_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2002_ Inst_RegFile_switch_matrix.JW2BEG0 Inst_RegFile_switch_matrix.JS2BEG0 _1030_
+ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__mux2_1
XFILLER_35_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2904_ net70 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_61_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2835_ EE4END[15] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_1
X_2766_ clknet_4_0_0_UserCLK_regs _0102_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2697_ net758 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1717_ net86 net90 net88 net114 Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q
+ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__mux4_1
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1648_ net77 net20 net105 net133 Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q
+ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__mux4_2
X_1579_ Inst_RegFile_32x4.mem\[26\]\[2\] Inst_RegFile_32x4.mem\[27\]\[2\] net628 VGND
+ VGND VPWR VPWR _0499_ sky130_fd_sc_hd__mux2_1
XFILLER_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer41 _1072_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__buf_6
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2620_ net773 net721 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2551_ net29 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1502_ net417 _0427_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__and2b_1
X_2482_ net751 net702 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1433_ Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q Inst_RegFile_switch_matrix.JS2BEG4
+ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a21o_1
X_1364_ Inst_RegFile_32x4.mem\[18\]\[3\] Inst_RegFile_32x4.mem\[19\]\[3\] net617 VGND
+ VGND VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
X_1295_ net446 _0230_ _0232_ net662 VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3034_ WW4END[9] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__buf_4
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2818_ E6END[8] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_1
X_2749_ clknet_4_13_0_UserCLK_regs _0085_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[31\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_7_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput19 E2MID[6] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1080_ net128 VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__inv_1
XFILLER_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1982_ net62 net90 Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q VGND VGND VPWR VPWR
+ _0836_ sky130_fd_sc_hd__mux2_1
XFILLER_60_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2603_ net50 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2534_ net762 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2465_ net40 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1416_ net650 net684 net431 net642 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__mux4_2
X_2396_ net773 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1347_ Inst_RegFile_32x4.mem\[18\]\[2\] Inst_RegFile_32x4.mem\[19\]\[2\] net618 VGND
+ VGND VPWR VPWR _0283_ sky130_fd_sc_hd__mux2_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1278_ Inst_RegFile_32x4.mem\[16\]\[0\] Inst_RegFile_32x4.mem\[17\]\[0\] net618 VGND
+ VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux2_1
X_3017_ W6END[2] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2250_ clknet_4_12_0_UserCLK_regs _0008_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[26\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1201_ net416 _0144_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__nand2b_1
XFILLER_77_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2181_ _0920_ _0929_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__nand2_8
X_1132_ Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__inv_1
XFILLER_80_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1965_ net406 net689 Inst_RegFile_switch_matrix.JN2BEG1 _0377_ Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E1BEG2
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_31_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1896_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q net404 VGND VGND VPWR VPWR _0781_
+ sky130_fd_sc_hd__nor2_4
X_2517_ net747 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2448_ net52 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2379_ net755 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_71_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1750_ net690 net407 net415 net647 Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q
+ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__mux4_1
XFILLER_30_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1681_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q _0590_ VGND VGND VPWR VPWR _0591_
+ sky130_fd_sc_hd__nor2_1
X_2302_ clknet_4_11_0_UserCLK_regs _0060_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[18\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2233_ net608 net510 _0966_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__mux2_4
XFILLER_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2164_ net629 net517 _0951_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__mux2_4
X_1115_ Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__inv_2
X_2095_ net604 net483 _0931_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__mux2_4
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2997_ Inst_RegFile_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__buf_6
X_1948_ Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q _0826_ _0825_ VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.NN4BEG0 sky130_fd_sc_hd__o21ba_4
X_1879_ _1044_ net689 Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _0766_ sky130_fd_sc_hd__mux2_1
XFILLER_79_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2920_ N4END[12] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2851_ net778 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2782_ clknet_4_5_0_UserCLK_regs _0118_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1802_ _1044_ net689 Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q VGND VGND VPWR VPWR
+ _0699_ sky130_fd_sc_hd__mux2_1
X_1733_ _0636_ _0635_ Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR VPWR
+ _0637_ sky130_fd_sc_hd__mux2_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1664_ _0576_ _0573_ Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JS2BEG2 sky130_fd_sc_hd__mux2_4
X_1595_ Inst_RegFile_32x4.mem\[10\]\[2\] Inst_RegFile_32x4.mem\[11\]\[2\] net623 VGND
+ VGND VPWR VPWR _0515_ sky130_fd_sc_hd__mux2_1
Xfanout718 FrameStrobe[4] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__buf_2
Xfanout707 net708 VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__buf_2
Xfanout729 net730 VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__buf_2
X_2216_ net600 net535 _0962_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__mux2_4
XFILLER_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2147_ net608 net516 _0948_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__mux2_4
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2078_ _0885_ _0879_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_64_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1380_ Inst_RegFile_32x4.mem\[2\]\[3\] Inst_RegFile_32x4.mem\[3\]\[3\] net614 VGND
+ VGND VPWR VPWR _0314_ sky130_fd_sc_hd__mux2_1
X_2001_ net437 _0847_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_18_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2903_ Inst_RegFile_switch_matrix.JN2BEG7 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_61_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2834_ EE4END[14] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_1
X_2765_ clknet_4_2_0_UserCLK_regs _0101_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1716_ _0620_ _0621_ Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q VGND VGND VPWR VPWR
+ _0622_ sky130_fd_sc_hd__mux2_2
X_2696_ net759 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1647_ net76 net19 net132 Inst_RegFile_switch_matrix.JN2BEG5 Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__mux4_1
X_1578_ Inst_RegFile_32x4.BD_comb\[3\] Inst_RegFile_32x4.BD_reg\[3\] Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q
+ VGND VGND VPWR VPWR BD3 sky130_fd_sc_hd__mux2_4
XFILLER_58_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer20 BD3 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__buf_6
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer42 net433 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_15_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2550_ net28 net711 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1501_ _0426_ _0425_ net687 VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux2_1
X_2481_ net53 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1432_ Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q _0984_ Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q
+ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__o21ai_1
X_1363_ Inst_RegFile_32x4.mem\[16\]\[3\] Inst_RegFile_32x4.mem\[17\]\[3\] net617 VGND
+ VGND VPWR VPWR _0297_ sky130_fd_sc_hd__mux2_1
X_1294_ _0231_ net445 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_66_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3033_ WW4END[8] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__buf_4
XFILLER_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2817_ E6END[7] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_1
X_2748_ clknet_4_13_0_UserCLK_regs _0084_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[31\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_52_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2679_ net778 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1981_ _1028_ _0128_ _0834_ Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q VGND VGND VPWR
+ VPWR _0835_ sky130_fd_sc_hd__o211a_1
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2602_ net49 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2533_ net763 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2464_ net768 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1415_ Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q _0345_ VGND VGND VPWR VPWR _0346_
+ sky130_fd_sc_hd__or2_1
X_2395_ net33 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1346_ Inst_RegFile_32x4.mem\[16\]\[2\] Inst_RegFile_32x4.mem\[17\]\[2\] net618 VGND
+ VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_1
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1277_ _0213_ _0216_ net663 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__mux2_1
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3016_ net133 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1200_ _0143_ _1063_ net444 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__mux2_1
X_2180_ net569 net602 _0954_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__mux2_4
X_1131_ Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_48_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1964_ net635 _0407_ Inst_RegFile_switch_matrix.JN2BEG2 _0827_ Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E1BEG3
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_31_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1895_ Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q _0779_ VGND VGND VPWR VPWR _0780_
+ sky130_fd_sc_hd__nand2_1
X_2516_ net55 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2447_ net754 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2378_ net756 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_39_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1329_ _0264_ _0263_ net676 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__mux2_4
XFILLER_71_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput290 net290 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1680_ net691 net414 net407 net646 Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q
+ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__mux4_1
X_2301_ clknet_4_11_0_UserCLK_regs _0059_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[16\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2232_ _0926_ _0937_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__nand2_8
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2163_ net605 net518 _0951_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux2_2
X_1114_ Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__inv_1
X_2094_ net609 net488 _0931_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__mux2_4
XFILLER_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2996_ clknet_1_0__leaf_UserCLK VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__buf_2
X_1947_ net60 net784 net693 net660 Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q
+ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__mux4_2
X_1878_ _0762_ _0763_ _0764_ Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q VGND VGND
+ VPWR VPWR _0765_ sky130_fd_sc_hd__o22a_1
XFILLER_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2850_ net779 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
X_1801_ net73 net16 net101 net129 Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q
+ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__mux4_2
X_2781_ clknet_4_7_0_UserCLK_regs _0117_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1732_ net58 net1 net62 net5 Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q
+ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__mux4_1
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1663_ _0574_ _0575_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q VGND VGND VPWR VPWR
+ _0576_ sky130_fd_sc_hd__mux2_1
X_1594_ Inst_RegFile_32x4.mem\[8\]\[2\] Inst_RegFile_32x4.mem\[9\]\[2\] net623 VGND
+ VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux2_1
Xfanout708 net709 VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__clkbuf_2
Xfanout719 FrameStrobe[3] VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2215_ net630 net491 _0962_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__mux2_4
XFILLER_81_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2146_ _0926_ _0939_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__nand2_8
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2077_ _0885_ _0879_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nor2_8
XFILLER_53_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2979_ Inst_RegFile_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2000_ Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q _0852_ _0850_ VGND VGND VPWR VPWR
+ _0854_ sky130_fd_sc_hd__a21o_4
XFILLER_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2833_ EE4END[13] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
X_2764_ clknet_4_0_0_UserCLK_regs _0100_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1715_ net649 net684 net668 net637 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__mux4_1
X_2695_ net45 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1646_ _0559_ _0560_ Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q VGND VGND VPWR VPWR
+ _0561_ sky130_fd_sc_hd__mux2_4
X_1577_ _0498_ _0483_ _0409_ VGND VGND VPWR VPWR Inst_RegFile_32x4.BD_comb\[3\] sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_69_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer10 _0352_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer43 _0334_ VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__buf_6
X_2129_ net575 net602 _0943_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_52_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1500_ Inst_RegFile_32x4.mem\[0\]\[0\] Inst_RegFile_32x4.mem\[1\]\[0\] net624 VGND
+ VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
X_2480_ net52 net703 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1431_ _0360_ _0357_ Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JS2BEG4 sky130_fd_sc_hd__mux2_4
X_1362_ _0292_ _0295_ net664 VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__mux2_1
X_1293_ Inst_RegFile_32x4.mem\[12\]\[1\] Inst_RegFile_32x4.mem\[13\]\[1\] net612 VGND
+ VGND VPWR VPWR _0231_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3032_ WW4END[7] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__buf_4
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2816_ E6END[6] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2747_ clknet_4_9_0_UserCLK_regs _0083_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[29\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2678_ net779 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1629_ Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q _0543_ _0545_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q
+ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__a211o_1
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ _1039_ _1040_ _1042_ Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q VGND VGND VPWR
+ VPWR _0834_ sky130_fd_sc_hd__a211o_1
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2601_ net758 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2532_ net764 net710 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2463_ net770 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1414_ net692 net674 net660 net656 Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__mux4_1
X_2394_ net32 net742 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1345_ _0277_ _0280_ net663 VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
XFILLER_83_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1276_ _0214_ _0215_ net446 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__mux2_1
X_3015_ net132 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_3_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_69_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1130_ Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_48_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1963_ net682 Inst_RegFile_switch_matrix.E2BEG3 _0829_ _0828_ Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S1BEG0
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_31_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1894_ net689 _0778_ Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _0779_ sky130_fd_sc_hd__mux2_1
X_2515_ net749 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2446_ net757 net698 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2377_ net758 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_39_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1328_ Inst_RegFile_32x4.mem\[14\]\[2\] Inst_RegFile_32x4.mem\[15\]\[2\] net614 VGND
+ VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux2_1
XFILLER_56_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1259_ _0198_ _0199_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q VGND VGND VPWR VPWR
+ _0200_ sky130_fd_sc_hd__mux2_1
Xclone6 BD2 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__buf_6
XFILLER_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput280 Inst_RegFile_switch_matrix.NN4BEG1 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__buf_8
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput291 net291 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2300_ clknet_4_14_0_UserCLK_regs _0058_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[16\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2231_ net601 net468 _0965_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__mux2_4
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2162_ net609 net524 _0951_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux2_4
X_2093_ _0886_ _0929_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__nand2_8
X_1113_ Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__inv_1
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2995_ Inst_RegFile_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__buf_6
X_1946_ Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q _0824_ _0822_ Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q
+ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__o211a_1
X_1877_ net82 net110 net783 net692 Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q
+ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__mux4_1
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2429_ net772 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_76_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1800_ net73 net16 net101 net129 Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q
+ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux4_2
X_2780_ clknet_4_4_0_UserCLK_regs _0116_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1731_ net86 net90 net110 net114 Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__mux4_1
XFILLER_7_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1662_ net781 net93 net109 net121 Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q
+ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__mux4_1
X_1593_ _0505_ _0512_ _0394_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__mux2_4
Xfanout709 net710 VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__clkbuf_2
X_2214_ net604 net509 _0962_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__mux2_4
X_2145_ net600 net514 _0947_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__mux2_4
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2076_ net571 net602 _0922_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__mux2_4
XFILLER_81_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2978_ Inst_RegFile_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_6
X_1929_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q net404 VGND VGND VPWR VPWR _0810_
+ sky130_fd_sc_hd__nor2_1
XFILLER_1_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold90 Inst_RegFile_32x4.mem\[2\]\[1\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2901_ Inst_RegFile_switch_matrix.JN2BEG5 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__buf_1
XFILLER_50_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2832_ EE4END[12] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_1
X_2763_ clknet_4_2_0_UserCLK_regs _0099_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1714_ net136 net673 net659 net655 Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q
+ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__mux4_1
X_2694_ net761 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1645_ net81 net8 net121 Inst_RegFile_switch_matrix.JN2BEG3 Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__mux4_2
X_1576_ _0490_ _0497_ _0394_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_69_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer11 net402 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlymetal6s2s_1
X_2128_ net565 net631 _0943_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__mux2_4
Xrebuffer44 _1071_ VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_6
XFILLER_81_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2059_ _0986_ Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q VGND VGND VPWR VPWR _0910_
+ sky130_fd_sc_hd__nand2_1
XFILLER_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1430_ _0358_ _0359_ Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q VGND VGND VPWR VPWR
+ _0360_ sky130_fd_sc_hd__mux2_1
XFILLER_49_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1361_ _0293_ _0294_ net678 VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__mux2_1
X_1292_ Inst_RegFile_32x4.mem\[14\]\[1\] Inst_RegFile_32x4.mem\[15\]\[1\] A_ADR0 VGND
+ VGND VPWR VPWR _0230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3031_ WW4END[6] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_4
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2815_ E6END[5] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_1
X_2746_ clknet_4_13_0_UserCLK_regs _0082_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[29\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2677_ net747 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1628_ Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q _0544_ VGND VGND VPWR VPWR _0545_
+ sky130_fd_sc_hd__and2b_1
XFILLER_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1559_ _0479_ _0480_ net688 VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux2_1
XFILLER_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_UserCLK_regs clknet_0_UserCLK_regs VGND VGND VPWR VPWR clknet_4_11_0_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2600_ net759 net717 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2531_ net765 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2462_ net36 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2393_ net31 net742 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1413_ Inst_RegFile_32x4.mem\[26\]\[0\] Inst_RegFile_32x4.mem\[27\]\[0\] net628 VGND
+ VGND VPWR VPWR _0344_ sky130_fd_sc_hd__mux2_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1344_ _0278_ _0279_ net676 VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_1
XFILLER_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1275_ Inst_RegFile_32x4.mem\[28\]\[0\] Inst_RegFile_32x4.mem\[29\]\[0\] net615 VGND
+ VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3014_ net131 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2729_ net47 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ net666 _0563_ Inst_RegFile_switch_matrix.E2BEG0 net396 Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q
+ Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S1BEG1
+ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1893_ net85 net11 net96 net124 Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q
+ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_31_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2514_ net751 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2445_ net769 net701 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2376_ net759 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1327_ Inst_RegFile_32x4.mem\[12\]\[2\] Inst_RegFile_32x4.mem\[13\]\[2\] net614 VGND
+ VGND VPWR VPWR _0263_ sky130_fd_sc_hd__mux2_1
XFILLER_71_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1258_ net24 net87 net89 net97 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux4_1
X_1189_ _0133_ _1001_ Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q VGND VGND VPWR VPWR
+ _0134_ sky130_fd_sc_hd__o21a_1
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput270 net270 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_58_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput281 net281 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__buf_8
Xoutput292 net292 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_58_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2230_ net629 net465 _0965_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__mux2_4
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2161_ _0920_ _0933_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__nand2_4
X_2092_ _0854_ _0847_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nand2_8
X_1112_ Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_85_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2994_ Inst_RegFile_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__buf_4
X_1945_ _0823_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__inv_1
X_1876_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q _0760_ Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q
+ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2428_ net773 net695 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2359_ net29 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1730_ _0632_ _0633_ Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR VPWR
+ _0634_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_13_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1661_ net65 net8 net2 net25 Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q
+ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__mux4_1
XFILLER_7_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1592_ _0508_ _0511_ net645 VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__mux2_1
XFILLER_85_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2213_ net608 net492 _0962_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_4
X_2144_ net629 net455 _0947_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__mux2_4
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2075_ net564 net631 _0922_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_64_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2977_ Inst_RegFile_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__buf_4
X_1928_ Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q _0808_ VGND VGND VPWR VPWR _0809_
+ sky130_fd_sc_hd__nand2_1
X_1859_ Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q _0747_ _0746_ VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.SS4BEG0 sky130_fd_sc_hd__o21ba_4
XFILLER_1_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold91 Inst_RegFile_32x4.mem\[28\]\[1\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 Inst_RegFile_32x4.mem\[26\]\[2\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
X_2900_ Inst_RegFile_switch_matrix.JN2BEG4 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_26_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2831_ EE4END[11] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__buf_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2762_ clknet_4_0_0_UserCLK_regs _0098_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1713_ _0614_ _0616_ _0619_ _1016_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.JN2BEG1
+ sky130_fd_sc_hd__a22o_4
X_2693_ net763 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1644_ net69 net97 net25 net125 Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q
+ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__mux4_1
X_1575_ _0493_ _0496_ net644 VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer45 _0853_ VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__buf_12
X_2127_ net528 net606 _0943_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__mux2_4
X_2058_ net98 Inst_RegFile_switch_matrix.JW2BEG3 Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q
+ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__mux2_1
XFILLER_81_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1360_ Inst_RegFile_32x4.mem\[28\]\[3\] Inst_RegFile_32x4.mem\[29\]\[3\] net615 VGND
+ VGND VPWR VPWR _0294_ sky130_fd_sc_hd__mux2_1
X_1291_ net416 _0228_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_66_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3030_ WW4END[5] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__buf_2
XFILLER_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2814_ E6END[4] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_1
X_2745_ clknet_4_9_0_UserCLK_regs _0081_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[29\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2676_ net748 net728 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1627_ net76 net19 Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q VGND VGND VPWR VPWR
+ _0544_ sky130_fd_sc_hd__mux2_1
XFILLER_86_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1558_ Inst_RegFile_32x4.mem\[22\]\[3\] Inst_RegFile_32x4.mem\[23\]\[3\] net626 VGND
+ VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux2_1
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1489_ _0413_ _0414_ _0343_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
XFILLER_86_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2530_ net766 net709 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2461_ net772 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1412_ _0323_ _0326_ _0340_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a22o_4
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2392_ net30 net742 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_79_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1343_ Inst_RegFile_32x4.mem\[28\]\[2\] Inst_RegFile_32x4.mem\[29\]\[2\] net615 VGND
+ VGND VPWR VPWR _0279_ sky130_fd_sc_hd__mux2_1
XFILLER_83_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1274_ Inst_RegFile_32x4.mem\[30\]\[0\] Inst_RegFile_32x4.mem\[31\]\[0\] net615 VGND
+ VGND VPWR VPWR _0214_ sky130_fd_sc_hd__mux2_1
X_3013_ net130 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2728_ net759 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2659_ net42 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout690 net135 VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__buf_2
XFILLER_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1961_ net635 net689 Inst_RegFile_switch_matrix.E2BEG1 _0377_ Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S1BEG2
+ sky130_fd_sc_hd__mux4_2
X_1892_ Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q _0772_ _0774_ _0777_ VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix.EE4BEG3 sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_31_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2513_ net752 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2444_ net780 net699 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2375_ net760 net737 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1326_ _0260_ _0261_ net444 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__mux2_4
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1257_ net61 net69 net783 net12 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux4_1
XFILLER_71_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1188_ net681 net634 net406 net639 Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q
+ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__mux4_2
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput271 net271 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput260 net260 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_79_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput282 net282 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__buf_6
Xoutput293 Inst_RegFile_switch_matrix.S1BEG1 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__buf_6
XFILLER_58_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2160_ net457 net602 _0950_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__mux2_4
X_1111_ Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__inv_2
X_2091_ _0847_ _0854_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__and2_4
XFILLER_65_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2993_ Inst_RegFile_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__buf_8
X_1944_ net668 _0697_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q VGND VGND VPWR VPWR
+ _0823_ sky130_fd_sc_hd__mux2_1
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1875_ Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q _0761_ VGND VGND VPWR VPWR _0762_
+ sky130_fd_sc_hd__and2b_1
X_2427_ net774 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2358_ net779 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1309_ _0245_ _0246_ net678 VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__mux2_1
X_2289_ clknet_4_8_0_UserCLK_regs _0047_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[23\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1660_ _0571_ _0572_ Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q VGND VGND VPWR VPWR
+ _0573_ sky130_fd_sc_hd__mux2_4
X_1591_ _0509_ _0510_ net688 VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__mux2_1
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2212_ _0926_ _0958_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__nand2_8
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2143_ net604 net534 _0947_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__mux2_4
XFILLER_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2074_ net551 net606 _0922_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__mux2_4
XFILLER_81_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2976_ Inst_RegFile_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__buf_4
X_1927_ net689 _0807_ Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR
+ _0808_ sky130_fd_sc_hd__mux2_1
X_1858_ net60 net3 net693 net661 Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q
+ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__mux4_1
X_1789_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q net434 _0686_ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__o211a_1
XFILLER_1_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold81 Inst_RegFile_32x4.mem\[20\]\[1\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 Inst_RegFile_32x4.mem\[2\]\[3\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 Inst_RegFile_32x4.mem\[26\]\[1\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2830_ EE4END[10] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_26_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2761_ clknet_4_0_0_UserCLK_regs _0097_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1712_ _0617_ _0618_ Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q VGND VGND VPWR VPWR
+ _0619_ sky130_fd_sc_hd__mux2_1
X_2692_ net764 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_1 E6END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1643_ _0558_ _0555_ Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.JN2BEG3 sky130_fd_sc_hd__mux2_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1574_ _0494_ _0495_ net686 VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__mux2_1
XFILLER_58_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ net560 net610 _0943_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux2_4
X_2057_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q _0726_ _0904_ _0907_ Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q
+ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__o221a_1
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2959_ net101 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1290_ _0226_ _0227_ net444 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__mux2_1
X_2813_ E6END[3] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_1
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2744_ clknet_4_6_0_UserCLK_regs _0080_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[29\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2675_ net749 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1626_ net104 Inst_RegFile_switch_matrix.JN2BEG6 Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q
+ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__mux2_1
X_1557_ Inst_RegFile_32x4.mem\[20\]\[3\] Inst_RegFile_32x4.mem\[21\]\[3\] net626 VGND
+ VGND VPWR VPWR _0479_ sky130_fd_sc_hd__mux2_1
X_1488_ Inst_RegFile_32x4.mem\[22\]\[0\] Inst_RegFile_32x4.mem\[23\]\[0\] net626 VGND
+ VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
X_2109_ net493 net602 _0935_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__mux2_4
XFILLER_54_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer4 _0139_ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_6
XFILLER_61_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2460_ net773 net700 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_54_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1411_ Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q _0341_ Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q
+ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o21a_1
X_2391_ net778 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_79_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1342_ Inst_RegFile_32x4.mem\[30\]\[2\] Inst_RegFile_32x4.mem\[31\]\[2\] net615 VGND
+ VGND VPWR VPWR _0278_ sky130_fd_sc_hd__mux2_1
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1273_ _0211_ _0212_ net678 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_1
XFILLER_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3012_ net129 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__buf_1
XFILLER_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2727_ net760 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2658_ net41 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2589_ net772 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1609_ _0528_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__inv_1
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout680 net682 VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__buf_2
XFILLER_18_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout691 net134 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1960_ net640 _0407_ Inst_RegFile_switch_matrix.E2BEG2 _0827_ Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q
+ Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.S1BEG3
+ sky130_fd_sc_hd__mux4_2
X_1891_ Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q _0776_ Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q
+ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_31_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2512_ net753 net708 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2443_ net755 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2374_ net761 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1325_ Inst_RegFile_32x4.mem\[8\]\[2\] Inst_RegFile_32x4.mem\[9\]\[2\] net614 VGND
+ VGND VPWR VPWR _0261_ sky130_fd_sc_hd__mux2_1
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1256_ _0972_ _0196_ Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q VGND VGND VPWR VPWR
+ _0197_ sky130_fd_sc_hd__o21a_1
XFILLER_56_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1187_ _0131_ Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q VGND VGND VPWR VPWR _0132_
+ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_82_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput261 net261 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput250 Inst_RegFile_switch_matrix.JN2BEG6 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_8
XFILLER_79_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput272 net272 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput283 net283 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput294 Inst_RegFile_switch_matrix.S1BEG2 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__buf_6
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__inv_1
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2090_ net572 net602 _0928_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__mux2_4
XFILLER_80_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1943_ Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q _0821_ VGND VGND VPWR VPWR _0822_
+ sky130_fd_sc_hd__nand2_1
X_1874_ net674 net660 Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _0761_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_UserCLK UserCLK VGND VGND VPWR VPWR clknet_0_UserCLK sky130_fd_sc_hd__clkbuf_16
X_2426_ net775 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2357_ net56 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2288_ clknet_4_10_0_UserCLK_regs _0046_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[23\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1308_ Inst_RegFile_32x4.mem\[24\]\[1\] Inst_RegFile_32x4.mem\[25\]\[1\] net619 VGND
+ VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux2_1
XFILLER_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1239_ net445 _0180_ _0179_ net416 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__o211ai_1
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1590_ Inst_RegFile_32x4.mem\[22\]\[2\] Inst_RegFile_32x4.mem\[23\]\[2\] net626 VGND
+ VGND VPWR VPWR _0510_ sky130_fd_sc_hd__mux2_1
XFILLER_7_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2211_ net600 net500 _0961_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__mux2_4
XFILLER_59_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2142_ net608 net478 _0947_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__mux2_4
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2073_ net532 net610 _0922_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__mux2_4
XFILLER_81_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2975_ S4END[15] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_2
X_1926_ net64 net92 net7 net138 Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q
+ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_12_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1857_ Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q _0745_ _0743_ Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q
+ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__o211a_1
X_1788_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q net403 VGND VGND VPWR VPWR _0686_
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2409_ net758 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold60 Inst_RegFile_32x4.mem\[20\]\[0\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 Inst_RegFile_32x4.mem\[16\]\[2\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 Inst_RegFile_32x4.mem\[18\]\[1\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold93 Inst_RegFile_32x4.mem\[24\]\[2\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2760_ clknet_4_0_0_UserCLK_regs _0096_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2691_ net42 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1711_ net24 net782 net92 net120 Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q
+ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__mux4_1
XANTENNA_2 E6END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ _0556_ _0557_ Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q VGND VGND VPWR VPWR
+ _0558_ sky130_fd_sc_hd__mux2_1
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1573_ Inst_RegFile_32x4.mem\[6\]\[3\] Inst_RegFile_32x4.mem\[7\]\[3\] net620 VGND
+ VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux2_1
XFILLER_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ _0942_ _0921_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__nor2_8
X_2056_ Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q _0906_ Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__o21ai_1
Xrebuffer47 _0958_ VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__buf_8
XFILLER_81_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2958_ net100 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__buf_1
X_1909_ _0698_ _0541_ Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q VGND VGND VPWR VPWR
+ _0792_ sky130_fd_sc_hd__mux2_1
X_2889_ FrameStrobe[17] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__buf_1
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2812_ E6END[2] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_1
X_2743_ clknet_4_15_0_UserCLK_regs _0079_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[19\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2674_ net751 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1625_ _0541_ _0540_ Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR VPWR
+ _0542_ sky130_fd_sc_hd__mux2_4
X_1556_ _0476_ _0477_ net688 VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux2_1
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1487_ Inst_RegFile_32x4.mem\[20\]\[0\] Inst_RegFile_32x4.mem\[21\]\[0\] net626 VGND
+ VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2108_ net464 net630 _0935_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__mux2_4
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2039_ net105 net133 Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q VGND VGND VPWR VPWR
+ _0893_ sky130_fd_sc_hd__mux2_1
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer5 _0394_ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1410_ net65 net8 net110 net121 Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q
+ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux4_2
XFILLER_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2390_ net779 net741 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1341_ _0275_ _0276_ net678 VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__mux2_1
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1272_ Inst_RegFile_32x4.mem\[24\]\[0\] Inst_RegFile_32x4.mem\[25\]\[0\] net619 VGND
+ VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3011_ net128 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2726_ net761 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2657_ net767 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1608_ Inst_RegFile_32x4.mem\[6\]\[2\] Inst_RegFile_32x4.mem\[7\]\[2\] net620 VGND
+ VGND VPWR VPWR _0528_ sky130_fd_sc_hd__mux2_1
X_2588_ net773 net716 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1539_ net686 _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__or2_1
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout692 net117 VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__buf_2
Xfanout670 net671 VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__buf_8
Xfanout681 net682 VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__buf_6
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1890_ net402 _0775_ Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q VGND VGND VPWR VPWR
+ _0776_ sky130_fd_sc_hd__mux2_1
XFILLER_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2511_ net754 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2442_ net756 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2373_ net763 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1324_ Inst_RegFile_32x4.mem\[10\]\[2\] Inst_RegFile_32x4.mem\[11\]\[2\] net616 VGND
+ VGND VPWR VPWR _0260_ sky130_fd_sc_hd__mux2_1
X_1255_ net405 net684 net668 net404 Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q
+ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ net691 net671 net657 net653 Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q
+ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_82_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2709_ net56 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput262 net262 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput251 net251 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__buf_8
Xoutput240 net240 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__buf_6
Xoutput284 net284 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput273 net273 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput295 Inst_RegFile_switch_matrix.S1BEG3 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__buf_8
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2991_ SS4END[15] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_2
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1942_ _0698_ _0341_ Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q VGND VGND VPWR VPWR
+ _0821_ sky130_fd_sc_hd__mux2_1
X_1873_ net655 net650 Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _0760_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_54_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2425_ net776 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_63_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2356_ net748 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1307_ Inst_RegFile_32x4.mem\[26\]\[1\] Inst_RegFile_32x4.mem\[27\]\[1\] net619 VGND
+ VGND VPWR VPWR _0245_ sky130_fd_sc_hd__mux2_1
XFILLER_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2287_ clknet_4_10_0_UserCLK_regs _0045_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[23\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1238_ Inst_RegFile_32x4.mem\[6\]\[0\] Inst_RegFile_32x4.mem\[7\]\[0\] net394 VGND
+ VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux2_1
XFILLER_56_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1169_ Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q _1060_ Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q
+ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__o21a_1
XFILLER_52_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2210_ net630 net460 _0961_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__mux2_4
XFILLER_78_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2141_ _0939_ _0923_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__nand2_8
XFILLER_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2072_ _0921_ _0855_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__nor2_8
XFILLER_81_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2974_ S4END[14] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_2
X_1925_ _0801_ _0806_ Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.NN4BEG3 sky130_fd_sc_hd__mux2_1
X_1856_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__inv_1
X_1787_ _0681_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q _0684_ VGND VGND VPWR VPWR
+ _0685_ sky130_fd_sc_hd__o21a_1
XFILLER_69_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2408_ net759 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_4_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2339_ net42 net731 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold61 Inst_RegFile_32x4.mem\[4\]\[2\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold83 Inst_RegFile_32x4.mem\[28\]\[2\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 Inst_RegFile_32x4.mem\[30\]\[2\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold94 Inst_RegFile_32x4.mem\[0\]\[3\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2690_ net41 net729 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_77_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1710_ net64 net1 net80 net7 Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q
+ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__mux4_1
XANTENNA_3 E6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1641_ net782 net94 net122 net139 Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__mux4_1
X_1572_ Inst_RegFile_32x4.mem\[4\]\[3\] Inst_RegFile_32x4.mem\[5\]\[3\] net620 VGND
+ VGND VPWR VPWR _0494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _0941_ net437 VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__nand2_8
XFILLER_81_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2055_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__inv_1
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2957_ net99 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__buf_1
X_2888_ FrameStrobe[16] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_1
X_1908_ Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q _0790_ _0791_ _0788_ VGND VGND
+ VPWR VPWR Inst_RegFile_switch_matrix.EE4BEG1 sky130_fd_sc_hd__o22a_4
X_1839_ Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q _0729_ VGND VGND VPWR VPWR _0730_
+ sky130_fd_sc_hd__nand2_1
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2811_ net20 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_1
X_2742_ clknet_4_15_0_UserCLK_regs _0078_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[19\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2673_ net752 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1624_ net69 net12 net97 net136 Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q
+ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__mux4_2
X_1555_ Inst_RegFile_32x4.mem\[18\]\[3\] Inst_RegFile_32x4.mem\[19\]\[3\] net626 VGND
+ VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1486_ _0410_ _0411_ net688 VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2107_ net506 net606 _0935_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__mux2_4
X_2038_ Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q _0891_ VGND VGND VPWR VPWR _0892_
+ sky130_fd_sc_hd__or2_1
XFILLER_52_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ Inst_RegFile_32x4.mem\[24\]\[2\] Inst_RegFile_32x4.mem\[25\]\[2\] net619 VGND
+ VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1271_ Inst_RegFile_32x4.mem\[26\]\[0\] Inst_RegFile_32x4.mem\[27\]\[0\] net619 VGND
+ VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
XFILLER_83_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3010_ net127 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__buf_1
XFILLER_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2725_ net44 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2656_ net768 net725 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1607_ net686 _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__or2_1
X_2587_ net774 net715 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1538_ Inst_RegFile_32x4.mem\[4\]\[1\] Inst_RegFile_32x4.mem\[5\]\[1\] net432 VGND
+ VGND VPWR VPWR _0462_ sky130_fd_sc_hd__mux2_1
XFILLER_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1469_ Inst_RegFile_32x4.mem\[30\]\[0\] Inst_RegFile_32x4.mem\[31\]\[0\] net624 VGND
+ VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_1
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold180 Inst_RegFile_32x4.mem\[27\]\[3\] VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout660 net661 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__buf_4
Xfanout693 net116 VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__buf_4
Xfanout671 AD0 VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__buf_8
Xfanout682 BD0 VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__buf_8
XFILLER_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2510_ net757 net707 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2441_ net47 net697 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2372_ net764 net736 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1323_ Inst_RegFile_32x4.AD_comb\[1\] Inst_RegFile_32x4.AD_reg\[1\] Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q
+ VGND VGND VPWR VPWR AD1 sky130_fd_sc_hd__mux2_4
X_1254_ Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q _0194_ VGND VGND VPWR VPWR _0195_
+ sky130_fd_sc_hd__or2_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1185_ _1072_ Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q _0129_ VGND VGND VPWR VPWR
+ _0130_ sky130_fd_sc_hd__o21ai_1
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2708_ net55 net745 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput252 net252 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput241 net241 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__buf_8
Xoutput230 net230 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
X_2639_ net754 net724 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput285 net285 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput263 net263 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__buf_6
Xoutput274 net274 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput296 net296 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_8
XFILLER_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2990_ SS4END[14] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1941_ _0816_ _0820_ Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q VGND VGND VPWR VPWR
+ Inst_RegFile_switch_matrix.NN4BEG1 sky130_fd_sc_hd__mux2_4
X_1872_ _1023_ _0751_ _0755_ _0759_ VGND VGND VPWR VPWR Inst_RegFile_switch_matrix.E6BEG1
+ sky130_fd_sc_hd__a31o_4
XFILLER_80_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2424_ net777 net694 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2355_ net750 net735 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1306_ net393 _0239_ _0243_ _0209_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a31o_1
X_2286_ clknet_4_10_0_UserCLK_regs _0044_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[23\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1237_ _0178_ net445 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__nand2b_1
X_1168_ net65 net8 net93 net137 Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q
+ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__mux4_2
X_1099_ Inst_RegFile_32x4.mem\[10\]\[1\] VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_50_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2140_ net574 net603 _0946_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__mux2_4
X_2071_ _0884_ _0919_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__or2_4
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2973_ S4END[13] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_2
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1924_ _0802_ _0803_ _0805_ Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q VGND VGND
+ VPWR VPWR _0806_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1855_ net666 _0697_ Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q VGND VGND VPWR VPWR
+ _0744_ sky130_fd_sc_hd__mux2_1
X_1786_ Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q _0683_ Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2407_ net760 net739 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_4_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2338_ net766 net732 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2269_ clknet_4_12_0_UserCLK_regs _0027_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[30\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold62 Inst_RegFile_32x4.mem\[12\]\[2\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 Inst_RegFile_32x4.mem\[10\]\[2\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold95 Inst_RegFile_32x4.mem\[16\]\[1\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 Inst_RegFile_32x4.mem\[0\]\[0\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1640_ net66 net78 net784 net9 Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q
+ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__mux4_1
XANTENNA_4 E6END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1571_ _0491_ _0492_ net686 VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux2_1
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2123_ _0838_ _0846_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__nor2_8
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2054_ net78 net782 Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q VGND VGND VPWR VPWR
+ _0905_ sky130_fd_sc_hd__mux2_1
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2956_ net98 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_60_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2887_ FrameStrobe[15] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_1
X_1907_ Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q _0789_ Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q
+ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__a21bo_1
X_1838_ net689 _0191_ Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q VGND VGND VPWR VPWR
+ _0729_ sky130_fd_sc_hd__mux2_1
X_1769_ _0666_ _0667_ Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q VGND VGND VPWR VPWR
+ _0668_ sky130_fd_sc_hd__mux2_4
XFILLER_57_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput130 W2MID[4] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_2
XFILLER_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2810_ net19 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_1
XFILLER_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2741_ clknet_4_15_0_UserCLK_regs _0077_ VGND VGND VPWR VPWR Inst_RegFile_32x4.mem\[19\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2672_ net753 net727 VGND VGND VPWR VPWR Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_1623_ net81 net23 net109 Inst_RegFile_switch_matrix.JN2BEG4 Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q
+ Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__mux4_2
X_1554_ Inst_RegFile_32x4.mem\[16\]\[3\] Inst_RegFile_32x4.mem\[17\]\[3\] net626 VGND
+ VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux2_1
X_1485_ Inst_RegFile_32x4.mem\[18\]\[0\] Inst_RegFile_32x4.mem\[19\]\[0\] net627 VGND
+ VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux2_1
.ends

