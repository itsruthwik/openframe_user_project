module LUT4AB (Ci,
    Co,
    UserCLK,
    UserCLKo,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input Ci;
 output Co;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire A;
 wire B;
 wire C;
 wire net141;
 wire D;
 wire E;
 wire net142;
 wire net143;
 wire net412;
 wire net475;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net547;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net525;
 wire net474;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net179;
 wire net512;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire F;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire G;
 wire H;
 wire \Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.M_AB ;
 wire \Inst_LUT4AB_switch_matrix.M_AD ;
 wire \Inst_LUT4AB_switch_matrix.M_AH ;
 wire \Inst_LUT4AB_switch_matrix.M_EF ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG3 ;
 wire net242;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net251;
 wire net252;
 wire net545;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net542;
 wire net543;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net283;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net541;
 wire net546;
 wire net429;
 wire net476;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net548;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net526;
 wire net411;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net544;
 wire net384;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net427;
 wire net428;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;

 sky130_fd_sc_hd__inv_2 _0711_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_1 _0712_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .Y(_0564_));
 sky130_fd_sc_hd__inv_1 _0713_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .Y(_0565_));
 sky130_fd_sc_hd__inv_1 _0714_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .Y(_0566_));
 sky130_fd_sc_hd__inv_1 _0715_ (.A(net75),
    .Y(_0567_));
 sky130_fd_sc_hd__inv_1 _0716_ (.A(net18),
    .Y(_0568_));
 sky130_fd_sc_hd__inv_2 _0717_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .Y(_0569_));
 sky130_fd_sc_hd__inv_1 _0718_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .Y(_0570_));
 sky130_fd_sc_hd__inv_1 _0719_ (.A(net131),
    .Y(_0571_));
 sky130_fd_sc_hd__inv_2 _0720_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .Y(_0572_));
 sky130_fd_sc_hd__inv_1 _0721_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .Y(_0573_));
 sky130_fd_sc_hd__inv_2 _0722_ (.A(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .Y(_0574_));
 sky130_fd_sc_hd__inv_1 _0723_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_0575_));
 sky130_fd_sc_hd__inv_1 _0724_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .Y(_0576_));
 sky130_fd_sc_hd__inv_1 _0725_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0577_));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .Y(_0578_));
 sky130_fd_sc_hd__inv_1 _0727_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .Y(_0579_));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .Y(_0580_));
 sky130_fd_sc_hd__inv_1 _0729_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .Y(_0581_));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .Y(_0582_));
 sky130_fd_sc_hd__inv_1 _0731_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .Y(_0583_));
 sky130_fd_sc_hd__inv_1 _0732_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .Y(_0584_));
 sky130_fd_sc_hd__inv_1 _0733_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ),
    .Y(_0585_));
 sky130_fd_sc_hd__inv_1 _0734_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ),
    .Y(_0586_));
 sky130_fd_sc_hd__mux4_2 _0735_ (.A0(net433),
    .A1(net648),
    .A2(net463),
    .A3(net643),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0587_));
 sky130_fd_sc_hd__mux4_1 _0736_ (.A0(net462),
    .A1(net628),
    .A2(net619),
    .A3(net404),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0588_));
 sky130_fd_sc_hd__or2_1 _0737_ (.A(_0563_),
    .B(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__o21a_1 _0738_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_0587_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0590_));
 sky130_fd_sc_hd__mux4_1 _0739_ (.A0(net805),
    .A1(net95),
    .A2(net123),
    .A3(net135),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0591_));
 sky130_fd_sc_hd__mux4_1 _0740_ (.A0(net61),
    .A1(net67),
    .A2(net79),
    .A3(net10),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _0741_ (.A0(_0591_),
    .A1(_0592_),
    .S(_0563_),
    .X(_0593_));
 sky130_fd_sc_hd__a22o_4 _0742_ (.A1(_0590_),
    .A2(_0589_),
    .B1(_0593_),
    .B2(_0564_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__mux4_2 _0743_ (.A0(net16),
    .A1(net101),
    .A2(net129),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_0594_));
 sky130_fd_sc_hd__mux4_2 _0744_ (.A0(net74),
    .A1(net17),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .X(_0595_));
 sky130_fd_sc_hd__mux4_1 _0745_ (.A0(net433),
    .A1(net639),
    .A2(net624),
    .A3(net645),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_0596_));
 sky130_fd_sc_hd__or2_1 _0746_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .B(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__mux4_1 _0747_ (.A0(net415),
    .A1(net629),
    .A2(net620),
    .A3(net618),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0598_));
 sky130_fd_sc_hd__o21a_1 _0748_ (.A1(_0565_),
    .A2(_0598_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0599_));
 sky130_fd_sc_hd__mux4_1 _0749_ (.A0(net59),
    .A1(net65),
    .A2(net81),
    .A3(net8),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0600_));
 sky130_fd_sc_hd__mux4_1 _0750_ (.A0(net22),
    .A1(net93),
    .A2(net121),
    .A3(net140),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _0751_ (.A0(_0600_),
    .A1(_0601_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0602_));
 sky130_fd_sc_hd__a22o_1 _0752_ (.A1(_0599_),
    .A2(_0597_),
    .B1(_0602_),
    .B2(_0566_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0753_ (.A0(net26),
    .A1(net109),
    .A2(net126),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_0603_));
 sky130_fd_sc_hd__mux4_2 _0754_ (.A0(net83),
    .A1(net93),
    .A2(net8),
    .A3(net121),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_0604_));
 sky130_fd_sc_hd__mux4_2 _0755_ (.A0(_0594_),
    .A1(_0595_),
    .A2(_0604_),
    .A3(_0603_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .X(_0605_));
 sky130_fd_sc_hd__mux4_2 _0756_ (.A0(net634),
    .A1(net411),
    .A2(net412),
    .A3(net416),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0606_));
 sky130_fd_sc_hd__mux4_1 _0757_ (.A0(net653),
    .A1(net649),
    .A2(net624),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0607_));
 sky130_fd_sc_hd__and2b_1 _0758_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .B(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__a21bo_1 _0759_ (.A1(_0606_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0609_));
 sky130_fd_sc_hd__mux4_1 _0760_ (.A0(net67),
    .A1(net807),
    .A2(net79),
    .A3(net10),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0610_));
 sky130_fd_sc_hd__mux4_1 _0761_ (.A0(net805),
    .A1(net95),
    .A2(net123),
    .A3(net135),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _0762_ (.A0(_0610_),
    .A1(_0611_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .X(_0612_));
 sky130_fd_sc_hd__o22a_4 _0763_ (.A1(_0608_),
    .A2(_0609_),
    .B1(_0612_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0764_ (.A0(net77),
    .A1(net105),
    .A2(net133),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_0613_));
 sky130_fd_sc_hd__mux4_2 _0765_ (.A0(net78),
    .A1(net21),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0614_));
 sky130_fd_sc_hd__inv_1 _0766_ (.A(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(_0613_),
    .A1(_0614_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .X(_0616_));
 sky130_fd_sc_hd__mux4_2 _0768_ (.A0(net634),
    .A1(net629),
    .A2(net620),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .X(_0617_));
 sky130_fd_sc_hd__mux4_1 _0769_ (.A0(net434),
    .A1(net638),
    .A2(net624),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_0618_));
 sky130_fd_sc_hd__nand2b_1 _0770_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .B(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__a21boi_2 _0771_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_0617_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .Y(_0620_));
 sky130_fd_sc_hd__mux4_1 _0772_ (.A0(net65),
    .A1(net2),
    .A2(net81),
    .A3(net8),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_0621_));
 sky130_fd_sc_hd__mux4_1 _0773_ (.A0(net805),
    .A1(net93),
    .A2(net121),
    .A3(net135),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _0774_ (.A0(_0621_),
    .A1(_0622_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_0623_));
 sky130_fd_sc_hd__o2bb2a_4 _0775_ (.A1_N(_0619_),
    .A2_N(_0620_),
    .B1(_0623_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _0776_ (.A0(net86),
    .A1(net137),
    .A2(net110),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ),
    .X(_0624_));
 sky130_fd_sc_hd__mux4_2 _0777_ (.A0(net69),
    .A1(net114),
    .A2(net12),
    .A3(net125),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _0778_ (.A0(_0625_),
    .A1(_0624_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(_0616_),
    .A1(_0626_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_4 _0780_ (.A0(_0627_),
    .A1(net1),
    .S(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _0781_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .S(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__mux4_2 _0782_ (.A0(net633),
    .A1(net628),
    .A2(net619),
    .A3(net523),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0630_));
 sky130_fd_sc_hd__mux4_2 _0783_ (.A0(net653),
    .A1(net648),
    .A2(net623),
    .A3(net643),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0631_));
 sky130_fd_sc_hd__or2_4 _0784_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .B(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__o21a_1 _0785_ (.A1(_0630_),
    .A2(_0569_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0633_));
 sky130_fd_sc_hd__mux4_1 _0786_ (.A0(net95),
    .A1(net123),
    .A2(net107),
    .A3(net139),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .X(_0634_));
 sky130_fd_sc_hd__mux4_1 _0787_ (.A0(net67),
    .A1(net807),
    .A2(net10),
    .A3(net805),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _0788_ (.A0(_0634_),
    .A1(_0635_),
    .S(_0569_),
    .X(_0636_));
 sky130_fd_sc_hd__a22o_4 _0789_ (.A1(_0633_),
    .A2(_0632_),
    .B1(_0636_),
    .B2(_0570_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__inv_1 _0790_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .Y(_0637_));
 sky130_fd_sc_hd__mux4_2 _0791_ (.A0(_0567_),
    .A1(_0568_),
    .A2(_0571_),
    .A3(_0637_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_0638_));
 sky130_fd_sc_hd__mux4_2 _0792_ (.A0(net75),
    .A1(net18),
    .A2(net131),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_0639_));
 sky130_fd_sc_hd__mux4_2 _0793_ (.A0(net76),
    .A1(net19),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_0640_));
 sky130_fd_sc_hd__mux4_2 _0794_ (.A0(net653),
    .A1(net444),
    .A2(net623),
    .A3(net643),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_0641_));
 sky130_fd_sc_hd__or2_4 _0795_ (.A(_0641_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0642_));
 sky130_fd_sc_hd__mux4_2 _0796_ (.A0(net462),
    .A1(net411),
    .A2(net619),
    .A3(net416),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_0643_));
 sky130_fd_sc_hd__o21a_1 _0797_ (.A1(_0572_),
    .A2(_0643_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0644_));
 sky130_fd_sc_hd__mux4_1 _0798_ (.A0(net109),
    .A1(net113),
    .A2(net121),
    .A3(net135),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_0645_));
 sky130_fd_sc_hd__mux4_1 _0799_ (.A0(net85),
    .A1(net26),
    .A2(net2),
    .A3(net805),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _0800_ (.A0(_0645_),
    .A1(_0646_),
    .S(_0572_),
    .X(_0647_));
 sky130_fd_sc_hd__a22o_4 _0801_ (.A1(_0644_),
    .A2(_0642_),
    .B1(_0647_),
    .B2(_0573_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG1 ));
 sky130_fd_sc_hd__mux4_2 _0802_ (.A0(net80),
    .A1(net804),
    .A2(net136),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_0648_));
 sky130_fd_sc_hd__mux4_2 _0803_ (.A0(net67),
    .A1(net95),
    .A2(net24),
    .A3(net123),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_0649_));
 sky130_fd_sc_hd__mux4_2 _0804_ (.A0(_0639_),
    .A1(_0640_),
    .A2(_0649_),
    .A3(_0648_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _0805_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S(_0628_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_4 _0806_ (.A0(_0629_),
    .A1(_0651_),
    .S(_0605_),
    .X(_0652_));
 sky130_fd_sc_hd__mux4_1 _0807_ (.A0(net434),
    .A1(net638),
    .A2(net623),
    .A3(net643),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0653_));
 sky130_fd_sc_hd__and2b_1 _0808_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .B(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__mux4_2 _0809_ (.A0(net633),
    .A1(net628),
    .A2(net620),
    .A3(net404),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .X(_0655_));
 sky130_fd_sc_hd__a21bo_1 _0810_ (.A1(_0655_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0656_));
 sky130_fd_sc_hd__mux4_1 _0811_ (.A0(net59),
    .A1(net8),
    .A2(net65),
    .A3(net805),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0657_));
 sky130_fd_sc_hd__mux4_1 _0812_ (.A0(net93),
    .A1(net121),
    .A2(net109),
    .A3(net135),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _0813_ (.A0(_0657_),
    .A1(_0658_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0659_));
 sky130_fd_sc_hd__o22a_4 _0814_ (.A1(_0656_),
    .A2(_0654_),
    .B1(_0659_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG1 ));
 sky130_fd_sc_hd__mux4_1 _0815_ (.A0(net79),
    .A1(net22),
    .A2(net107),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_0660_));
 sky130_fd_sc_hd__mux4_2 _0816_ (.A0(net63),
    .A1(net91),
    .A2(net6),
    .A3(net140),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ),
    .X(_0661_));
 sky130_fd_sc_hd__mux4_2 _0817_ (.A0(net433),
    .A1(net648),
    .A2(net463),
    .A3(net643),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0662_));
 sky130_fd_sc_hd__and2b_1 _0818_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .B(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__mux4_1 _0819_ (.A0(net462),
    .A1(net628),
    .A2(net619),
    .A3(net618),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .X(_0664_));
 sky130_fd_sc_hd__a21bo_1 _0820_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0664_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0665_));
 sky130_fd_sc_hd__mux4_1 _0821_ (.A0(net61),
    .A1(net10),
    .A2(net67),
    .A3(net805),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0666_));
 sky130_fd_sc_hd__mux4_1 _0822_ (.A0(net95),
    .A1(net123),
    .A2(net107),
    .A3(net139),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _0823_ (.A0(_0666_),
    .A1(_0667_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0668_));
 sky130_fd_sc_hd__o22a_4 _0824_ (.A1(_0665_),
    .A2(_0663_),
    .B1(_0668_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG3 ));
 sky130_fd_sc_hd__mux4_1 _0825_ (.A0(net71),
    .A1(net14),
    .A2(net99),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .X(_0669_));
 sky130_fd_sc_hd__mux4_1 _0826_ (.A0(net72),
    .A1(net15),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _0827_ (.A0(_0669_),
    .A1(_0670_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _0828_ (.A0(_0661_),
    .A1(_0660_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _0829_ (.A0(_0671_),
    .A1(_0672_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _0830_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .S(_0628_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _0831_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .S(_0628_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _0832_ (.A0(_0674_),
    .A1(_0675_),
    .S(_0605_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_4 _0833_ (.A0(_0676_),
    .A1(_0652_),
    .S(_0650_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _0834_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .S(_0628_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _0835_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S(_0628_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _0836_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .S(_0628_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _0837_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .S(_0628_),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _0838_ (.A0(_0681_),
    .A1(_0680_),
    .S(_0605_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _0839_ (.A0(_0678_),
    .A1(_0679_),
    .S(_0605_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _0840_ (.A0(_0682_),
    .A1(_0683_),
    .S(_0650_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_4 _0841_ (.A0(_0677_),
    .A1(_0684_),
    .S(_0673_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_4 _0842_ (.A0(_0685_),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(A));
 sky130_fd_sc_hd__mux2_1 _0843_ (.A0(_0669_),
    .A1(_0670_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(_0661_),
    .A1(_0660_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _0845_ (.A0(_0686_),
    .A1(_0687_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _0846_ (.A0(_0613_),
    .A1(_0614_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _0847_ (.A0(_0625_),
    .A1(_0624_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(_0689_),
    .A1(_0690_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ),
    .X(_0691_));
 sky130_fd_sc_hd__o21ai_4 _0849_ (.A1(net1),
    .A2(_0605_),
    .B1(_0650_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_8 _0850_ (.A(_0605_),
    .B(net1),
    .Y(_0693_));
 sky130_fd_sc_hd__nand2_2 _0851_ (.A(_0693_),
    .B(_0692_),
    .Y(_0694_));
 sky130_fd_sc_hd__mux2_4 _0852_ (.A0(_0691_),
    .A1(_0694_),
    .S(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0695_));
 sky130_fd_sc_hd__mux4_2 _0853_ (.A0(_0639_),
    .A1(_0640_),
    .A2(_0649_),
    .A3(_0648_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_0696_));
 sky130_fd_sc_hd__mux4_2 _0854_ (.A0(_0594_),
    .A1(_0595_),
    .A2(_0604_),
    .A3(_0603_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ),
    .X(_0697_));
 sky130_fd_sc_hd__nand2_1 _0855_ (.A(_0696_),
    .B(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__nor2_1 _0856_ (.A(_0696_),
    .B(_0697_),
    .Y(_0699_));
 sky130_fd_sc_hd__mux2_4 _0857_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S(_0695_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_4 _0858_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .S(_0695_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_4 _0859_ (.A0(_0701_),
    .A1(_0700_),
    .S(_0697_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _0860_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .S(_0695_),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _0861_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .S(_0695_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _0862_ (.A0(_0704_),
    .A1(_0703_),
    .S(_0697_),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_4 _0863_ (.A0(_0705_),
    .A1(_0702_),
    .S(_0696_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _0864_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S(_0695_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _0865_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .S(_0695_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _0866_ (.A0(_0708_),
    .A1(_0707_),
    .S(_0697_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _0867_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .S(_0695_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _0868_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .S(_0695_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0869_ (.A0(_0710_),
    .A1(_0008_),
    .S(_0697_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0870_ (.A0(_0009_),
    .A1(_0709_),
    .S(_0696_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_4 _0871_ (.A0(_0706_),
    .A1(_0010_),
    .S(_0688_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_4 _0872_ (.A0(_0011_),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(B));
 sky130_fd_sc_hd__mux4_2 _0873_ (.A0(net656),
    .A1(net649),
    .A2(net639),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0012_));
 sky130_fd_sc_hd__mux4_1 _0874_ (.A0(net636),
    .A1(net630),
    .A2(net622),
    .A3(net402),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_4 _0875_ (.A0(_0012_),
    .A1(_0013_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0014_));
 sky130_fd_sc_hd__mux4_1 _0876_ (.A0(net60),
    .A1(net82),
    .A2(net66),
    .A3(net9),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .X(_0015_));
 sky130_fd_sc_hd__mux4_1 _0877_ (.A0(net804),
    .A1(net94),
    .A2(net122),
    .A3(net136),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0878_ (.A0(_0015_),
    .A1(_0016_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_4 _0879_ (.A0(_0017_),
    .A1(_0014_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _0880_ (.A0(net81),
    .A1(net8),
    .A2(net126),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ),
    .X(_0018_));
 sky130_fd_sc_hd__mux4_2 _0881_ (.A0(net65),
    .A1(net8),
    .A2(net93),
    .A3(net139),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ),
    .X(_0019_));
 sky130_fd_sc_hd__mux4_1 _0882_ (.A0(net654),
    .A1(net650),
    .A2(net625),
    .A3(net641),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0020_));
 sky130_fd_sc_hd__and2b_1 _0883_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .B(_0020_),
    .X(_0021_));
 sky130_fd_sc_hd__mux4_2 _0884_ (.A0(net635),
    .A1(net630),
    .A2(net621),
    .A3(net617),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0022_));
 sky130_fd_sc_hd__a21bo_1 _0885_ (.A1(_0022_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_0023_));
 sky130_fd_sc_hd__mux4_1 _0886_ (.A0(net88),
    .A1(net96),
    .A2(net90),
    .A3(net116),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0024_));
 sky130_fd_sc_hd__mux4_1 _0887_ (.A0(net60),
    .A1(net68),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _0888_ (.A0(_0025_),
    .A1(_0024_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .X(_0026_));
 sky130_fd_sc_hd__o22ai_4 _0889_ (.A1(_0023_),
    .A2(_0021_),
    .B1(_0026_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_6 _0890_ (.A(net474),
    .Y(\Inst_LUT4AB_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _0891_ (.A0(net73),
    .A1(net129),
    .A2(net16),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0028_));
 sky130_fd_sc_hd__mux4_2 _0892_ (.A0(net74),
    .A1(net17),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0029_));
 sky130_fd_sc_hd__mux4_2 _0893_ (.A0(_0028_),
    .A1(_0029_),
    .A2(_0019_),
    .A3(_0018_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ),
    .X(_0030_));
 sky130_fd_sc_hd__mux4_2 _0894_ (.A0(net653),
    .A1(net649),
    .A2(net639),
    .A3(net645),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0031_));
 sky130_fd_sc_hd__and2b_1 _0895_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .B(_0031_),
    .X(_0032_));
 sky130_fd_sc_hd__mux4_2 _0896_ (.A0(net634),
    .A1(net629),
    .A2(net620),
    .A3(net483),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0033_));
 sky130_fd_sc_hd__a21bo_1 _0897_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(_0033_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0034_));
 sky130_fd_sc_hd__mux4_1 _0898_ (.A0(net94),
    .A1(net122),
    .A2(net110),
    .A3(net136),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0035_));
 sky130_fd_sc_hd__mux4_1 _0899_ (.A0(net86),
    .A1(net3),
    .A2(net9),
    .A3(net23),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0900_ (.A0(_0036_),
    .A1(_0035_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0037_));
 sky130_fd_sc_hd__o22a_4 _0901_ (.A1(_0034_),
    .A2(_0032_),
    .B1(_0037_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _0902_ (.A0(net84),
    .A1(net25),
    .A2(net108),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ),
    .X(_0038_));
 sky130_fd_sc_hd__mux4_2 _0903_ (.A0(net67),
    .A1(net10),
    .A2(net113),
    .A3(net123),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ),
    .X(_0039_));
 sky130_fd_sc_hd__mux4_1 _0904_ (.A0(net654),
    .A1(net650),
    .A2(net625),
    .A3(net641),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0040_));
 sky130_fd_sc_hd__mux4_2 _0905_ (.A0(net635),
    .A1(net630),
    .A2(net621),
    .A3(net403),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_4 _0906_ (.A0(_0040_),
    .A1(_0041_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0042_));
 sky130_fd_sc_hd__mux4_1 _0907_ (.A0(net60),
    .A1(net68),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0043_));
 sky130_fd_sc_hd__mux4_1 _0908_ (.A0(net88),
    .A1(net96),
    .A2(net116),
    .A3(net659),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0909_ (.A0(_0043_),
    .A1(_0044_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_4 _0910_ (.A0(_0045_),
    .A1(_0042_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__mux4_2 _0911_ (.A0(net75),
    .A1(net18),
    .A2(net103),
    .A3(net488),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_0046_));
 sky130_fd_sc_hd__mux4_1 _0912_ (.A0(net76),
    .A1(net19),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ),
    .X(_0047_));
 sky130_fd_sc_hd__mux4_2 _0913_ (.A0(net525),
    .A1(_0047_),
    .A2(_0039_),
    .A3(_0038_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_0048_));
 sky130_fd_sc_hd__inv_2 _0914_ (.A(_0048_),
    .Y(_0049_));
 sky130_fd_sc_hd__or2_4 _0915_ (.A(_0030_),
    .B(_0048_),
    .X(_0050_));
 sky130_fd_sc_hd__nand2_1 _0916_ (.A(_0030_),
    .B(_0048_),
    .Y(_0051_));
 sky130_fd_sc_hd__mux4_2 _0917_ (.A0(_0028_),
    .A1(_0029_),
    .A2(_0019_),
    .A3(_0018_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_2 _0918_ (.A0(net525),
    .A1(_0047_),
    .A2(_0039_),
    .A3(_0038_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .X(_0053_));
 sky130_fd_sc_hd__inv_2 _0919_ (.A(_0053_),
    .Y(_0054_));
 sky130_fd_sc_hd__or2_2 _0920_ (.A(_0052_),
    .B(_0053_),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(_0052_),
    .B(_0053_),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_1 _0922_ (.A(_0052_),
    .B(_0053_),
    .Y(_0057_));
 sky130_fd_sc_hd__a31oi_4 _0923_ (.A1(_0692_),
    .A2(_0693_),
    .A3(_0698_),
    .B1(_0699_),
    .Y(_0058_));
 sky130_fd_sc_hd__a21o_1 _0924_ (.A1(_0058_),
    .A2(_0055_),
    .B1(_0056_),
    .X(_0059_));
 sky130_fd_sc_hd__a221o_1 _0925_ (.A1(_0048_),
    .A2(_0030_),
    .B1(_0055_),
    .B2(_0058_),
    .C1(_0056_),
    .X(_0060_));
 sky130_fd_sc_hd__mux4_1 _0926_ (.A0(net655),
    .A1(net650),
    .A2(net625),
    .A3(net640),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0061_));
 sky130_fd_sc_hd__mux4_2 _0927_ (.A0(net646),
    .A1(net631),
    .A2(net621),
    .A3(net524),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_4 _0928_ (.A0(_0061_),
    .A1(_0062_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0063_));
 sky130_fd_sc_hd__mux4_1 _0929_ (.A0(net61),
    .A1(net69),
    .A2(net807),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .X(_0064_));
 sky130_fd_sc_hd__mux4_1 _0930_ (.A0(net89),
    .A1(net115),
    .A2(net97),
    .A3(net660),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0931_ (.A0(_0064_),
    .A1(_0065_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_4 _0932_ (.A0(_0066_),
    .A1(_0063_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0933_ (.A0(net77),
    .A1(net133),
    .A2(net20),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0067_));
 sky130_fd_sc_hd__mux4_2 _0934_ (.A0(net78),
    .A1(net21),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0068_));
 sky130_fd_sc_hd__mux4_2 _0935_ (.A0(net82),
    .A1(net122),
    .A2(net9),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_0069_));
 sky130_fd_sc_hd__mux4_1 _0936_ (.A0(net70),
    .A1(net98),
    .A2(net26),
    .A3(net126),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0070_));
 sky130_fd_sc_hd__a21bo_1 _0937_ (.A1(_0060_),
    .A2(_0050_),
    .B1_N(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0071_));
 sky130_fd_sc_hd__mux4_2 _0938_ (.A0(_0067_),
    .A1(_0068_),
    .A2(_0070_),
    .A3(_0069_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_0072_));
 sky130_fd_sc_hd__o21ai_4 _0939_ (.A1(_0072_),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .B1(_0071_),
    .Y(_0073_));
 sky130_fd_sc_hd__mux4_1 _0940_ (.A0(net654),
    .A1(net650),
    .A2(net626),
    .A3(net640),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0074_));
 sky130_fd_sc_hd__nand2b_1 _0941_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .B(_0074_),
    .Y(_0075_));
 sky130_fd_sc_hd__mux4_2 _0942_ (.A0(net646),
    .A1(net631),
    .A2(net621),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0076_));
 sky130_fd_sc_hd__a21boi_2 _0943_ (.A1(_0076_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0077_));
 sky130_fd_sc_hd__mux4_1 _0944_ (.A0(net61),
    .A1(net69),
    .A2(net807),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .X(_0078_));
 sky130_fd_sc_hd__mux4_1 _0945_ (.A0(net89),
    .A1(net115),
    .A2(net97),
    .A3(net660),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(_0078_),
    .A1(_0079_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_0080_));
 sky130_fd_sc_hd__a2bb2o_4 _0947_ (.A1_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .A2_N(_0080_),
    .B1(_0075_),
    .B2(_0077_),
    .X(_0081_));
 sky130_fd_sc_hd__inv_2 _0948_ (.A(_0081_),
    .Y(\Inst_LUT4AB_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _0949_ (.A0(net75),
    .A1(net131),
    .A2(net103),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_0082_));
 sky130_fd_sc_hd__mux4_1 _0950_ (.A0(net76),
    .A1(net19),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ),
    .X(_0083_));
 sky130_fd_sc_hd__mux4_2 _0951_ (.A0(net80),
    .A1(net112),
    .A2(net123),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ),
    .X(_0084_));
 sky130_fd_sc_hd__mux4_2 _0952_ (.A0(net68),
    .A1(net11),
    .A2(net112),
    .A3(net124),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .X(_0085_));
 sky130_fd_sc_hd__mux4_2 _0953_ (.A0(_0082_),
    .A1(_0083_),
    .A2(_0085_),
    .A3(_0084_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0086_));
 sky130_fd_sc_hd__mux4_2 _0954_ (.A0(net85),
    .A1(net109),
    .A2(net8),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0087_));
 sky130_fd_sc_hd__mux4_2 _0955_ (.A0(net66),
    .A1(net94),
    .A2(net9),
    .A3(net138),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .X(_0088_));
 sky130_fd_sc_hd__mux4_1 _0956_ (.A0(net657),
    .A1(net652),
    .A2(net627),
    .A3(net642),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0089_));
 sky130_fd_sc_hd__and2b_1 _0957_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .B(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__mux4_1 _0958_ (.A0(net647),
    .A1(net632),
    .A2(net622),
    .A3(net618),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0091_));
 sky130_fd_sc_hd__a21bo_1 _0959_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0091_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0092_));
 sky130_fd_sc_hd__mux4_1 _0960_ (.A0(net61),
    .A1(net69),
    .A2(net807),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0093_));
 sky130_fd_sc_hd__mux4_1 _0961_ (.A0(net87),
    .A1(net89),
    .A2(net97),
    .A3(net660),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0962_ (.A0(_0093_),
    .A1(_0094_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0095_));
 sky130_fd_sc_hd__o22a_4 _0963_ (.A1(_0090_),
    .A2(_0092_),
    .B1(_0095_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__mux4_1 _0964_ (.A0(net73),
    .A1(net101),
    .A2(net16),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0096_));
 sky130_fd_sc_hd__mux4_2 _0965_ (.A0(net74),
    .A1(net17),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_0097_));
 sky130_fd_sc_hd__mux4_2 _0966_ (.A0(_0096_),
    .A1(_0097_),
    .A2(_0088_),
    .A3(_0087_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .X(_0098_));
 sky130_fd_sc_hd__inv_2 _0967_ (.A(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__or2_1 _0968_ (.A(_0086_),
    .B(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_4 _0969_ (.A(_0098_),
    .B(_0086_),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__o22a_1 _0971_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0100_),
    .B1(_0101_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .X(_0103_));
 sky130_fd_sc_hd__nand2_1 _0972_ (.A(_0086_),
    .B(_0099_),
    .Y(_0104_));
 sky130_fd_sc_hd__or2_2 _0973_ (.A(_0086_),
    .B(_0098_),
    .X(_0105_));
 sky130_fd_sc_hd__o22a_1 _0974_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0104_),
    .B1(_0105_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .X(_0106_));
 sky130_fd_sc_hd__a21bo_1 _0975_ (.A1(_0103_),
    .A2(_0106_),
    .B1_N(_0073_),
    .X(_0107_));
 sky130_fd_sc_hd__o22a_1 _0976_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0101_),
    .B1(_0104_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .X(_0108_));
 sky130_fd_sc_hd__o22a_1 _0977_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0100_),
    .B1(_0105_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .X(_0109_));
 sky130_fd_sc_hd__a21o_1 _0978_ (.A1(_0108_),
    .A2(_0109_),
    .B1(_0073_),
    .X(_0110_));
 sky130_fd_sc_hd__mux4_1 _0979_ (.A0(net654),
    .A1(net650),
    .A2(net625),
    .A3(net640),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0111_));
 sky130_fd_sc_hd__and2b_1 _0980_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .B(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__mux4_1 _0981_ (.A0(net646),
    .A1(net630),
    .A2(net621),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0113_));
 sky130_fd_sc_hd__a21bo_1 _0982_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(_0113_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0114_));
 sky130_fd_sc_hd__mux4_1 _0983_ (.A0(net61),
    .A1(net69),
    .A2(net807),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0115_));
 sky130_fd_sc_hd__mux4_1 _0984_ (.A0(net87),
    .A1(net89),
    .A2(net97),
    .A3(net660),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0985_ (.A0(_0115_),
    .A1(_0116_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0117_));
 sky130_fd_sc_hd__o22a_2 _0986_ (.A1(_0112_),
    .A2(_0114_),
    .B1(_0117_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG5 ));
 sky130_fd_sc_hd__mux4_2 _0987_ (.A0(net14),
    .A1(net99),
    .A2(net127),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ),
    .X(_0118_));
 sky130_fd_sc_hd__mux4_1 _0988_ (.A0(net72),
    .A1(net15),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_0119_));
 sky130_fd_sc_hd__mux4_2 _0989_ (.A0(net27),
    .A1(net138),
    .A2(net107),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_0120_));
 sky130_fd_sc_hd__mux4_2 _0990_ (.A0(net85),
    .A1(net7),
    .A2(net92),
    .A3(net120),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(_0118_),
    .A1(_0119_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_4 _0992_ (.A0(_0121_),
    .A1(_0120_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_4 _0993_ (.A0(_0122_),
    .A1(_0123_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_0124_));
 sky130_fd_sc_hd__o22a_1 _0994_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0100_),
    .B1(_0101_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .X(_0125_));
 sky130_fd_sc_hd__o22a_1 _0995_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0104_),
    .B1(_0105_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .X(_0126_));
 sky130_fd_sc_hd__a21bo_1 _0996_ (.A1(_0125_),
    .A2(_0126_),
    .B1_N(_0073_),
    .X(_0127_));
 sky130_fd_sc_hd__o22a_1 _0997_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0100_),
    .B1(_0101_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .X(_0128_));
 sky130_fd_sc_hd__o221a_1 _0998_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0104_),
    .B1(_0105_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .C1(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__o21ba_1 _0999_ (.A1(_0073_),
    .A2(_0129_),
    .B1_N(_0124_),
    .X(_0130_));
 sky130_fd_sc_hd__a32o_1 _1000_ (.A1(_0124_),
    .A2(_0110_),
    .A3(_0107_),
    .B1(_0127_),
    .B2(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_4 _1001_ (.A0(_0131_),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(E));
 sky130_fd_sc_hd__mux4_1 _1002_ (.A0(net654),
    .A1(net650),
    .A2(net625),
    .A3(net641),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0132_));
 sky130_fd_sc_hd__mux4_1 _1003_ (.A0(net478),
    .A1(net630),
    .A2(net621),
    .A3(net618),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(_0132_),
    .A1(_0133_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .X(_0134_));
 sky130_fd_sc_hd__mux4_1 _1005_ (.A0(net88),
    .A1(net96),
    .A2(net116),
    .A3(net659),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0135_));
 sky130_fd_sc_hd__mux4_1 _1006_ (.A0(net60),
    .A1(net68),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _1007_ (.A0(_0136_),
    .A1(_0135_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_4 _1008_ (.A0(_0137_),
    .A1(_0134_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _1009_ (.A0(net20),
    .A1(net133),
    .A2(net105),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0138_));
 sky130_fd_sc_hd__mux4_1 _1010_ (.A0(net78),
    .A1(net21),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _1011_ (.A0(_0138_),
    .A1(_0139_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_0140_));
 sky130_fd_sc_hd__mux4_1 _1012_ (.A0(net656),
    .A1(net651),
    .A2(net642),
    .A3(net647),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0141_));
 sky130_fd_sc_hd__and2b_1 _1013_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .B(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__mux4_2 _1014_ (.A0(net637),
    .A1(net630),
    .A2(net622),
    .A3(net407),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0143_));
 sky130_fd_sc_hd__a21bo_1 _1015_ (.A1(_0143_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0144_));
 sky130_fd_sc_hd__mux4_1 _1016_ (.A0(net66),
    .A1(net82),
    .A2(net3),
    .A3(net9),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0145_));
 sky130_fd_sc_hd__mux4_1 _1017_ (.A0(net804),
    .A1(net94),
    .A2(net122),
    .A3(net138),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _1018_ (.A0(_0145_),
    .A1(_0146_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0147_));
 sky130_fd_sc_hd__o22a_4 _1019_ (.A1(_0144_),
    .A2(_0142_),
    .B1(_0147_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1020_ (.A0(net9),
    .A1(net139),
    .A2(net114),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_0148_));
 sky130_fd_sc_hd__mux4_1 _1021_ (.A0(net86),
    .A1(net97),
    .A2(net12),
    .A3(net125),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _1022_ (.A0(_0149_),
    .A1(_0148_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _1023_ (.A0(_0140_),
    .A1(_0150_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _1024_ (.A0(_0151_),
    .A1(_0058_),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0152_));
 sky130_fd_sc_hd__nand2_1 _1025_ (.A(_0052_),
    .B(_0054_),
    .Y(_0153_));
 sky130_fd_sc_hd__o22a_1 _1026_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0057_),
    .B1(_0153_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .X(_0154_));
 sky130_fd_sc_hd__or2_1 _1027_ (.A(_0052_),
    .B(_0054_),
    .X(_0155_));
 sky130_fd_sc_hd__or2_1 _1028_ (.A(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .B(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__o211a_1 _1029_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0055_),
    .B1(_0154_),
    .C1(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__mux4_1 _1030_ (.A0(net654),
    .A1(net650),
    .A2(net625),
    .A3(net641),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0158_));
 sky130_fd_sc_hd__mux4_2 _1031_ (.A0(net478),
    .A1(net630),
    .A2(net621),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_4 _1032_ (.A0(_0158_),
    .A1(_0159_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0160_));
 sky130_fd_sc_hd__mux4_1 _1033_ (.A0(net60),
    .A1(net68),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0161_));
 sky130_fd_sc_hd__mux4_1 _1034_ (.A0(net88),
    .A1(net96),
    .A2(net90),
    .A3(net116),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _1035_ (.A0(_0161_),
    .A1(_0162_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_4 _1036_ (.A0(_0163_),
    .A1(_0160_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG4 ));
 sky130_fd_sc_hd__mux4_1 _1037_ (.A0(net71),
    .A1(net99),
    .A2(net127),
    .A3(net479),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_0164_));
 sky130_fd_sc_hd__mux4_2 _1038_ (.A0(net72),
    .A1(net15),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ),
    .X(_0165_));
 sky130_fd_sc_hd__mux4_2 _1039_ (.A0(net653),
    .A1(net648),
    .A2(net444),
    .A3(net644),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0166_));
 sky130_fd_sc_hd__mux4_1 _1040_ (.A0(net462),
    .A1(net628),
    .A2(net412),
    .A3(net416),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_4 _1041_ (.A0(_0166_),
    .A1(_0167_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0168_));
 sky130_fd_sc_hd__mux4_1 _1042_ (.A0(net110),
    .A1(net122),
    .A2(net114),
    .A3(net136),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .X(_0169_));
 sky130_fd_sc_hd__mux4_1 _1043_ (.A0(net60),
    .A1(net66),
    .A2(net27),
    .A3(net804),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _1044_ (.A0(_0170_),
    .A1(_0169_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_4 _1045_ (.A0(_0171_),
    .A1(_0168_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1046_ (.A0(net79),
    .A1(net135),
    .A2(net111),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_0172_));
 sky130_fd_sc_hd__mux4_2 _1047_ (.A0(net63),
    .A1(net91),
    .A2(net25),
    .A3(net119),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .X(_0173_));
 sky130_fd_sc_hd__mux4_2 _1048_ (.A0(_0164_),
    .A1(_0165_),
    .A2(_0173_),
    .A3(_0172_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .X(_0174_));
 sky130_fd_sc_hd__o22a_1 _1049_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(_0057_),
    .B1(_0153_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _1050_ (.A(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .B(_0155_),
    .X(_0176_));
 sky130_fd_sc_hd__o211a_1 _1051_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0055_),
    .B1(_0175_),
    .C1(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _1052_ (.A0(_0177_),
    .A1(_0157_),
    .S(_0152_),
    .X(_0178_));
 sky130_fd_sc_hd__o22a_1 _1053_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0055_),
    .B1(_0153_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .X(_0179_));
 sky130_fd_sc_hd__o22a_1 _1054_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0057_),
    .B1(_0155_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .X(_0180_));
 sky130_fd_sc_hd__a21oi_1 _1055_ (.A1(_0179_),
    .A2(_0180_),
    .B1(_0152_),
    .Y(_0181_));
 sky130_fd_sc_hd__o22a_1 _1056_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0057_),
    .B1(_0155_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .X(_0182_));
 sky130_fd_sc_hd__o22a_1 _1057_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0055_),
    .B1(_0153_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_1 _1058_ (.A(_0182_),
    .B(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__a21oi_1 _1059_ (.A1(_0152_),
    .A2(_0184_),
    .B1(_0181_),
    .Y(_0185_));
 sky130_fd_sc_hd__mux2_4 _1060_ (.A0(_0178_),
    .A1(_0185_),
    .S(_0174_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_4 _1061_ (.A0(_0186_),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(C));
 sky130_fd_sc_hd__mux4_2 _1062_ (.A0(_0067_),
    .A1(_0068_),
    .A2(_0070_),
    .A3(_0069_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_0187_));
 sky130_fd_sc_hd__a31o_1 _1063_ (.A1(_0105_),
    .A2(_0060_),
    .A3(_0050_),
    .B1(_0102_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_4 _1064_ (.A0(_0187_),
    .A1(_0188_),
    .S(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0189_));
 sky130_fd_sc_hd__mux4_2 _1065_ (.A0(_0082_),
    .A1(_0083_),
    .A2(_0085_),
    .A3(_0084_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .X(_0190_));
 sky130_fd_sc_hd__mux4_2 _1066_ (.A0(_0096_),
    .A1(_0097_),
    .A2(_0088_),
    .A3(_0087_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .X(_0191_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__nand2_1 _1068_ (.A(_0190_),
    .B(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__or2_1 _1069_ (.A(_0190_),
    .B(_0192_),
    .X(_0194_));
 sky130_fd_sc_hd__or2_1 _1070_ (.A(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__nand2_1 _1071_ (.A(_0190_),
    .B(_0191_),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_1 _1072_ (.A(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__or2_4 _1073_ (.A(_0190_),
    .B(_0191_),
    .X(_0198_));
 sky130_fd_sc_hd__o22a_1 _1074_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0193_),
    .B1(_0196_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .X(_0199_));
 sky130_fd_sc_hd__o211a_1 _1075_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0198_),
    .B1(_0199_),
    .C1(_0195_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _1076_ (.A0(_0118_),
    .A1(_0119_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_4 _1077_ (.A0(_0121_),
    .A1(_0120_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_4 _1078_ (.A0(_0201_),
    .A1(_0202_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0203_));
 sky130_fd_sc_hd__o22a_1 _1079_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A2(_0193_),
    .B1(_0194_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .X(_0204_));
 sky130_fd_sc_hd__o221a_1 _1080_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0196_),
    .B1(_0198_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .C1(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_4 _1081_ (.A0(_0200_),
    .A1(_0205_),
    .S(_0189_),
    .X(_0206_));
 sky130_fd_sc_hd__o22a_1 _1082_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0193_),
    .B1(_0194_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .X(_0207_));
 sky130_fd_sc_hd__o221a_1 _1083_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0196_),
    .B1(_0198_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .C1(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__or2_1 _1084_ (.A(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .B(_0194_),
    .X(_0209_));
 sky130_fd_sc_hd__o22a_1 _1085_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0193_),
    .B1(_0198_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .X(_0210_));
 sky130_fd_sc_hd__o211a_1 _1086_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(_0196_),
    .B1(_0209_),
    .C1(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _1087_ (.A0(_0211_),
    .A1(_0208_),
    .S(_0189_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_4 _1088_ (.A0(_0212_),
    .A1(_0206_),
    .S(_0203_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_4 _1089_ (.A0(_0213_),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(F));
 sky130_fd_sc_hd__a311o_1 _1090_ (.A1(_0050_),
    .A2(_0060_),
    .A3(_0105_),
    .B1(_0102_),
    .C1(_0197_),
    .X(_0214_));
 sky130_fd_sc_hd__mux4_1 _1091_ (.A0(net655),
    .A1(net650),
    .A2(net626),
    .A3(net641),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0215_));
 sky130_fd_sc_hd__mux4_2 _1092_ (.A0(net646),
    .A1(net621),
    .A2(net477),
    .A3(net405),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_4 _1093_ (.A0(_0215_),
    .A1(_0216_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0217_));
 sky130_fd_sc_hd__mux4_1 _1094_ (.A0(net90),
    .A1(net116),
    .A2(net98),
    .A3(net659),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .X(_0218_));
 sky130_fd_sc_hd__mux4_1 _1095_ (.A0(net62),
    .A1(net70),
    .A2(net5),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(_0219_),
    .A1(_0218_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_4 _1097_ (.A0(_0220_),
    .A1(_0217_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1098_ (.A0(net77),
    .A1(net105),
    .A2(net20),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_0221_));
 sky130_fd_sc_hd__mux4_1 _1099_ (.A0(net78),
    .A1(net21),
    .A2(net106),
    .A3(net134),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_0222_));
 sky130_fd_sc_hd__mux4_1 _1100_ (.A0(net82),
    .A1(net24),
    .A2(net110),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0223_));
 sky130_fd_sc_hd__mux4_2 _1101_ (.A0(net70),
    .A1(net13),
    .A2(net98),
    .A3(net137),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_0224_));
 sky130_fd_sc_hd__mux4_2 _1102_ (.A0(_0221_),
    .A1(_0222_),
    .A2(_0224_),
    .A3(_0223_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_0225_));
 sky130_fd_sc_hd__and2b_1 _1103_ (.A_N(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ),
    .B(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__a31o_1 _1104_ (.A1(_0214_),
    .A2(_0198_),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ),
    .B1(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__mux4_1 _1105_ (.A0(net657),
    .A1(net651),
    .A2(net626),
    .A3(net640),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0228_));
 sky130_fd_sc_hd__and2b_1 _1106_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .B(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__mux4_2 _1107_ (.A0(net646),
    .A1(net427),
    .A2(net635),
    .A3(net430),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0230_));
 sky130_fd_sc_hd__a21bo_1 _1108_ (.A1(_0230_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_0231_));
 sky130_fd_sc_hd__mux4_1 _1109_ (.A0(net62),
    .A1(net70),
    .A2(net806),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .X(_0232_));
 sky130_fd_sc_hd__mux4_1 _1110_ (.A0(net90),
    .A1(net116),
    .A2(net98),
    .A3(net659),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _1111_ (.A0(_0232_),
    .A1(_0233_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_0234_));
 sky130_fd_sc_hd__o22a_1 _1112_ (.A1(_0231_),
    .A2(_0229_),
    .B1(_0234_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__mux4_2 _1113_ (.A0(net18),
    .A1(net131),
    .A2(net103),
    .A3(net429),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0235_));
 sky130_fd_sc_hd__mux4_1 _1114_ (.A0(net76),
    .A1(net19),
    .A2(net104),
    .A3(net132),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .X(_0236_));
 sky130_fd_sc_hd__mux4_2 _1115_ (.A0(net23),
    .A1(net108),
    .A2(net140),
    .A3(net489),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_0237_));
 sky130_fd_sc_hd__mux4_2 _1116_ (.A0(net84),
    .A1(net96),
    .A2(net11),
    .A3(net124),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ),
    .X(_0238_));
 sky130_fd_sc_hd__mux4_2 _1117_ (.A0(_0235_),
    .A1(_0236_),
    .A2(_0238_),
    .A3(_0237_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ),
    .X(_0239_));
 sky130_fd_sc_hd__mux4_1 _1118_ (.A0(net656),
    .A1(net652),
    .A2(net627),
    .A3(net640),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0240_));
 sky130_fd_sc_hd__mux4_2 _1119_ (.A0(net647),
    .A1(net485),
    .A2(net637),
    .A3(net402),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_4 _1120_ (.A0(_0240_),
    .A1(_0241_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_0242_));
 sky130_fd_sc_hd__mux4_1 _1121_ (.A0(net88),
    .A1(net90),
    .A2(net98),
    .A3(net659),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0243_));
 sky130_fd_sc_hd__mux4_1 _1122_ (.A0(net62),
    .A1(net70),
    .A2(net806),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _1123_ (.A0(_0244_),
    .A1(_0243_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_4 _1124_ (.A0(_0245_),
    .A1(_0242_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _1125_ (.A0(net73),
    .A1(net129),
    .A2(net101),
    .A3(net413),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_0246_));
 sky130_fd_sc_hd__mux4_2 _1126_ (.A0(net74),
    .A1(net17),
    .A2(net102),
    .A3(net130),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ),
    .X(_0247_));
 sky130_fd_sc_hd__mux4_2 _1127_ (.A0(net81),
    .A1(net121),
    .A2(net113),
    .A3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_0248_));
 sky130_fd_sc_hd__mux4_2 _1128_ (.A0(net66),
    .A1(net111),
    .A2(net9),
    .A3(net122),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ),
    .X(_0249_));
 sky130_fd_sc_hd__mux4_2 _1129_ (.A0(_0246_),
    .A1(_0247_),
    .A2(_0249_),
    .A3(_0248_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .X(_0250_));
 sky130_fd_sc_hd__or2_1 _1130_ (.A(_0239_),
    .B(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__and2_1 _1131_ (.A(_0239_),
    .B(_0250_),
    .X(_0252_));
 sky130_fd_sc_hd__inv_1 _1132_ (.A(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__mux4_1 _1133_ (.A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S0(_0250_),
    .S1(_0239_),
    .X(_0254_));
 sky130_fd_sc_hd__mux4_2 _1134_ (.A0(net83),
    .A1(net119),
    .A2(net805),
    .A3(net479),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0255_));
 sky130_fd_sc_hd__mux4_2 _1135_ (.A0(net64),
    .A1(net92),
    .A2(net27),
    .A3(net120),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .X(_0256_));
 sky130_fd_sc_hd__mux4_1 _1136_ (.A0(net655),
    .A1(net651),
    .A2(net625),
    .A3(net640),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0257_));
 sky130_fd_sc_hd__and2b_1 _1137_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .B(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__mux4_2 _1138_ (.A0(net646),
    .A1(net621),
    .A2(net635),
    .A3(net417),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0259_));
 sky130_fd_sc_hd__a21bo_1 _1139_ (.A1(_0259_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0260_));
 sky130_fd_sc_hd__mux4_1 _1140_ (.A0(net62),
    .A1(net70),
    .A2(net806),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0261_));
 sky130_fd_sc_hd__mux4_1 _1141_ (.A0(net88),
    .A1(net90),
    .A2(net98),
    .A3(net659),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _1142_ (.A0(_0261_),
    .A1(_0262_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_0263_));
 sky130_fd_sc_hd__o22a_4 _1143_ (.A1(_0260_),
    .A2(_0258_),
    .B1(_0263_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__mux4_1 _1144_ (.A0(net71),
    .A1(net14),
    .A2(net127),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .X(_0264_));
 sky130_fd_sc_hd__mux4_1 _1145_ (.A0(net72),
    .A1(net15),
    .A2(net100),
    .A3(net128),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .X(_0265_));
 sky130_fd_sc_hd__mux4_2 _1146_ (.A0(_0264_),
    .A1(_0265_),
    .A2(_0256_),
    .A3(_0255_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .X(_0266_));
 sky130_fd_sc_hd__mux4_1 _1147_ (.A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .S0(_0250_),
    .S1(_0239_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_4 _1148_ (.A0(_0267_),
    .A1(_0254_),
    .S(_0227_),
    .X(_0268_));
 sky130_fd_sc_hd__mux4_1 _1149_ (.A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S0(_0250_),
    .S1(_0239_),
    .X(_0269_));
 sky130_fd_sc_hd__or3b_1 _1150_ (.A(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .B(_0239_),
    .C_N(_0250_),
    .X(_0270_));
 sky130_fd_sc_hd__or3b_1 _1151_ (.A(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .B(_0250_),
    .C_N(_0239_),
    .X(_0271_));
 sky130_fd_sc_hd__o22a_1 _1152_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0251_),
    .B1(_0253_),
    .B2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .X(_0272_));
 sky130_fd_sc_hd__and3_1 _1153_ (.A(_0270_),
    .B(_0271_),
    .C(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _1154_ (.A0(_0269_),
    .A1(_0273_),
    .S(_0227_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_4 _1155_ (.A0(_0274_),
    .A1(_0268_),
    .S(_0266_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_4 _1156_ (.A0(_0275_),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(G));
 sky130_fd_sc_hd__a31o_4 _1157_ (.A1(_0251_),
    .A2(_0214_),
    .A3(_0198_),
    .B1(_0252_),
    .X(_0276_));
 sky130_fd_sc_hd__mux4_1 _1158_ (.A0(_0221_),
    .A1(_0222_),
    .A2(_0224_),
    .A3(_0223_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .X(_0277_));
 sky130_fd_sc_hd__nand2b_1 _1159_ (.A_N(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .B(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _1160_ (.A(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__a21oi_4 _1161_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0276_),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__mux4_2 _1162_ (.A0(_0235_),
    .A1(_0236_),
    .A2(_0238_),
    .A3(_0237_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_0281_));
 sky130_fd_sc_hd__mux4_2 _1163_ (.A0(_0246_),
    .A1(_0247_),
    .A2(_0249_),
    .A3(_0248_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .X(_0282_));
 sky130_fd_sc_hd__nand2b_1 _1164_ (.A_N(_0281_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2b_1 _1165_ (.A_N(_0282_),
    .B(_0281_),
    .Y(_0284_));
 sky130_fd_sc_hd__o22a_1 _1166_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0283_),
    .B1(_0284_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .X(_0285_));
 sky130_fd_sc_hd__nand2_1 _1167_ (.A(_0281_),
    .B(_0282_),
    .Y(_0286_));
 sky130_fd_sc_hd__or2_4 _1168_ (.A(_0282_),
    .B(_0281_),
    .X(_0287_));
 sky130_fd_sc_hd__o221a_1 _1169_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0286_),
    .B1(_0287_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .C1(_0285_),
    .X(_0288_));
 sky130_fd_sc_hd__mux4_2 _1170_ (.A0(_0264_),
    .A1(_0265_),
    .A2(_0256_),
    .A3(_0255_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _1171_ (.A(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .B(_0284_),
    .X(_0290_));
 sky130_fd_sc_hd__or2_1 _1172_ (.A(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .B(_0286_),
    .X(_0291_));
 sky130_fd_sc_hd__o221a_1 _1173_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0283_),
    .B1(_0287_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .C1(_0290_),
    .X(_0292_));
 sky130_fd_sc_hd__a221o_1 _1174_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0276_),
    .B1(_0291_),
    .B2(_0292_),
    .C1(_0279_),
    .X(_0293_));
 sky130_fd_sc_hd__o211ai_2 _1175_ (.A1(_0280_),
    .A2(_0288_),
    .B1(_0289_),
    .C1(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__o22a_1 _1176_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0284_),
    .B1(_0286_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .X(_0295_));
 sky130_fd_sc_hd__o22a_1 _1177_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0283_),
    .B1(_0287_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_1 _1178_ (.A(_0295_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__o22a_1 _1179_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0284_),
    .B1(_0286_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .X(_0298_));
 sky130_fd_sc_hd__o22a_1 _1180_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0283_),
    .B1(_0287_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _1181_ (.A(_0298_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__mux2_1 _1182_ (.A0(_0297_),
    .A1(_0300_),
    .S(_0280_),
    .X(_0301_));
 sky130_fd_sc_hd__o211a_1 _1183_ (.A1(_0289_),
    .A2(_0301_),
    .B1(_0574_),
    .C1(_0294_),
    .X(_0302_));
 sky130_fd_sc_hd__o21ba_4 _1184_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0574_),
    .B1_N(_0302_),
    .X(H));
 sky130_fd_sc_hd__mux2_4 _1185_ (.A0(net481),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_4 _1186_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_4 _1187_ (.A0(_0304_),
    .A1(_0303_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ),
    .X(_0305_));
 sky130_fd_sc_hd__inv_2 _1188_ (.A(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__nor2_1 _1189_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .B(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .Y(_0307_));
 sky130_fd_sc_hd__a211oi_4 _1190_ (.A1(_0027_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .B1(_0307_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_0308_));
 sky130_fd_sc_hd__mux2_4 _1191_ (.A0(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .X(_0309_));
 sky130_fd_sc_hd__a21oi_4 _1192_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ),
    .A2(_0309_),
    .B1(_0308_),
    .Y(_0310_));
 sky130_fd_sc_hd__mux2_4 _1193_ (.A0(_0306_),
    .A1(net475),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_4 _1194_ (.A0(net484),
    .A1(net646),
    .S(_0311_),
    .X(\Inst_LUT4AB_switch_matrix.M_EF ));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(_0149_),
    .A1(_0148_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _1196_ (.A0(_0138_),
    .A1(_0139_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _1197_ (.A0(_0313_),
    .A1(_0312_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_4 _1198_ (.A0(_0314_),
    .A1(_0059_),
    .S(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_1 _1199_ (.A(_0030_),
    .B(_0049_),
    .Y(_0316_));
 sky130_fd_sc_hd__or2_1 _1200_ (.A(_0030_),
    .B(_0049_),
    .X(_0317_));
 sky130_fd_sc_hd__o22a_1 _1201_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0316_),
    .B1(_0317_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .X(_0318_));
 sky130_fd_sc_hd__o221a_1 _1202_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0050_),
    .B1(_0051_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .C1(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__mux4_1 _1203_ (.A0(_0164_),
    .A1(_0165_),
    .A2(_0173_),
    .A3(_0172_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .X(_0320_));
 sky130_fd_sc_hd__or2_1 _1204_ (.A(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .B(_0051_),
    .X(_0321_));
 sky130_fd_sc_hd__o22a_1 _1205_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0316_),
    .B1(_0317_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .X(_0322_));
 sky130_fd_sc_hd__o211a_1 _1206_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0050_),
    .B1(_0321_),
    .C1(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_4 _1207_ (.A0(_0319_),
    .A1(_0323_),
    .S(_0315_),
    .X(_0324_));
 sky130_fd_sc_hd__o22a_1 _1208_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0316_),
    .B1(_0317_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .X(_0325_));
 sky130_fd_sc_hd__o221a_1 _1209_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0050_),
    .B1(_0051_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .C1(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _1210_ (.A(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .B(_0051_),
    .X(_0327_));
 sky130_fd_sc_hd__o22a_1 _1211_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0316_),
    .B1(_0317_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .X(_0328_));
 sky130_fd_sc_hd__o211a_1 _1212_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0050_),
    .B1(_0327_),
    .C1(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _1213_ (.A0(_0329_),
    .A1(_0326_),
    .S(_0315_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_4 _1214_ (.A0(_0324_),
    .A1(_0330_),
    .S(_0320_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_4 _1215_ (.A0(_0331_),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ),
    .X(D));
 sky130_fd_sc_hd__mux2_4 _1216_ (.A0(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_4 _1217_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_0333_));
 sky130_fd_sc_hd__and2b_1 _1218_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ),
    .B(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__a21oi_4 _1219_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ),
    .A2(_0332_),
    .B1(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__mux2_4 _1220_ (.A0(_0335_),
    .A1(net475),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_4 _1221_ (.A0(net640),
    .A1(net625),
    .S(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_4 _1222_ (.A0(_0337_),
    .A1(net483),
    .S(net522),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_4 _1223_ (.A0(_0337_),
    .A1(_0338_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(\Inst_LUT4AB_switch_matrix.M_AD ));
 sky130_fd_sc_hd__mux4_1 _1224_ (.A0(net656),
    .A1(net652),
    .A2(net627),
    .A3(net642),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0339_));
 sky130_fd_sc_hd__nand2b_1 _1225_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__mux4_1 _1226_ (.A0(net647),
    .A1(net632),
    .A2(net637),
    .A3(net408),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_0341_));
 sky130_fd_sc_hd__nand2_1 _1227_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__mux4_1 _1228_ (.A0(net59),
    .A1(net63),
    .A2(net2),
    .A3(net6),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0343_));
 sky130_fd_sc_hd__mux4_1 _1229_ (.A0(net87),
    .A1(net89),
    .A2(net111),
    .A3(net137),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _1230_ (.A0(_0343_),
    .A1(_0344_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_0345_));
 sky130_fd_sc_hd__nor2_1 _1231_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__a31o_1 _1232_ (.A1(_0342_),
    .A2(_0340_),
    .A3(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .B1(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__inv_4 _1233_ (.A(_0347_),
    .Y(\Inst_LUT4AB_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__mux4_2 _1234_ (.A0(net646),
    .A1(net631),
    .A2(net477),
    .A3(net417),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0348_));
 sky130_fd_sc_hd__mux4_1 _1235_ (.A0(net655),
    .A1(net650),
    .A2(net625),
    .A3(net640),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0349_));
 sky130_fd_sc_hd__and2b_1 _1236_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .B(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__a21bo_1 _1237_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A2(_0348_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0351_));
 sky130_fd_sc_hd__mux4_1 _1238_ (.A0(net59),
    .A1(net63),
    .A2(net2),
    .A3(net24),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .X(_0352_));
 sky130_fd_sc_hd__mux4_1 _1239_ (.A0(net87),
    .A1(net115),
    .A2(net91),
    .A3(net660),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _1240_ (.A0(_0352_),
    .A1(_0353_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .X(_0354_));
 sky130_fd_sc_hd__o22a_1 _1241_ (.A1(_0351_),
    .A2(_0350_),
    .B1(_0354_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG7 ));
 sky130_fd_sc_hd__mux4_1 _1242_ (.A0(net655),
    .A1(net651),
    .A2(net626),
    .A3(net640),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0355_));
 sky130_fd_sc_hd__mux4_1 _1243_ (.A0(net646),
    .A1(net631),
    .A2(net636),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _1244_ (.A0(_0355_),
    .A1(_0356_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0357_));
 sky130_fd_sc_hd__mux4_1 _1245_ (.A0(net59),
    .A1(net63),
    .A2(net2),
    .A3(net6),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0358_));
 sky130_fd_sc_hd__mux4_1 _1246_ (.A0(net87),
    .A1(net115),
    .A2(net91),
    .A3(net117),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _1247_ (.A0(_0358_),
    .A1(_0359_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_4 _1248_ (.A0(_0360_),
    .A1(_0357_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG7 ));
 sky130_fd_sc_hd__mux4_2 _1249_ (.A0(net654),
    .A1(net649),
    .A2(net624),
    .A3(net638),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0361_));
 sky130_fd_sc_hd__mux4_2 _1250_ (.A0(net464),
    .A1(net630),
    .A2(net478),
    .A3(net480),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_4 _1251_ (.A0(_0361_),
    .A1(_0362_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_0363_));
 sky130_fd_sc_hd__mux4_1 _1252_ (.A0(net59),
    .A1(net83),
    .A2(net2),
    .A3(net6),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0364_));
 sky130_fd_sc_hd__mux4_1 _1253_ (.A0(net87),
    .A1(net89),
    .A2(net91),
    .A3(net115),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _1254_ (.A0(_0364_),
    .A1(_0365_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_4 _1255_ (.A0(_0366_),
    .A1(_0363_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG7 ));
 sky130_fd_sc_hd__nand2b_1 _1256_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .B(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .Y(_0367_));
 sky130_fd_sc_hd__a21oi_1 _1257_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_0368_));
 sky130_fd_sc_hd__mux2_4 _1258_ (.A0(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_0369_));
 sky130_fd_sc_hd__a2bb2o_4 _1259_ (.A1_N(_0575_),
    .A2_N(_0369_),
    .B1(_0368_),
    .B2(_0367_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_4 _1260_ (.A0(_0370_),
    .A1(_0335_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _1261_ (.A0(_0371_),
    .A1(_0311_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _1262_ (.A0(net622),
    .A1(net631),
    .S(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_4 _1263_ (.A0(_0373_),
    .A1(net617),
    .S(_0371_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_4 _1264_ (.A0(_0373_),
    .A1(_0374_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _1265_ (.A0(_0374_),
    .A1(_0338_),
    .S(_0370_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_4 _1266_ (.A0(_0375_),
    .A1(_0376_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.M_AH ));
 sky130_fd_sc_hd__mux2_4 _1267_ (.A0(net650),
    .A1(net654),
    .S(net520),
    .X(\Inst_LUT4AB_switch_matrix.M_AB ));
 sky130_fd_sc_hd__mux4_1 _1268_ (.A0(net648),
    .A1(net638),
    .A2(net623),
    .A3(net643),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0377_));
 sky130_fd_sc_hd__or2_1 _1269_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__mux4_1 _1270_ (.A0(net633),
    .A1(net628),
    .A2(net619),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .X(_0379_));
 sky130_fd_sc_hd__o21a_1 _1271_ (.A1(_0576_),
    .A2(_0379_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0380_));
 sky130_fd_sc_hd__mux4_1 _1272_ (.A0(net62),
    .A1(net7),
    .A2(net64),
    .A3(net804),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0381_));
 sky130_fd_sc_hd__mux4_1 _1273_ (.A0(net92),
    .A1(net120),
    .A2(net108),
    .A3(net136),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _1274_ (.A0(_0381_),
    .A1(_0382_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0383_));
 sky130_fd_sc_hd__a22o_1 _1275_ (.A1(_0378_),
    .A2(_0380_),
    .B1(_0383_),
    .B2(_0577_),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1276_ (.A0(net446),
    .A1(net444),
    .A2(net463),
    .A3(net643),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0384_));
 sky130_fd_sc_hd__mux4_2 _1277_ (.A0(net633),
    .A1(net628),
    .A2(net619),
    .A3(net404),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .X(_0385_));
 sky130_fd_sc_hd__or2_4 _1278_ (.A(_0578_),
    .B(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__o21a_1 _1279_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0384_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_0387_));
 sky130_fd_sc_hd__mux4_1 _1280_ (.A0(net92),
    .A1(net120),
    .A2(net108),
    .A3(net136),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0388_));
 sky130_fd_sc_hd__mux4_1 _1281_ (.A0(net84),
    .A1(net7),
    .A2(net806),
    .A3(net804),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _1282_ (.A0(_0388_),
    .A1(_0389_),
    .S(_0578_),
    .X(_0390_));
 sky130_fd_sc_hd__a22o_1 _1283_ (.A1(_0386_),
    .A2(_0387_),
    .B1(_0390_),
    .B2(_0579_),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1284_ (.A0(net634),
    .A1(net629),
    .A2(net619),
    .A3(net416),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0391_));
 sky130_fd_sc_hd__or2_4 _1285_ (.A(_0580_),
    .B(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__mux4_1 _1286_ (.A0(net446),
    .A1(net444),
    .A2(net463),
    .A3(net643),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0393_));
 sky130_fd_sc_hd__o21a_1 _1287_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .A2(_0393_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0394_));
 sky130_fd_sc_hd__mux4_1 _1288_ (.A0(net804),
    .A1(net120),
    .A2(net92),
    .A3(net136),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .X(_0395_));
 sky130_fd_sc_hd__mux4_1 _1289_ (.A0(net62),
    .A1(net64),
    .A2(net80),
    .A3(net25),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _1290_ (.A0(_0395_),
    .A1(_0396_),
    .S(_0580_),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _1291_ (.A1(_0392_),
    .A2(_0394_),
    .B1(_0397_),
    .B2(_0581_),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1292_ (.A0(net446),
    .A1(net638),
    .A2(net623),
    .A3(net643),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .X(_0398_));
 sky130_fd_sc_hd__or2_1 _1293_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__mux4_1 _1294_ (.A0(net633),
    .A1(net628),
    .A2(net619),
    .A3(net618),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_0400_));
 sky130_fd_sc_hd__o21a_1 _1295_ (.A1(_0582_),
    .A2(_0400_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .X(_0401_));
 sky130_fd_sc_hd__mux4_1 _1296_ (.A0(net804),
    .A1(net112),
    .A2(net120),
    .A3(net136),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_0402_));
 sky130_fd_sc_hd__mux4_1 _1297_ (.A0(net64),
    .A1(net806),
    .A2(net80),
    .A3(net7),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _1298_ (.A0(_0402_),
    .A1(_0403_),
    .S(_0582_),
    .X(_0404_));
 sky130_fd_sc_hd__a22o_1 _1299_ (.A1(_0401_),
    .A2(_0399_),
    .B1(_0404_),
    .B2(_0583_),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1300_ (.A0(_0639_),
    .A1(_0046_),
    .A2(_0082_),
    .A3(_0235_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0405_));
 sky130_fd_sc_hd__nand2b_4 _1301_ (.A_N(_0405_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .Y(_0406_));
 sky130_fd_sc_hd__mux4_1 _1302_ (.A0(net628),
    .A1(net619),
    .A2(net523),
    .A3(net416),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0407_));
 sky130_fd_sc_hd__o211a_1 _1303_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0407_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .C1(_0406_),
    .X(_0408_));
 sky130_fd_sc_hd__nand2b_1 _1304_ (.A_N(net660),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .Y(_0409_));
 sky130_fd_sc_hd__o21ba_1 _1305_ (.A1(net807),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _1306_ (.A0(net433),
    .A1(net446),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_0411_));
 sky130_fd_sc_hd__a221o_1 _1307_ (.A1(_0409_),
    .A2(_0410_),
    .B1(_0411_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _1308_ (.A0(net414),
    .A1(net444),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_0413_));
 sky130_fd_sc_hd__inv_1 _1309_ (.A(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__mux2_1 _1310_ (.A0(net464),
    .A1(net415),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_0415_));
 sky130_fd_sc_hd__o21ai_1 _1311_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .A2(_0414_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .Y(_0416_));
 sky130_fd_sc_hd__a21o_1 _1312_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .A2(_0415_),
    .B1(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__a31o_1 _1313_ (.A1(_0584_),
    .A2(_0412_),
    .A3(_0417_),
    .B1(_0408_),
    .X(\Inst_LUT4AB_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1314_ (.A0(net806),
    .A1(net659),
    .A2(net654),
    .A3(net651),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0418_));
 sky130_fd_sc_hd__mux4_1 _1315_ (.A0(net626),
    .A1(net640),
    .A2(net646),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _1316_ (.A0(_0418_),
    .A1(_0419_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_0420_));
 sky130_fd_sc_hd__mux4_2 _1317_ (.A0(net631),
    .A1(net622),
    .A2(net482),
    .A3(net406),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _1318_ (.A0(_0595_),
    .A1(_0029_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_0422_));
 sky130_fd_sc_hd__and2b_1 _1319_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .B(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _1320_ (.A0(_0097_),
    .A1(net658),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_0424_));
 sky130_fd_sc_hd__a21bo_1 _1321_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .A2(_0424_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_0425_));
 sky130_fd_sc_hd__o221a_1 _1322_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_0421_),
    .B1(_0423_),
    .B2(_0425_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ),
    .X(_0426_));
 sky130_fd_sc_hd__a21o_1 _1323_ (.A1(_0585_),
    .A2(_0420_),
    .B1(_0426_),
    .X(\Inst_LUT4AB_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1324_ (.A0(net60),
    .A1(net88),
    .A2(net116),
    .A3(net445),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0427_));
 sky130_fd_sc_hd__mux4_2 _1325_ (.A0(net644),
    .A1(_0082_),
    .A2(_0235_),
    .A3(_0649_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_4 _1326_ (.A0(_0427_),
    .A1(_0428_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__mux2_1 _1327_ (.A0(net658),
    .A1(_0039_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0429_));
 sky130_fd_sc_hd__nand2_1 _1328_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__mux2_1 _1329_ (.A0(net414),
    .A1(_0097_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0431_));
 sky130_fd_sc_hd__inv_1 _1330_ (.A(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__o211a_1 _1331_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_0432_),
    .B1(_0430_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .X(_0433_));
 sky130_fd_sc_hd__mux4_1 _1332_ (.A0(net59),
    .A1(net115),
    .A2(net87),
    .A3(net446),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_0434_));
 sky130_fd_sc_hd__o21ba_1 _1333_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .A2(_0434_),
    .B1_N(_0433_),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1334_ (.A0(net62),
    .A1(net90),
    .A2(net118),
    .A3(net654),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0435_));
 sky130_fd_sc_hd__mux4_2 _1335_ (.A0(net621),
    .A1(_0639_),
    .A2(_0046_),
    .A3(_0085_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_4 _1336_ (.A0(_0435_),
    .A1(_0436_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1337_ (.A0(_0029_),
    .A1(_0238_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_0437_));
 sky130_fd_sc_hd__nand2_1 _1338_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__mux2_1 _1339_ (.A0(net630),
    .A1(_0595_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_0439_));
 sky130_fd_sc_hd__inv_1 _1340_ (.A(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__o211a_1 _1341_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .A2(_0440_),
    .B1(_0438_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .X(_0441_));
 sky130_fd_sc_hd__mux4_2 _1342_ (.A0(net61),
    .A1(net89),
    .A2(net660),
    .A3(net478),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0442_));
 sky130_fd_sc_hd__o21ba_1 _1343_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(_0442_),
    .B1_N(_0441_),
    .X(\Inst_LUT4AB_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1344_ (.A0(net60),
    .A1(net3),
    .A2(net116),
    .A3(net445),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .X(_0443_));
 sky130_fd_sc_hd__mux4_1 _1345_ (.A0(net645),
    .A1(_0082_),
    .A2(_0235_),
    .A3(_0661_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _1346_ (.A0(_0443_),
    .A1(_0444_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Inst_LUT4AB_switch_matrix.SS4BEG3 ));
 sky130_fd_sc_hd__mux2_1 _1347_ (.A0(net658),
    .A1(_0173_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_0445_));
 sky130_fd_sc_hd__nand2_1 _1348_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__mux2_1 _1349_ (.A0(net414),
    .A1(_0097_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_0447_));
 sky130_fd_sc_hd__inv_1 _1350_ (.A(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__o211a_1 _1351_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .A2(_0448_),
    .B1(_0446_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .X(_0449_));
 sky130_fd_sc_hd__mux4_1 _1352_ (.A0(net59),
    .A1(net115),
    .A2(net2),
    .A3(net649),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_0450_));
 sky130_fd_sc_hd__o21ba_1 _1353_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .A2(_0450_),
    .B1_N(_0449_),
    .X(\Inst_LUT4AB_switch_matrix.SS4BEG2 ));
 sky130_fd_sc_hd__mux2_1 _1354_ (.A0(net525),
    .A1(_0121_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_0451_));
 sky130_fd_sc_hd__nand2_1 _1355_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .B(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__nor2_1 _1356_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .B(net412),
    .Y(_0453_));
 sky130_fd_sc_hd__a211o_1 _1357_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_0638_),
    .B1(_0453_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0454_));
 sky130_fd_sc_hd__and3_1 _1358_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .B(_0452_),
    .C(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__mux4_1 _1359_ (.A0(net62),
    .A1(net806),
    .A2(net659),
    .A3(net434),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0456_));
 sky130_fd_sc_hd__o21ba_4 _1360_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .A2(_0456_),
    .B1_N(_0455_),
    .X(\Inst_LUT4AB_switch_matrix.SS4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1361_ (.A0(_0029_),
    .A1(_0256_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_1 _1362_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .B(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__mux2_1 _1363_ (.A0(net411),
    .A1(_0595_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_0459_));
 sky130_fd_sc_hd__inv_1 _1364_ (.A(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__o211a_1 _1365_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .A2(_0460_),
    .B1(_0458_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .X(_0461_));
 sky130_fd_sc_hd__mux4_1 _1366_ (.A0(net61),
    .A1(net660),
    .A2(net807),
    .A3(net415),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_0462_));
 sky130_fd_sc_hd__o21ba_1 _1367_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .A2(_0462_),
    .B1_N(_0461_),
    .X(\Inst_LUT4AB_switch_matrix.SS4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1368_ (.A0(net625),
    .A1(net641),
    .A2(net647),
    .A3(net477),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0463_));
 sky130_fd_sc_hd__mux4_1 _1369_ (.A0(net4),
    .A1(net660),
    .A2(net656),
    .A3(net651),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _1370_ (.A0(_0464_),
    .A1(_0463_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .X(_0465_));
 sky130_fd_sc_hd__mux4_1 _1371_ (.A0(_0639_),
    .A1(_0046_),
    .A2(_0082_),
    .A3(_0235_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0466_));
 sky130_fd_sc_hd__mux4_2 _1372_ (.A0(net630),
    .A1(net622),
    .A2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .A3(net416),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_4 _1373_ (.A0(_0467_),
    .A1(_0466_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_4 _1374_ (.A0(_0465_),
    .A1(_0468_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1375_ (.A0(net806),
    .A1(net659),
    .A2(net656),
    .A3(net651),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0469_));
 sky130_fd_sc_hd__mux4_1 _1376_ (.A0(net627),
    .A1(net642),
    .A2(net647),
    .A3(net636),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _1377_ (.A0(_0469_),
    .A1(_0470_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .X(_0471_));
 sky130_fd_sc_hd__mux4_2 _1378_ (.A0(net632),
    .A1(net622),
    .A2(net482),
    .A3(net408),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _1379_ (.A0(_0595_),
    .A1(_0029_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .X(_0473_));
 sky130_fd_sc_hd__and2b_1 _1380_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .B(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _1381_ (.A0(_0097_),
    .A1(net658),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .X(_0475_));
 sky130_fd_sc_hd__a21bo_1 _1382_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_0475_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .X(_0476_));
 sky130_fd_sc_hd__o221a_1 _1383_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .A2(_0472_),
    .B1(_0474_),
    .B2(_0476_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ),
    .X(_0477_));
 sky130_fd_sc_hd__a21o_1 _1384_ (.A1(_0586_),
    .A2(_0471_),
    .B1(_0477_),
    .X(\Inst_LUT4AB_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1385_ (.A0(net60),
    .A1(net3),
    .A2(net88),
    .A3(net642),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_4 _1386_ (.A0(net647),
    .A1(_0082_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_4 _1387_ (.A0(_0235_),
    .A1(_0625_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_4 _1388_ (.A0(_0479_),
    .A1(_0480_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_4 _1389_ (.A0(_0478_),
    .A1(_0481_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .X(\Inst_LUT4AB_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__mux2_1 _1390_ (.A0(net658),
    .A1(_0149_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _1391_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__mux2_1 _1392_ (.A0(net627),
    .A1(_0097_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .X(_0484_));
 sky130_fd_sc_hd__inv_1 _1393_ (.A(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__o211a_1 _1394_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .A2(_0485_),
    .B1(_0483_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .X(_0486_));
 sky130_fd_sc_hd__mux4_1 _1395_ (.A0(net59),
    .A1(net87),
    .A2(net2),
    .A3(net651),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .X(_0487_));
 sky130_fd_sc_hd__o21ba_1 _1396_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .A2(_0487_),
    .B1_N(_0486_),
    .X(\Inst_LUT4AB_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1397_ (.A0(net62),
    .A1(net806),
    .A2(net90),
    .A3(net656),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .X(_0488_));
 sky130_fd_sc_hd__nor2_1 _1398_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .B(net622),
    .Y(_0489_));
 sky130_fd_sc_hd__a211oi_1 _1399_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .A2(_0638_),
    .B1(_0489_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .Y(_0490_));
 sky130_fd_sc_hd__mux2_1 _1400_ (.A0(net525),
    .A1(_0070_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .X(_0491_));
 sky130_fd_sc_hd__a21bo_1 _1401_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .A2(_0491_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .X(_0492_));
 sky130_fd_sc_hd__o22a_4 _1402_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .A2(_0488_),
    .B1(_0490_),
    .B2(_0492_),
    .X(\Inst_LUT4AB_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1403_ (.A0(_0029_),
    .A1(_0224_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .X(_0493_));
 sky130_fd_sc_hd__nand2_1 _1404_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__mux2_1 _1405_ (.A0(net632),
    .A1(_0595_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .X(_0495_));
 sky130_fd_sc_hd__inv_1 _1406_ (.A(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__o211a_1 _1407_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .A2(_0496_),
    .B1(_0494_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _1408_ (.A0(net61),
    .A1(net807),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .X(_0498_));
 sky130_fd_sc_hd__nand2b_1 _1409_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .B(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__mux2_1 _1410_ (.A0(net89),
    .A1(net477),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .X(_0500_));
 sky130_fd_sc_hd__a21oi_1 _1411_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .A2(_0500_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .Y(_0501_));
 sky130_fd_sc_hd__a21oi_1 _1412_ (.A1(_0499_),
    .A2(_0501_),
    .B1(_0497_),
    .Y(\Inst_LUT4AB_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1413_ (.A0(net60),
    .A1(net3),
    .A2(net116),
    .A3(net642),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .X(_0502_));
 sky130_fd_sc_hd__mux4_2 _1414_ (.A0(net647),
    .A1(_0082_),
    .A2(_0235_),
    .A3(_0604_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_4 _1415_ (.A0(_0502_),
    .A1(_0503_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.NN4BEG3 ));
 sky130_fd_sc_hd__mux2_1 _1416_ (.A0(net658),
    .A1(_0019_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_1 _1417_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__mux2_1 _1418_ (.A0(net627),
    .A1(_0097_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .X(_0506_));
 sky130_fd_sc_hd__inv_1 _1419_ (.A(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__o211a_1 _1420_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .A2(_0507_),
    .B1(_0505_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _1421_ (.A0(net59),
    .A1(net2),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .X(_0509_));
 sky130_fd_sc_hd__nand2b_1 _1422_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .B(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__mux2_1 _1423_ (.A0(net115),
    .A1(net651),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .X(_0511_));
 sky130_fd_sc_hd__a21oi_1 _1424_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .A2(_0511_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .Y(_0512_));
 sky130_fd_sc_hd__a21oi_1 _1425_ (.A1(_0510_),
    .A2(_0512_),
    .B1(_0508_),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1426_ (.A0(net62),
    .A1(net806),
    .A2(net659),
    .A3(net656),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .X(_0513_));
 sky130_fd_sc_hd__nor2_1 _1427_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .B(net622),
    .Y(_0514_));
 sky130_fd_sc_hd__a211oi_1 _1428_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .A2(_0638_),
    .B1(_0514_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .Y(_0515_));
 sky130_fd_sc_hd__mux2_1 _1429_ (.A0(net525),
    .A1(_0088_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .X(_0516_));
 sky130_fd_sc_hd__a21bo_1 _1430_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .A2(_0516_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ),
    .X(_0517_));
 sky130_fd_sc_hd__o22a_1 _1431_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ),
    .A2(_0513_),
    .B1(_0515_),
    .B2(_0517_),
    .X(\Inst_LUT4AB_switch_matrix.NN4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(_0029_),
    .A1(_0249_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .X(_0518_));
 sky130_fd_sc_hd__nand2_1 _1433_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__mux2_1 _1434_ (.A0(net632),
    .A1(_0595_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .X(_0520_));
 sky130_fd_sc_hd__inv_1 _1435_ (.A(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__o211a_1 _1436_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .A2(_0521_),
    .B1(_0519_),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .X(_0522_));
 sky130_fd_sc_hd__mux4_1 _1437_ (.A0(net61),
    .A1(net660),
    .A2(net807),
    .A3(net477),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .X(_0523_));
 sky130_fd_sc_hd__o21ba_1 _1438_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .A2(_0523_),
    .B1_N(_0522_),
    .X(\Inst_LUT4AB_switch_matrix.NN4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1439_ (.A0(net434),
    .A1(_0640_),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A3(_0624_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1440_ (.A0(net619),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .A2(net658),
    .A3(_0255_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1441_ (.A0(net628),
    .A1(_0068_),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .A3(_0084_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1442_ (.A0(net462),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .A2(_0165_),
    .A3(_0018_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1443_ (.A0(net92),
    .A1(net107),
    .A2(net135),
    .A3(net445),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_1 _1444_ (.A0(net91),
    .A1(net136),
    .A2(net110),
    .A3(net414),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1445_ (.A0(net805),
    .A1(net109),
    .A2(net94),
    .A3(net649),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1446_ (.A0(net804),
    .A1(net108),
    .A2(net93),
    .A3(net433),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1447_ (.A0(net412),
    .A1(_0640_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .A3(_0624_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1448_ (.A0(net411),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .A2(net658),
    .A3(_0255_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1449_ (.A0(net415),
    .A1(_0068_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .A3(_0084_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1450_ (.A0(net643),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .A2(_0165_),
    .A3(_0018_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1451_ (.A0(net411),
    .A1(_0640_),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A3(_0624_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1452_ (.A0(net415),
    .A1(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .A2(net658),
    .A3(_0255_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1453_ (.A0(net645),
    .A1(_0068_),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .A3(_0084_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1454_ (.A0(net445),
    .A1(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .A2(_0165_),
    .A3(_0018_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__mux4_1 _1455_ (.A0(net64),
    .A1(net135),
    .A2(net79),
    .A3(net412),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1456_ (.A0(net63),
    .A1(net82),
    .A2(net136),
    .A3(net631),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__mux4_2 _1457_ (.A0(net66),
    .A1(net81),
    .A2(net805),
    .A3(net478),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__mux4_1 _1458_ (.A0(net65),
    .A1(net80),
    .A2(net804),
    .A3(net464),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__mux4_2 _1459_ (.A0(net637),
    .A1(_0640_),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .A3(_0624_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_2 _1460_ (.A0(net464),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .A2(net658),
    .A3(_0255_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _1461_ (.A0(net641),
    .A1(_0068_),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .A3(_0084_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux4_2 _1462_ (.A0(net463),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .A2(_0165_),
    .A3(_0018_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__a21bo_4 _1463_ (.A1(_0287_),
    .A2(_0276_),
    .B1_N(_0286_),
    .X(net141));
 sky130_fd_sc_hd__mux2_1 _1464_ (.A0(_0264_),
    .A1(_0670_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(_0165_),
    .A1(_0119_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0525_));
 sky130_fd_sc_hd__mux4_2 _1466_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(_0524_),
    .A1(_0525_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_0527_));
 sky130_fd_sc_hd__and2b_1 _1468_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .B(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__a21oi_4 _1469_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0526_),
    .B1(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__or2_1 _1470_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .B(_0221_),
    .X(_0530_));
 sky130_fd_sc_hd__a21oi_1 _1471_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_0615_),
    .B1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0531_));
 sky130_fd_sc_hd__mux2_1 _1472_ (.A0(_0139_),
    .A1(_0068_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0532_));
 sky130_fd_sc_hd__a221o_1 _1473_ (.A1(_0530_),
    .A2(_0531_),
    .B1(_0532_),
    .B2(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .C1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_2 _1474_ (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0534_));
 sky130_fd_sc_hd__and2b_1 _1475_ (.A_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .B(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _1476_ (.A0(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_0536_));
 sky130_fd_sc_hd__a21bo_1 _1477_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_0536_),
    .B1_N(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .X(_0537_));
 sky130_fd_sc_hd__o21a_4 _1478_ (.A1(_0537_),
    .A2(_0535_),
    .B1(_0533_),
    .X(_0538_));
 sky130_fd_sc_hd__nand2_2 _1479_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__o211ai_1 _1480_ (.A1(_0289_),
    .A2(_0301_),
    .B1(_0539_),
    .C1(_0294_),
    .Y(_0540_));
 sky130_fd_sc_hd__o2bb2a_1 _1481_ (.A1_N(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2_N(_0529_),
    .B1(_0539_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ),
    .X(_0541_));
 sky130_fd_sc_hd__a32o_1 _1482_ (.A1(net548),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A3(_0529_),
    .B1(_0540_),
    .B2(_0541_),
    .X(_0000_));
 sky130_fd_sc_hd__nand2_2 _1483_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ),
    .B(_0538_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_1 _1484_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ),
    .B(_0529_),
    .Y(_0543_));
 sky130_fd_sc_hd__mux2_2 _1485_ (.A0(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0685_),
    .S(_0542_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(net546),
    .A1(_0544_),
    .S(_0543_),
    .X(_0001_));
 sky130_fd_sc_hd__nand2_1 _1487_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .B(_0529_),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_4 _1488_ (.A(_0538_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ),
    .Y(_0546_));
 sky130_fd_sc_hd__mux2_2 _1489_ (.A0(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0011_),
    .S(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _1490_ (.A0(net545),
    .A1(_0547_),
    .S(_0545_),
    .X(_0002_));
 sky130_fd_sc_hd__nand2_1 _1491_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .B(_0529_),
    .Y(_0548_));
 sky130_fd_sc_hd__nand2_2 _1492_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ),
    .B(_0538_),
    .Y(_0549_));
 sky130_fd_sc_hd__mux2_2 _1493_ (.A0(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0186_),
    .S(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _1494_ (.A0(net544),
    .A1(_0550_),
    .S(_0548_),
    .X(_0003_));
 sky130_fd_sc_hd__nand2_1 _1495_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .B(_0529_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_4 _1496_ (.A(_0538_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ),
    .Y(_0552_));
 sky130_fd_sc_hd__mux2_2 _1497_ (.A0(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0331_),
    .S(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _1498_ (.A0(net542),
    .A1(_0553_),
    .S(_0551_),
    .X(_0004_));
 sky130_fd_sc_hd__nand2_1 _1499_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .B(_0529_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_4 _1500_ (.A(_0538_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ),
    .Y(_0555_));
 sky130_fd_sc_hd__mux2_2 _1501_ (.A0(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0131_),
    .S(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _1502_ (.A0(net541),
    .A1(_0556_),
    .S(_0554_),
    .X(_0005_));
 sky130_fd_sc_hd__nand2_1 _1503_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .B(_0529_),
    .Y(_0557_));
 sky130_fd_sc_hd__nand2_4 _1504_ (.A(_0538_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ),
    .Y(_0558_));
 sky130_fd_sc_hd__mux2_2 _1505_ (.A0(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0213_),
    .S(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_2 _1506_ (.A0(net547),
    .A1(_0559_),
    .S(_0557_),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _1507_ (.A(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .B(_0529_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_4 _1508_ (.A(_0538_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_0561_));
 sky130_fd_sc_hd__mux2_2 _1509_ (.A0(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ),
    .A1(_0275_),
    .S(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _1510_ (.A0(net543),
    .A1(_0562_),
    .S(_0560_),
    .X(_0007_));
 sky130_fd_sc_hd__dlxtp_1 _1511_ (.D(net770),
    .GATE(net56),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1512_ (.D(net769),
    .GATE(net56),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1513_ (.D(net766),
    .GATE(net56),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1514_ (.D(net764),
    .GATE(net56),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1515_ (.D(net762),
    .GATE(net56),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1516_ (.D(net760),
    .GATE(net56),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1517_ (.D(net757),
    .GATE(net56),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1518_ (.D(net755),
    .GATE(net56),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1519_ (.D(net803),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1520_ (.D(net781),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1521_ (.D(net759),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1522_ (.D(net753),
    .GATE(net700),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1523_ (.D(net751),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1524_ (.D(net749),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1525_ (.D(net747),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1526_ (.D(net745),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1527_ (.D(net743),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1528_ (.D(net740),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1529_ (.D(net800),
    .GATE(net701),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1530_ (.D(net798),
    .GATE(net700),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1531_ (.D(net796),
    .GATE(net702),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1532_ (.D(net794),
    .GATE(net702),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1533_ (.D(net792),
    .GATE(net702),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1534_ (.D(net790),
    .GATE(net700),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1535_ (.D(net788),
    .GATE(net703),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1536_ (.D(net787),
    .GATE(net703),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1537_ (.D(net784),
    .GATE(net700),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1538_ (.D(net782),
    .GATE(net700),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1539_ (.D(net778),
    .GATE(net700),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1540_ (.D(net776),
    .GATE(net702),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1541_ (.D(net775),
    .GATE(net702),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1542_ (.D(net773),
    .GATE(net702),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1543_ (.D(net770),
    .GATE(net702),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1544_ (.D(net769),
    .GATE(net700),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1545_ (.D(net766),
    .GATE(net700),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1546_ (.D(net764),
    .GATE(net700),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1547_ (.D(net762),
    .GATE(net702),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1548_ (.D(net760),
    .GATE(net700),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1549_ (.D(net757),
    .GATE(net703),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1550_ (.D(net755),
    .GATE(net702),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1551_ (.D(net802),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1552_ (.D(net781),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1553_ (.D(net759),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1554_ (.D(net752),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1555_ (.D(net751),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1556_ (.D(net748),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1557_ (.D(net747),
    .GATE(net705),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1558_ (.D(net745),
    .GATE(net705),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1559_ (.D(net743),
    .GATE(net705),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1560_ (.D(net740),
    .GATE(net705),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1561_ (.D(net800),
    .GATE(net705),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1562_ (.D(net798),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1563_ (.D(net796),
    .GATE(net705),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1564_ (.D(net794),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1565_ (.D(net792),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1566_ (.D(net790),
    .GATE(net705),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1567_ (.D(net788),
    .GATE(net704),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1568_ (.D(net787),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1569_ (.D(net784),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1570_ (.D(net782),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1571_ (.D(net778),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1572_ (.D(net776),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1573_ (.D(net775),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1574_ (.D(net773),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1575_ (.D(net770),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1576_ (.D(net769),
    .GATE(net707),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1577_ (.D(net43),
    .GATE(net707),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1578_ (.D(net765),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1579_ (.D(net763),
    .GATE(net707),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1580_ (.D(net761),
    .GATE(net706),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1581_ (.D(net48),
    .GATE(net707),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1582_ (.D(net49),
    .GATE(net707),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1583_ (.D(net803),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1584_ (.D(net781),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1585_ (.D(net758),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1586_ (.D(net752),
    .GATE(net709),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1587_ (.D(net751),
    .GATE(net710),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1588_ (.D(net749),
    .GATE(net709),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1589_ (.D(net747),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1590_ (.D(net745),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1591_ (.D(net743),
    .GATE(net710),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1592_ (.D(net740),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1593_ (.D(net800),
    .GATE(net709),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1594_ (.D(net798),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1595_ (.D(net796),
    .GATE(net710),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1596_ (.D(net794),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1597_ (.D(net792),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1598_ (.D(net790),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1599_ (.D(net788),
    .GATE(net710),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1600_ (.D(net787),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1601_ (.D(net784),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1602_ (.D(net782),
    .GATE(net708),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1603_ (.D(net778),
    .GATE(net710),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1604_ (.D(net776),
    .GATE(net709),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1605_ (.D(net775),
    .GATE(net710),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1606_ (.D(net773),
    .GATE(net711),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1607_ (.D(net770),
    .GATE(net711),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1608_ (.D(net769),
    .GATE(net711),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1609_ (.D(net766),
    .GATE(net711),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1610_ (.D(net764),
    .GATE(net711),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1611_ (.D(net763),
    .GATE(net710),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1612_ (.D(net760),
    .GATE(net710),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1613_ (.D(net757),
    .GATE(net710),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1614_ (.D(net49),
    .GATE(net710),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1615_ (.D(net803),
    .GATE(net712),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1616_ (.D(net38),
    .GATE(net712),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1617_ (.D(net47),
    .GATE(net712),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1618_ (.D(net753),
    .GATE(net712),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1619_ (.D(net751),
    .GATE(net712),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1620_ (.D(net749),
    .GATE(net712),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1621_ (.D(net747),
    .GATE(net712),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1622_ (.D(net745),
    .GATE(net712),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1623_ (.D(net743),
    .GATE(net55),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1624_ (.D(net740),
    .GATE(net712),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1625_ (.D(net800),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1626_ (.D(net798),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1627_ (.D(net796),
    .GATE(net714),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1628_ (.D(net794),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1629_ (.D(net792),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1630_ (.D(net790),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1631_ (.D(net788),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1632_ (.D(net787),
    .GATE(net715),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1633_ (.D(net784),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1634_ (.D(net782),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1635_ (.D(net778),
    .GATE(net714),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1636_ (.D(net776),
    .GATE(net714),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1637_ (.D(net775),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1638_ (.D(net773),
    .GATE(net714),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1639_ (.D(net770),
    .GATE(net714),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1640_ (.D(net769),
    .GATE(net713),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1641_ (.D(net766),
    .GATE(net715),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1642_ (.D(net44),
    .GATE(net712),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1643_ (.D(net45),
    .GATE(net715),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1644_ (.D(net46),
    .GATE(net715),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ));
 sky130_fd_sc_hd__dlxtp_1 _1645_ (.D(net757),
    .GATE(net715),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ));
 sky130_fd_sc_hd__dlxtp_1 _1646_ (.D(net755),
    .GATE(net715),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ));
 sky130_fd_sc_hd__dlxtp_1 _1647_ (.D(net803),
    .GATE(net719),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ));
 sky130_fd_sc_hd__dlxtp_1 _1648_ (.D(net781),
    .GATE(net719),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ));
 sky130_fd_sc_hd__dlxtp_1 _1649_ (.D(net758),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ));
 sky130_fd_sc_hd__dlxtp_1 _1650_ (.D(net753),
    .GATE(net719),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ));
 sky130_fd_sc_hd__dlxtp_1 _1651_ (.D(net751),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ));
 sky130_fd_sc_hd__dlxtp_1 _1652_ (.D(net749),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ));
 sky130_fd_sc_hd__dlxtp_1 _1653_ (.D(net747),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ));
 sky130_fd_sc_hd__dlxtp_1 _1654_ (.D(net745),
    .GATE(net719),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ));
 sky130_fd_sc_hd__dlxtp_1 _1655_ (.D(net743),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ));
 sky130_fd_sc_hd__dlxtp_1 _1656_ (.D(net740),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ));
 sky130_fd_sc_hd__dlxtp_1 _1657_ (.D(net800),
    .GATE(net719),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ));
 sky130_fd_sc_hd__dlxtp_1 _1658_ (.D(net798),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ));
 sky130_fd_sc_hd__dlxtp_1 _1659_ (.D(net796),
    .GATE(net719),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ));
 sky130_fd_sc_hd__dlxtp_1 _1660_ (.D(net794),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ));
 sky130_fd_sc_hd__dlxtp_1 _1661_ (.D(net792),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ));
 sky130_fd_sc_hd__dlxtp_1 _1662_ (.D(net790),
    .GATE(net718),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ));
 sky130_fd_sc_hd__dlxtp_1 _1663_ (.D(net789),
    .GATE(net717),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1664_ (.D(net786),
    .GATE(net717),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1665_ (.D(net785),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1666_ (.D(net783),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1667_ (.D(net779),
    .GATE(net717),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1668_ (.D(net777),
    .GATE(net717),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1669_ (.D(net774),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1670_ (.D(net772),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1671_ (.D(net771),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1672_ (.D(net768),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1673_ (.D(net767),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1674_ (.D(net765),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1675_ (.D(net763),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1676_ (.D(net761),
    .GATE(net716),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1677_ (.D(net757),
    .GATE(net717),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1678_ (.D(net755),
    .GATE(net717),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1679_ (.D(net802),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1680_ (.D(net780),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1681_ (.D(net758),
    .GATE(net723),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1682_ (.D(net753),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1683_ (.D(net751),
    .GATE(net723),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1684_ (.D(net749),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1685_ (.D(net746),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1686_ (.D(net744),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1687_ (.D(net742),
    .GATE(net723),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1688_ (.D(net741),
    .GATE(net723),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1689_ (.D(net801),
    .GATE(net723),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1690_ (.D(net799),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1691_ (.D(net797),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1692_ (.D(net795),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1693_ (.D(net792),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1694_ (.D(net790),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1695_ (.D(net788),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1696_ (.D(net787),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1697_ (.D(net784),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1698_ (.D(net782),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1699_ (.D(net778),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1700_ (.D(net776),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1701_ (.D(net775),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1702_ (.D(net773),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1703_ (.D(net770),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1704_ (.D(net768),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1705_ (.D(net767),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1706_ (.D(net765),
    .GATE(net722),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1707_ (.D(net762),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1708_ (.D(net46),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1709_ (.D(net48),
    .GATE(net720),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1710_ (.D(net755),
    .GATE(net721),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1711_ (.D(net803),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1712_ (.D(net781),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1713_ (.D(net758),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1714_ (.D(net753),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1715_ (.D(net751),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1716_ (.D(net749),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1717_ (.D(net746),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1718_ (.D(net744),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1719_ (.D(net742),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1720_ (.D(net741),
    .GATE(net727),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1721_ (.D(net801),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1722_ (.D(net799),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1723_ (.D(net797),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1724_ (.D(net795),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1725_ (.D(net793),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1726_ (.D(net791),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1727_ (.D(net789),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1728_ (.D(net786),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1729_ (.D(net784),
    .GATE(net725),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1730_ (.D(net782),
    .GATE(net725),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1731_ (.D(net778),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1732_ (.D(net776),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1733_ (.D(net775),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1734_ (.D(net773),
    .GATE(net726),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1735_ (.D(net770),
    .GATE(net725),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1736_ (.D(net42),
    .GATE(net725),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1737_ (.D(net766),
    .GATE(net725),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1738_ (.D(net764),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1739_ (.D(net762),
    .GATE(net725),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1740_ (.D(net761),
    .GATE(net725),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1741_ (.D(net756),
    .GATE(net724),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1742_ (.D(net754),
    .GATE(net725),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1743_ (.D(net802),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1744_ (.D(net780),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1745_ (.D(net759),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1746_ (.D(net752),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1747_ (.D(net750),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1748_ (.D(net748),
    .GATE(net730),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1749_ (.D(net746),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1750_ (.D(net744),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1751_ (.D(net742),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1752_ (.D(net741),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1753_ (.D(net801),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1754_ (.D(net799),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1755_ (.D(net797),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1756_ (.D(net795),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1757_ (.D(net793),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1758_ (.D(net791),
    .GATE(net729),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1759_ (.D(net789),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1760_ (.D(net786),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1761_ (.D(net785),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1762_ (.D(net783),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1763_ (.D(net779),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1764_ (.D(net777),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1765_ (.D(net774),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1766_ (.D(net772),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1767_ (.D(net771),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1768_ (.D(net768),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1769_ (.D(net767),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1770_ (.D(net765),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1771_ (.D(net763),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1772_ (.D(net761),
    .GATE(net731),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1773_ (.D(net756),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1774_ (.D(net754),
    .GATE(net728),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1775_ (.D(net28),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1776_ (.D(net780),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1777_ (.D(net759),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1778_ (.D(net752),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1779_ (.D(net750),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1780_ (.D(net748),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1781_ (.D(net747),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1782_ (.D(net744),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1783_ (.D(net742),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1784_ (.D(net740),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1785_ (.D(net800),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1786_ (.D(net798),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1787_ (.D(net796),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1788_ (.D(net794),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1789_ (.D(net792),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1790_ (.D(net790),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1791_ (.D(net788),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1792_ (.D(net786),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1793_ (.D(net785),
    .GATE(net735),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1794_ (.D(net782),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1795_ (.D(net778),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1796_ (.D(net776),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1797_ (.D(net775),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1798_ (.D(net773),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1799_ (.D(net41),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1800_ (.D(net769),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1801_ (.D(net766),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1802_ (.D(net764),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1803_ (.D(net762),
    .GATE(net734),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1804_ (.D(net760),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1805_ (.D(net757),
    .GATE(net733),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1806_ (.D(net755),
    .GATE(net732),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1807_ (.D(net803),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1808_ (.D(net781),
    .GATE(net663),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1809_ (.D(net758),
    .GATE(net663),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1810_ (.D(net752),
    .GATE(net58),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1811_ (.D(net750),
    .GATE(net58),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1812_ (.D(net748),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1813_ (.D(net747),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1814_ (.D(net53),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1815_ (.D(net743),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1816_ (.D(net54),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1817_ (.D(net800),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1818_ (.D(net798),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1819_ (.D(net796),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1820_ (.D(net794),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1821_ (.D(net792),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1822_ (.D(net34),
    .GATE(net663),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1823_ (.D(net788),
    .GATE(net663),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1824_ (.D(net787),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1825_ (.D(net784),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1826_ (.D(net782),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1827_ (.D(net778),
    .GATE(net664),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1828_ (.D(net776),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1829_ (.D(net775),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1830_ (.D(net773),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1831_ (.D(net770),
    .GATE(net662),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1832_ (.D(net42),
    .GATE(net663),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1833_ (.D(net767),
    .GATE(net663),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1834_ (.D(net764),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1835_ (.D(net762),
    .GATE(net661),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1836_ (.D(net760),
    .GATE(net664),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1837_ (.D(net757),
    .GATE(net664),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1838_ (.D(net755),
    .GATE(net664),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1839_ (.D(net803),
    .GATE(net665),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1840_ (.D(net781),
    .GATE(net665),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1841_ (.D(net758),
    .GATE(net665),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1842_ (.D(net50),
    .GATE(net666),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1843_ (.D(net51),
    .GATE(net666),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1844_ (.D(net748),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1845_ (.D(net747),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1846_ (.D(net745),
    .GATE(net666),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1847_ (.D(net743),
    .GATE(net665),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1848_ (.D(net740),
    .GATE(net665),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1849_ (.D(net29),
    .GATE(net665),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1850_ (.D(net798),
    .GATE(net665),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1851_ (.D(net796),
    .GATE(net665),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1852_ (.D(net794),
    .GATE(net666),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1853_ (.D(net792),
    .GATE(net666),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1854_ (.D(net790),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1855_ (.D(net788),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1856_ (.D(net787),
    .GATE(net665),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1857_ (.D(net785),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1858_ (.D(net783),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1859_ (.D(net779),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1860_ (.D(net777),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1861_ (.D(net774),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1862_ (.D(net772),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1863_ (.D(net771),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1864_ (.D(net768),
    .GATE(net667),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1865_ (.D(net766),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1866_ (.D(net764),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1867_ (.D(net762),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1868_ (.D(net760),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1869_ (.D(net756),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1870_ (.D(net754),
    .GATE(net668),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1871_ (.D(net802),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1872_ (.D(net780),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1873_ (.D(net758),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1874_ (.D(net753),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1875_ (.D(net750),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1876_ (.D(net749),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1877_ (.D(net746),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1878_ (.D(net745),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1879_ (.D(net742),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1880_ (.D(net741),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1881_ (.D(net801),
    .GATE(net673),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1882_ (.D(net799),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1883_ (.D(net31),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1884_ (.D(net32),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1885_ (.D(net793),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1886_ (.D(net791),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1887_ (.D(net789),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1888_ (.D(net786),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1889_ (.D(net784),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1890_ (.D(net37),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1891_ (.D(net39),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1892_ (.D(net40),
    .GATE(net672),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1893_ (.D(net774),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1894_ (.D(net772),
    .GATE(net670),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1895_ (.D(net771),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1896_ (.D(net768),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1897_ (.D(net766),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1898_ (.D(net764),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1899_ (.D(net762),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1900_ (.D(net760),
    .GATE(net669),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1901_ (.D(net757),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1902_ (.D(net754),
    .GATE(net671),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1903_ (.D(net802),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1904_ (.D(net781),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1905_ (.D(net759),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1906_ (.D(net752),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1907_ (.D(net750),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1908_ (.D(net748),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1909_ (.D(net747),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1910_ (.D(net745),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1911_ (.D(net743),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1912_ (.D(net740),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1913_ (.D(net800),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1914_ (.D(net798),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1915_ (.D(net796),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1916_ (.D(net794),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1917_ (.D(net33),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1918_ (.D(net790),
    .GATE(net676),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1919_ (.D(net788),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1920_ (.D(net787),
    .GATE(net677),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1921_ (.D(net784),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1922_ (.D(net782),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1923_ (.D(net778),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1924_ (.D(net776),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1925_ (.D(net775),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1926_ (.D(net773),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1927_ (.D(net770),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1928_ (.D(net769),
    .GATE(net674),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1929_ (.D(net766),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1930_ (.D(net44),
    .GATE(net675),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1931_ (.D(net763),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1932_ (.D(net761),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1933_ (.D(net756),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1934_ (.D(net754),
    .GATE(net678),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1935_ (.D(net803),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1936_ (.D(net780),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1937_ (.D(net758),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1938_ (.D(net752),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1939_ (.D(net750),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1940_ (.D(net748),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1941_ (.D(net746),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1942_ (.D(net744),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1943_ (.D(net742),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1944_ (.D(net741),
    .GATE(net681),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1945_ (.D(net800),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1946_ (.D(net30),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1947_ (.D(net797),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1948_ (.D(net795),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1949_ (.D(net793),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1950_ (.D(net791),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1951_ (.D(net789),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1952_ (.D(net786),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1953_ (.D(net785),
    .GATE(net57),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1954_ (.D(net783),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1955_ (.D(net779),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1956_ (.D(net777),
    .GATE(net682),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1957_ (.D(net774),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1958_ (.D(net772),
    .GATE(net680),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1959_ (.D(net771),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1960_ (.D(net768),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1961_ (.D(net767),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1962_ (.D(net765),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1963_ (.D(net763),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1964_ (.D(net761),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1965_ (.D(net756),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1966_ (.D(net754),
    .GATE(net679),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1967_ (.D(net802),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1968_ (.D(net780),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1969_ (.D(net758),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1970_ (.D(net753),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1971_ (.D(net751),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1972_ (.D(net749),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1973_ (.D(net746),
    .GATE(net686),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1974_ (.D(net744),
    .GATE(net686),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1975_ (.D(net742),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1976_ (.D(net741),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1977_ (.D(net801),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1978_ (.D(net799),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1979_ (.D(net797),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1980_ (.D(net795),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1981_ (.D(net793),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1982_ (.D(net791),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1983_ (.D(net789),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1984_ (.D(net786),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1985_ (.D(net785),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1986_ (.D(net783),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1987_ (.D(net779),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1988_ (.D(net777),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1989_ (.D(net774),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1990_ (.D(net772),
    .GATE(net684),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1991_ (.D(net771),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1992_ (.D(net768),
    .GATE(net685),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1993_ (.D(net767),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1994_ (.D(net765),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1995_ (.D(net763),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1996_ (.D(net761),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1997_ (.D(net756),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1998_ (.D(net754),
    .GATE(net683),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _1999_ (.D(net802),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2000_ (.D(net780),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2001_ (.D(net759),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2002_ (.D(net752),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2003_ (.D(net750),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2004_ (.D(net52),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2005_ (.D(net746),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2006_ (.D(net744),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2007_ (.D(net742),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2008_ (.D(net741),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2009_ (.D(net801),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2010_ (.D(net799),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2011_ (.D(net797),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2012_ (.D(net795),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2013_ (.D(net793),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2014_ (.D(net791),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2015_ (.D(net35),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2016_ (.D(net787),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2017_ (.D(net785),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2018_ (.D(net783),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2019_ (.D(net779),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2020_ (.D(net777),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2021_ (.D(net774),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2022_ (.D(net772),
    .GATE(net689),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2023_ (.D(net771),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2024_ (.D(net768),
    .GATE(net690),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2025_ (.D(net767),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2026_ (.D(net765),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2027_ (.D(net763),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2028_ (.D(net761),
    .GATE(net687),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2029_ (.D(net756),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2030_ (.D(net754),
    .GATE(net688),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2031_ (.D(net802),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2032_ (.D(net780),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2033_ (.D(net759),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2034_ (.D(net752),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2035_ (.D(net750),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2036_ (.D(net748),
    .GATE(net692),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2037_ (.D(net746),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2038_ (.D(net744),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2039_ (.D(net742),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2040_ (.D(net741),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2041_ (.D(net801),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2042_ (.D(net799),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2043_ (.D(net797),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2044_ (.D(net795),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2045_ (.D(net793),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2046_ (.D(net791),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2047_ (.D(net789),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2048_ (.D(net786),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2049_ (.D(net785),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2050_ (.D(net783),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2051_ (.D(net779),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2052_ (.D(net777),
    .GATE(net694),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2053_ (.D(net774),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2054_ (.D(net772),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2055_ (.D(net771),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2056_ (.D(net769),
    .GATE(net693),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2057_ (.D(net767),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2058_ (.D(net765),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2059_ (.D(net763),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2060_ (.D(net761),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2061_ (.D(net756),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2062_ (.D(net754),
    .GATE(net691),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2063_ (.D(net802),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2064_ (.D(net780),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2065_ (.D(net759),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2066_ (.D(net752),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2067_ (.D(net750),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2068_ (.D(net748),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2069_ (.D(net746),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2070_ (.D(net744),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2071_ (.D(net742),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2072_ (.D(net741),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2073_ (.D(net801),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2074_ (.D(net799),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2075_ (.D(net797),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2076_ (.D(net795),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2077_ (.D(net793),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2078_ (.D(net791),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2079_ (.D(net789),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2080_ (.D(net786),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2081_ (.D(net785),
    .GATE(net699),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2082_ (.D(net783),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2083_ (.D(net779),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2084_ (.D(net777),
    .GATE(net698),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2085_ (.D(net774),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2086_ (.D(net772),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2087_ (.D(net771),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2088_ (.D(net768),
    .GATE(net696),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2089_ (.D(net767),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2090_ (.D(net765),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2091_ (.D(net762),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2092_ (.D(net760),
    .GATE(net697),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2093_ (.D(net756),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2094_ (.D(net754),
    .GATE(net695),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2095_ (.D(net802),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2096_ (.D(net780),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2097_ (.D(net759),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2098_ (.D(net753),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2099_ (.D(net750),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2100_ (.D(net748),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2101_ (.D(net746),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2102_ (.D(net744),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2103_ (.D(net743),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2104_ (.D(net740),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2105_ (.D(net801),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2106_ (.D(net799),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2107_ (.D(net797),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2108_ (.D(net795),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2109_ (.D(net793),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2110_ (.D(net791),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2111_ (.D(net789),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2112_ (.D(net786),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2113_ (.D(net36),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2114_ (.D(net783),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2115_ (.D(net779),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2116_ (.D(net777),
    .GATE(net738),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2117_ (.D(net774),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2118_ (.D(net772),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2119_ (.D(net771),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2120_ (.D(net768),
    .GATE(net736),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2121_ (.D(net43),
    .GATE(net739),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2122_ (.D(net764),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2123_ (.D(net762),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2124_ (.D(net760),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2125_ (.D(net756),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _2126_ (.D(net755),
    .GATE(net737),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__dfxtp_1 _2127_ (.CLK(clknet_1_1__leaf_UserCLK_regs),
    .D(_0000_),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2128_ (.CLK(clknet_1_0__leaf_UserCLK_regs),
    .D(_0001_),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2129_ (.CLK(clknet_1_0__leaf_UserCLK_regs),
    .D(_0002_),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2130_ (.CLK(clknet_1_0__leaf_UserCLK_regs),
    .D(_0003_),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2131_ (.CLK(clknet_1_0__leaf_UserCLK_regs),
    .D(_0004_),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2132_ (.CLK(clknet_1_1__leaf_UserCLK_regs),
    .D(_0005_),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2133_ (.CLK(clknet_1_1__leaf_UserCLK_regs),
    .D(_0006_),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__dfxtp_1 _2134_ (.CLK(clknet_1_1__leaf_UserCLK_regs),
    .D(_0007_),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__buf_1 _2135_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG0 ),
    .X(net142));
 sky130_fd_sc_hd__buf_4 _2136_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG1 ),
    .X(net143));
 sky130_fd_sc_hd__buf_8 clone18 (.A(net428),
    .X(net412));
 sky130_fd_sc_hd__buf_6 rebuffer81 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_6 _2139_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .X(net146));
 sky130_fd_sc_hd__buf_6 _2140_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .X(net147));
 sky130_fd_sc_hd__buf_4 _2141_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .X(net148));
 sky130_fd_sc_hd__buf_1 _2142_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .X(net149));
 sky130_fd_sc_hd__buf_8 _2143_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .X(net150));
 sky130_fd_sc_hd__buf_4 _2144_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .X(net151));
 sky130_fd_sc_hd__buf_4 _2145_ (.A(net413),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_2 _2147_ (.A(net14),
    .X(net154));
 sky130_fd_sc_hd__buf_1 _2148_ (.A(net15),
    .X(net155));
 sky130_fd_sc_hd__buf_1 _2149_ (.A(net16),
    .X(net156));
 sky130_fd_sc_hd__buf_1 _2150_ (.A(net17),
    .X(net157));
 sky130_fd_sc_hd__buf_1 _2151_ (.A(net18),
    .X(net158));
 sky130_fd_sc_hd__buf_1 _2152_ (.A(net19),
    .X(net159));
 sky130_fd_sc_hd__buf_1 _2153_ (.A(net20),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _2154_ (.A(net21),
    .X(net161));
 sky130_fd_sc_hd__buf_1 _2155_ (.A(E6END[2]),
    .X(net162));
 sky130_fd_sc_hd__buf_1 _2156_ (.A(E6END[3]),
    .X(net165));
 sky130_fd_sc_hd__buf_1 _2157_ (.A(E6END[4]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 _2158_ (.A(E6END[5]),
    .X(net167));
 sky130_fd_sc_hd__buf_1 _2159_ (.A(E6END[6]),
    .X(net168));
 sky130_fd_sc_hd__buf_1 _2160_ (.A(E6END[7]),
    .X(net169));
 sky130_fd_sc_hd__buf_1 _2161_ (.A(E6END[8]),
    .X(net170));
 sky130_fd_sc_hd__buf_1 _2162_ (.A(E6END[9]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 _2163_ (.A(E6END[10]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 _2164_ (.A(E6END[11]),
    .X(net173));
 sky130_fd_sc_hd__buf_6 rebuffer131 (.A(_0046_),
    .X(net525));
 sky130_fd_sc_hd__buf_6 rebuffer80 (.A(_0027_),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_1 _2167_ (.A(EE4END[4]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 _2168_ (.A(EE4END[5]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 _2169_ (.A(EE4END[6]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 _2170_ (.A(EE4END[7]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 _2171_ (.A(EE4END[8]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 _2172_ (.A(EE4END[9]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 _2173_ (.A(EE4END[10]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 _2174_ (.A(EE4END[11]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 _2175_ (.A(EE4END[12]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 _2176_ (.A(EE4END[13]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 _2177_ (.A(EE4END[14]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 _2178_ (.A(EE4END[15]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 _2179_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG0 ),
    .X(net177));
 sky130_fd_sc_hd__fill_1 FILLER_0_41 ();
 sky130_fd_sc_hd__clkbuf_2 _2181_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer118 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 _2183_ (.A(net803),
    .X(net190));
 sky130_fd_sc_hd__buf_1 _2184_ (.A(net781),
    .X(net201));
 sky130_fd_sc_hd__buf_1 _2185_ (.A(net758),
    .X(net212));
 sky130_fd_sc_hd__buf_1 _2186_ (.A(net753),
    .X(net215));
 sky130_fd_sc_hd__buf_1 _2187_ (.A(net751),
    .X(net216));
 sky130_fd_sc_hd__buf_1 _2188_ (.A(net749),
    .X(net217));
 sky130_fd_sc_hd__buf_1 _2189_ (.A(net747),
    .X(net218));
 sky130_fd_sc_hd__buf_1 _2190_ (.A(net745),
    .X(net219));
 sky130_fd_sc_hd__buf_1 _2191_ (.A(net743),
    .X(net220));
 sky130_fd_sc_hd__buf_1 _2192_ (.A(net740),
    .X(net221));
 sky130_fd_sc_hd__buf_1 _2193_ (.A(net800),
    .X(net191));
 sky130_fd_sc_hd__buf_1 _2194_ (.A(net798),
    .X(net192));
 sky130_fd_sc_hd__buf_1 _2195_ (.A(net796),
    .X(net193));
 sky130_fd_sc_hd__buf_1 _2196_ (.A(net794),
    .X(net194));
 sky130_fd_sc_hd__buf_1 _2197_ (.A(net792),
    .X(net195));
 sky130_fd_sc_hd__buf_1 _2198_ (.A(net790),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 _2199_ (.A(net788),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 _2200_ (.A(net787),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 _2201_ (.A(net784),
    .X(net199));
 sky130_fd_sc_hd__buf_1 _2202_ (.A(net782),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 _2203_ (.A(net778),
    .X(net202));
 sky130_fd_sc_hd__buf_1 _2204_ (.A(net776),
    .X(net203));
 sky130_fd_sc_hd__buf_1 _2205_ (.A(net775),
    .X(net204));
 sky130_fd_sc_hd__buf_1 _2206_ (.A(net773),
    .X(net205));
 sky130_fd_sc_hd__buf_1 _2207_ (.A(net770),
    .X(net206));
 sky130_fd_sc_hd__buf_1 _2208_ (.A(net769),
    .X(net207));
 sky130_fd_sc_hd__buf_1 _2209_ (.A(net766),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 _2210_ (.A(net764),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 _2211_ (.A(net45),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 _2212_ (.A(net760),
    .X(net211));
 sky130_fd_sc_hd__buf_1 _2213_ (.A(net757),
    .X(net213));
 sky130_fd_sc_hd__buf_1 _2214_ (.A(net755),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 _2215_ (.A(net739),
    .X(net222));
 sky130_fd_sc_hd__buf_1 _2216_ (.A(net699),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 _2217_ (.A(FrameStrobe[2]),
    .X(net234));
 sky130_fd_sc_hd__buf_1 _2218_ (.A(net690),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 _2219_ (.A(net686),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 _2220_ (.A(net682),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 _2221_ (.A(net676),
    .X(net238));
 sky130_fd_sc_hd__buf_1 _2222_ (.A(net672),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 _2223_ (.A(net665),
    .X(net240));
 sky130_fd_sc_hd__buf_1 _2224_ (.A(net664),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 _2225_ (.A(net734),
    .X(net223));
 sky130_fd_sc_hd__buf_2 _2226_ (.A(net731),
    .X(net224));
 sky130_fd_sc_hd__buf_1 _2227_ (.A(FrameStrobe[12]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 _2228_ (.A(FrameStrobe[13]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 _2229_ (.A(net719),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 _2230_ (.A(net714),
    .X(net228));
 sky130_fd_sc_hd__buf_1 _2231_ (.A(net711),
    .X(net229));
 sky130_fd_sc_hd__buf_1 _2232_ (.A(net707),
    .X(net230));
 sky130_fd_sc_hd__buf_1 _2233_ (.A(net702),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 _2234_ (.A(net56),
    .X(net232));
 sky130_fd_sc_hd__buf_6 _2235_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .X(net242));
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__clkbuf_2 _2237_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG2 ),
    .X(net244));
 sky130_fd_sc_hd__buf_6 _2238_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .X(net245));
 sky130_fd_sc_hd__buf_4 _2239_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .X(net246));
 sky130_fd_sc_hd__buf_2 _2240_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .X(net247));
 sky130_fd_sc_hd__buf_6 _2241_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .X(net248));
 sky130_fd_sc_hd__buf_1 _2242_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .X(net249));
 sky130_fd_sc_hd__decap_3 FILLER_0_141 ();
 sky130_fd_sc_hd__clkbuf_2 _2244_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .X(net251));
 sky130_fd_sc_hd__buf_1 _2245_ (.A(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_2 _2247_ (.A(net71),
    .X(net254));
 sky130_fd_sc_hd__buf_4 _2248_ (.A(net72),
    .X(net255));
 sky130_fd_sc_hd__buf_1 _2249_ (.A(net73),
    .X(net256));
 sky130_fd_sc_hd__buf_2 _2250_ (.A(net74),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 _2251_ (.A(net75),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 _2252_ (.A(net76),
    .X(net259));
 sky130_fd_sc_hd__buf_1 _2253_ (.A(net77),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_2 _2254_ (.A(net78),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 _2255_ (.A(N4END[4]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 _2256_ (.A(N4END[5]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 _2257_ (.A(N4END[6]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 _2258_ (.A(N4END[7]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 _2259_ (.A(N4END[8]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 _2260_ (.A(N4END[9]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 _2261_ (.A(N4END[10]),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 _2262_ (.A(N4END[11]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 _2263_ (.A(N4END[12]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 _2264_ (.A(N4END[13]),
    .X(net277));
 sky130_fd_sc_hd__buf_1 _2265_ (.A(N4END[14]),
    .X(net263));
 sky130_fd_sc_hd__buf_1 _2266_ (.A(N4END[15]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 _2267_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG0 ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net543));
 sky130_fd_sc_hd__buf_6 _2270_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 _2271_ (.A(NN4END[4]),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 _2272_ (.A(NN4END[5]),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 _2273_ (.A(NN4END[6]),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 _2274_ (.A(NN4END[7]),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 _2275_ (.A(NN4END[8]),
    .X(net288));
 sky130_fd_sc_hd__buf_1 _2276_ (.A(NN4END[9]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 _2277_ (.A(NN4END[10]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 _2278_ (.A(NN4END[11]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 _2279_ (.A(NN4END[12]),
    .X(net292));
 sky130_fd_sc_hd__buf_1 _2280_ (.A(NN4END[13]),
    .X(net293));
 sky130_fd_sc_hd__buf_1 _2281_ (.A(NN4END[14]),
    .X(net279));
 sky130_fd_sc_hd__buf_1 _2282_ (.A(NN4END[15]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 _2283_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG0 ),
    .X(net281));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__buf_4 _2285_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .X(net283));
 sky130_fd_sc_hd__fill_2 FILLER_0_265 ();
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_2 rebuffer35 (.A(net435),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_2 rebuffer82 (.A(net487),
    .X(net476));
 sky130_fd_sc_hd__buf_6 _2291_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 _2292_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .X(net299));
 sky130_fd_sc_hd__buf_6 _2293_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 _2294_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .X(net301));
 sky130_fd_sc_hd__buf_6 _2295_ (.A(net526),
    .X(net302));
 sky130_fd_sc_hd__buf_2 _2296_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .X(net303));
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__buf_6 _2298_ (.A(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .X(net305));
 sky130_fd_sc_hd__buf_1 _2299_ (.A(net99),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 _2300_ (.A(net100),
    .X(net307));
 sky130_fd_sc_hd__buf_1 _2301_ (.A(net101),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 _2302_ (.A(net102),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 _2303_ (.A(net103),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 _2304_ (.A(net104),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_2 _2305_ (.A(net105),
    .X(net312));
 sky130_fd_sc_hd__buf_1 _2306_ (.A(net106),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 _2307_ (.A(S4END[4]),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_2 _2308_ (.A(S4END[5]),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 _2309_ (.A(S4END[6]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 _2310_ (.A(S4END[7]),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 _2311_ (.A(S4END[8]),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 _2312_ (.A(S4END[9]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 _2313_ (.A(S4END[10]),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 _2314_ (.A(S4END[11]),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 _2315_ (.A(S4END[12]),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_2 _2316_ (.A(S4END[13]),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 _2317_ (.A(S4END[14]),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_2 _2318_ (.A(S4END[15]),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 _2319_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG0 ),
    .X(net317));
 sky130_fd_sc_hd__buf_1 _2320_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG1 ),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 _2321_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG2 ),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 _2322_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG3 ),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 _2323_ (.A(SS4END[4]),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 _2324_ (.A(SS4END[5]),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 _2325_ (.A(SS4END[6]),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 _2326_ (.A(SS4END[7]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_2 _2327_ (.A(SS4END[8]),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 _2328_ (.A(SS4END[9]),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_2 _2329_ (.A(SS4END[10]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 _2330_ (.A(SS4END[11]),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 _2331_ (.A(SS4END[12]),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 _2332_ (.A(SS4END[13]),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_2 _2333_ (.A(SS4END[14]),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_2 _2334_ (.A(SS4END[15]),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_1 _2335_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG0 ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net548));
 sky130_fd_sc_hd__buf_1 _2337_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG2 ),
    .X(net335));
 sky130_fd_sc_hd__buf_1 _2338_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG3 ),
    .X(net336));
 sky130_fd_sc_hd__buf_2 _2339_ (.A(clknet_1_0__leaf_UserCLK),
    .X(net346));
 sky130_fd_sc_hd__buf_1 _2340_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG0 ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer132 (.A(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .X(net526));
 sky130_fd_sc_hd__buf_6 clone17 (.A(G),
    .X(net411));
 sky130_fd_sc_hd__buf_6 _2343_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG3 ),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_1 _2344_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .X(net351));
 sky130_fd_sc_hd__buf_6 _2345_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .X(net352));
 sky130_fd_sc_hd__buf_1 _2346_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .X(net353));
 sky130_fd_sc_hd__buf_6 _2347_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .X(net354));
 sky130_fd_sc_hd__buf_6 _2348_ (.A(net479),
    .X(net355));
 sky130_fd_sc_hd__buf_1 _2349_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .X(net356));
 sky130_fd_sc_hd__buf_6 _2350_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .X(net357));
 sky130_fd_sc_hd__buf_1 _2351_ (.A(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .X(net358));
 sky130_fd_sc_hd__buf_1 _2352_ (.A(net127),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_2 _2353_ (.A(net128),
    .X(net360));
 sky130_fd_sc_hd__buf_2 _2354_ (.A(net129),
    .X(net361));
 sky130_fd_sc_hd__buf_1 _2355_ (.A(net130),
    .X(net362));
 sky130_fd_sc_hd__buf_1 _2356_ (.A(net131),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 _2357_ (.A(net132),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 _2358_ (.A(net133),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 _2359_ (.A(net134),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_2 _2360_ (.A(W6END[2]),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_2 _2361_ (.A(W6END[3]),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 _2362_ (.A(W6END[4]),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 _2363_ (.A(W6END[5]),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 _2364_ (.A(W6END[6]),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 _2365_ (.A(W6END[7]),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 _2366_ (.A(W6END[8]),
    .X(net375));
 sky130_fd_sc_hd__buf_4 _2367_ (.A(W6END[9]),
    .X(net376));
 sky130_fd_sc_hd__buf_4 _2368_ (.A(W6END[10]),
    .X(net377));
 sky130_fd_sc_hd__buf_4 _2369_ (.A(W6END[11]),
    .X(net378));
 sky130_fd_sc_hd__decap_3 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__clkbuf_2 _2372_ (.A(WW4END[4]),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_2 _2373_ (.A(WW4END[5]),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 _2374_ (.A(WW4END[6]),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_2 _2375_ (.A(WW4END[7]),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 _2376_ (.A(WW4END[8]),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 _2377_ (.A(WW4END[9]),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_2 _2378_ (.A(WW4END[10]),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_2 _2379_ (.A(WW4END[11]),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_2 _2380_ (.A(WW4END[12]),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_2 _2381_ (.A(WW4END[13]),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_2 _2382_ (.A(WW4END[14]),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_2 _2383_ (.A(WW4END[15]),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .X(net544));
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__buf_1 _2386_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG2 ),
    .X(net384));
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_679 ();
 sky130_fd_sc_hd__buf_8 fanout617 (.A(net431),
    .X(net617));
 sky130_fd_sc_hd__buf_12 fanout618 (.A(net480),
    .X(net618));
 sky130_fd_sc_hd__buf_6 fanout619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__buf_8 fanout620 (.A(net432),
    .X(net620));
 sky130_fd_sc_hd__buf_4 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_4 fanout622 (.A(H),
    .X(net622));
 sky130_fd_sc_hd__buf_8 fanout623 (.A(net624),
    .X(net623));
 sky130_fd_sc_hd__buf_8 fanout624 (.A(C),
    .X(net624));
 sky130_fd_sc_hd__buf_2 fanout625 (.A(net627),
    .X(net625));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__buf_8 fanout627 (.A(C),
    .X(net627));
 sky130_fd_sc_hd__buf_6 fanout628 (.A(net629),
    .X(net628));
 sky130_fd_sc_hd__buf_8 fanout629 (.A(G),
    .X(net629));
 sky130_fd_sc_hd__buf_2 fanout630 (.A(net632),
    .X(net630));
 sky130_fd_sc_hd__buf_6 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__buf_6 fanout632 (.A(G),
    .X(net632));
 sky130_fd_sc_hd__buf_8 fanout633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__buf_8 fanout634 (.A(net637),
    .X(net634));
 sky130_fd_sc_hd__buf_8 fanout635 (.A(net636),
    .X(net635));
 sky130_fd_sc_hd__buf_8 fanout636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__buf_8 fanout637 (.A(F),
    .X(net637));
 sky130_fd_sc_hd__buf_8 fanout638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__buf_8 fanout639 (.A(D),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_2 fanout640 (.A(net641),
    .X(net640));
 sky130_fd_sc_hd__buf_2 fanout641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_2 fanout642 (.A(D),
    .X(net642));
 sky130_fd_sc_hd__buf_2 fanout643 (.A(net645),
    .X(net643));
 sky130_fd_sc_hd__buf_8 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_8 fanout645 (.A(E),
    .X(net645));
 sky130_fd_sc_hd__buf_2 fanout646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__buf_2 fanout647 (.A(E),
    .X(net647));
 sky130_fd_sc_hd__buf_8 fanout648 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__buf_8 fanout649 (.A(net652),
    .X(net649));
 sky130_fd_sc_hd__buf_2 fanout650 (.A(net651),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 fanout651 (.A(net652),
    .X(net651));
 sky130_fd_sc_hd__buf_8 fanout652 (.A(B),
    .X(net652));
 sky130_fd_sc_hd__buf_8 fanout653 (.A(net657),
    .X(net653));
 sky130_fd_sc_hd__buf_2 fanout654 (.A(net656),
    .X(net654));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout655 (.A(net656),
    .X(net655));
 sky130_fd_sc_hd__buf_2 fanout656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__buf_12 fanout657 (.A(A),
    .X(net657));
 sky130_fd_sc_hd__buf_4 fanout658 (.A(_0247_),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_4 fanout659 (.A(net118),
    .X(net659));
 sky130_fd_sc_hd__buf_4 fanout660 (.A(net117),
    .X(net660));
 sky130_fd_sc_hd__buf_2 fanout661 (.A(net58),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_2 fanout662 (.A(net664),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_1 fanout663 (.A(net664),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_2 fanout664 (.A(net58),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_2 fanout665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_2 fanout666 (.A(net667),
    .X(net666));
 sky130_fd_sc_hd__buf_2 fanout667 (.A(FrameStrobe[8]),
    .X(net667));
 sky130_fd_sc_hd__buf_2 fanout668 (.A(FrameStrobe[8]),
    .X(net668));
 sky130_fd_sc_hd__buf_2 fanout669 (.A(net671),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_2 fanout670 (.A(net671),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_2 fanout671 (.A(net673),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_2 fanout672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_2 fanout673 (.A(FrameStrobe[7]),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_2 fanout674 (.A(net677),
    .X(net674));
 sky130_fd_sc_hd__clkbuf_2 fanout675 (.A(net677),
    .X(net675));
 sky130_fd_sc_hd__buf_1 fanout676 (.A(net677),
    .X(net676));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_2 fanout678 (.A(FrameStrobe[6]),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_2 fanout679 (.A(net681),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_2 fanout680 (.A(net681),
    .X(net680));
 sky130_fd_sc_hd__buf_2 fanout681 (.A(net57),
    .X(net681));
 sky130_fd_sc_hd__buf_2 fanout682 (.A(net57),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_2 fanout683 (.A(net686),
    .X(net683));
 sky130_fd_sc_hd__buf_2 fanout684 (.A(net686),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_2 fanout685 (.A(net686),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_2 fanout686 (.A(FrameStrobe[4]),
    .X(net686));
 sky130_fd_sc_hd__buf_2 fanout687 (.A(FrameStrobe[3]),
    .X(net687));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout688 (.A(FrameStrobe[3]),
    .X(net688));
 sky130_fd_sc_hd__buf_2 fanout689 (.A(FrameStrobe[3]),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_2 fanout690 (.A(FrameStrobe[3]),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_2 fanout691 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__buf_2 fanout692 (.A(FrameStrobe[2]),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_2 fanout693 (.A(net694),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_2 fanout694 (.A(FrameStrobe[2]),
    .X(net694));
 sky130_fd_sc_hd__buf_2 fanout695 (.A(net697),
    .X(net695));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout696 (.A(net697),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_2 fanout697 (.A(net699),
    .X(net697));
 sky130_fd_sc_hd__buf_2 fanout698 (.A(net699),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_2 fanout699 (.A(FrameStrobe[1]),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_2 fanout700 (.A(net703),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_2 fanout701 (.A(net703),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_2 fanout702 (.A(net703),
    .X(net702));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout703 (.A(FrameStrobe[18]),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_2 fanout704 (.A(FrameStrobe[17]),
    .X(net704));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout705 (.A(FrameStrobe[17]),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_2 fanout706 (.A(FrameStrobe[17]),
    .X(net706));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout707 (.A(FrameStrobe[17]),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_2 fanout708 (.A(net709),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_2 fanout709 (.A(FrameStrobe[16]),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_2 fanout710 (.A(FrameStrobe[16]),
    .X(net710));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout711 (.A(FrameStrobe[16]),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_2 fanout712 (.A(net55),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_2 fanout713 (.A(net714),
    .X(net713));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout714 (.A(net715),
    .X(net714));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout715 (.A(net55),
    .X(net715));
 sky130_fd_sc_hd__buf_2 fanout716 (.A(FrameStrobe[14]),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_2 fanout717 (.A(FrameStrobe[14]),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_2 fanout718 (.A(FrameStrobe[14]),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_2 fanout719 (.A(FrameStrobe[14]),
    .X(net719));
 sky130_fd_sc_hd__buf_2 fanout720 (.A(net721),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_2 fanout721 (.A(FrameStrobe[13]),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_2 fanout722 (.A(FrameStrobe[13]),
    .X(net722));
 sky130_fd_sc_hd__buf_1 fanout723 (.A(FrameStrobe[13]),
    .X(net723));
 sky130_fd_sc_hd__buf_2 fanout724 (.A(net726),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_2 fanout725 (.A(net726),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_2 fanout726 (.A(FrameStrobe[12]),
    .X(net726));
 sky130_fd_sc_hd__buf_2 fanout727 (.A(FrameStrobe[12]),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_2 fanout728 (.A(net729),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_4 fanout729 (.A(net730),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_2 fanout730 (.A(net731),
    .X(net730));
 sky130_fd_sc_hd__buf_2 fanout731 (.A(FrameStrobe[11]),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_2 fanout732 (.A(net733),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_2 fanout733 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_2 fanout734 (.A(net735),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_2 fanout735 (.A(FrameStrobe[10]),
    .X(net735));
 sky130_fd_sc_hd__buf_2 fanout736 (.A(net738),
    .X(net736));
 sky130_fd_sc_hd__buf_2 fanout737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_2 fanout738 (.A(net739),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_2 fanout739 (.A(FrameStrobe[0]),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_4 fanout740 (.A(net741),
    .X(net740));
 sky130_fd_sc_hd__buf_4 fanout741 (.A(net54),
    .X(net741));
 sky130_fd_sc_hd__buf_4 fanout742 (.A(FrameData[8]),
    .X(net742));
 sky130_fd_sc_hd__buf_4 fanout743 (.A(FrameData[8]),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_4 fanout744 (.A(net745),
    .X(net744));
 sky130_fd_sc_hd__buf_4 fanout745 (.A(net53),
    .X(net745));
 sky130_fd_sc_hd__buf_4 fanout746 (.A(FrameData[6]),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_4 fanout747 (.A(FrameData[6]),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_4 fanout748 (.A(net749),
    .X(net748));
 sky130_fd_sc_hd__buf_4 fanout749 (.A(net52),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_4 fanout750 (.A(net751),
    .X(net750));
 sky130_fd_sc_hd__buf_4 fanout751 (.A(net51),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_4 fanout752 (.A(net753),
    .X(net752));
 sky130_fd_sc_hd__buf_4 fanout753 (.A(net50),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_4 fanout754 (.A(net755),
    .X(net754));
 sky130_fd_sc_hd__buf_4 fanout755 (.A(net49),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 fanout756 (.A(net757),
    .X(net756));
 sky130_fd_sc_hd__buf_4 fanout757 (.A(net48),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_4 fanout758 (.A(net759),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_4 fanout759 (.A(net47),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_4 fanout760 (.A(net761),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_8 fanout761 (.A(net46),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_4 fanout762 (.A(net763),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_8 fanout763 (.A(net45),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_4 fanout764 (.A(net765),
    .X(net764));
 sky130_fd_sc_hd__buf_4 fanout765 (.A(net44),
    .X(net765));
 sky130_fd_sc_hd__buf_4 fanout766 (.A(net767),
    .X(net766));
 sky130_fd_sc_hd__buf_4 fanout767 (.A(net43),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_4 fanout768 (.A(net769),
    .X(net768));
 sky130_fd_sc_hd__buf_4 fanout769 (.A(net42),
    .X(net769));
 sky130_fd_sc_hd__buf_4 fanout770 (.A(net41),
    .X(net770));
 sky130_fd_sc_hd__buf_4 fanout771 (.A(net41),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_4 fanout772 (.A(FrameData[23]),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_4 fanout773 (.A(FrameData[23]),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_4 fanout774 (.A(FrameData[22]),
    .X(net774));
 sky130_fd_sc_hd__buf_4 fanout775 (.A(FrameData[22]),
    .X(net775));
 sky130_fd_sc_hd__buf_4 fanout776 (.A(net777),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_4 fanout777 (.A(net40),
    .X(net777));
 sky130_fd_sc_hd__buf_4 fanout778 (.A(net779),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_4 fanout779 (.A(net39),
    .X(net779));
 sky130_fd_sc_hd__buf_2 fanout780 (.A(net781),
    .X(net780));
 sky130_fd_sc_hd__buf_4 fanout781 (.A(net38),
    .X(net781));
 sky130_fd_sc_hd__buf_4 fanout782 (.A(net783),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_4 fanout783 (.A(net37),
    .X(net783));
 sky130_fd_sc_hd__buf_4 fanout784 (.A(net785),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_4 fanout785 (.A(net36),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_4 fanout786 (.A(FrameData[17]),
    .X(net786));
 sky130_fd_sc_hd__buf_4 fanout787 (.A(FrameData[17]),
    .X(net787));
 sky130_fd_sc_hd__buf_4 fanout788 (.A(net789),
    .X(net788));
 sky130_fd_sc_hd__buf_4 fanout789 (.A(net35),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_4 fanout790 (.A(net791),
    .X(net790));
 sky130_fd_sc_hd__buf_4 fanout791 (.A(net34),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_4 fanout792 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__buf_4 fanout793 (.A(net33),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_4 fanout794 (.A(net795),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_4 fanout795 (.A(net32),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_4 fanout796 (.A(net797),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_4 fanout797 (.A(net31),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_4 fanout798 (.A(net799),
    .X(net798));
 sky130_fd_sc_hd__buf_4 fanout799 (.A(net30),
    .X(net799));
 sky130_fd_sc_hd__buf_4 fanout800 (.A(net801),
    .X(net800));
 sky130_fd_sc_hd__buf_4 fanout801 (.A(net29),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_4 fanout802 (.A(net803),
    .X(net802));
 sky130_fd_sc_hd__buf_4 fanout803 (.A(net28),
    .X(net803));
 sky130_fd_sc_hd__buf_2 fanout804 (.A(net23),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_4 fanout805 (.A(net22),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_4 fanout806 (.A(net5),
    .X(net806));
 sky130_fd_sc_hd__buf_4 fanout807 (.A(net4),
    .X(net807));
 sky130_fd_sc_hd__buf_12 input1 (.A(Ci),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(E1END[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(E1END[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(E1END[2]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(E1END[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(E2END[0]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(E2END[1]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(E2END[2]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(E2END[3]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(E2END[4]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(E2END[5]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(E2END[6]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(E2END[7]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(E2MID[0]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(E2MID[1]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(E2MID[2]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(E2MID[3]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(E2MID[4]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(E2MID[5]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(E2MID[6]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(E2MID[7]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(E6END[0]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(E6END[1]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(EE4END[0]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(EE4END[1]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(EE4END[2]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(EE4END[3]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(FrameData[0]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(FrameData[10]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(FrameData[11]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(FrameData[12]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(FrameData[13]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(FrameData[14]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(FrameData[15]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(FrameData[16]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(FrameData[18]),
    .X(net36));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(FrameData[19]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(FrameData[1]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(FrameData[20]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(FrameData[21]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(FrameData[24]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(FrameData[25]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(FrameData[26]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(FrameData[27]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(FrameData[28]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(FrameData[29]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(FrameData[2]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(FrameData[30]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input49 (.A(FrameData[31]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(FrameData[3]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(FrameData[4]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(FrameData[5]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(FrameData[7]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(FrameData[9]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(FrameStrobe[15]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(FrameStrobe[19]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(FrameStrobe[5]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(FrameStrobe[9]),
    .X(net58));
 sky130_fd_sc_hd__buf_4 input59 (.A(N1END[0]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(N1END[1]),
    .X(net60));
 sky130_fd_sc_hd__buf_4 input61 (.A(N1END[2]),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input62 (.A(N1END[3]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(N2END[0]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(N2END[1]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(N2END[2]),
    .X(net65));
 sky130_fd_sc_hd__buf_2 input66 (.A(N2END[3]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(N2END[4]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(N2END[5]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input69 (.A(N2END[6]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input70 (.A(N2END[7]),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 input71 (.A(N2MID[0]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(N2MID[1]),
    .X(net72));
 sky130_fd_sc_hd__buf_2 input73 (.A(N2MID[2]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(N2MID[3]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(N2MID[4]),
    .X(net75));
 sky130_fd_sc_hd__buf_2 input76 (.A(N2MID[5]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(N2MID[6]),
    .X(net77));
 sky130_fd_sc_hd__buf_2 input78 (.A(N2MID[7]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(N4END[0]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(N4END[1]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(N4END[2]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(N4END[3]),
    .X(net82));
 sky130_fd_sc_hd__dlymetal6s2s_1 input83 (.A(NN4END[0]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(NN4END[1]),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 input85 (.A(NN4END[2]),
    .X(net85));
 sky130_fd_sc_hd__dlymetal6s2s_1 input86 (.A(NN4END[3]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(S1END[0]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(S1END[1]),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(S1END[2]),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input90 (.A(S1END[3]),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(S2END[0]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 input92 (.A(S2END[1]),
    .X(net92));
 sky130_fd_sc_hd__buf_2 input93 (.A(S2END[2]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(S2END[3]),
    .X(net94));
 sky130_fd_sc_hd__buf_2 input95 (.A(S2END[4]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(S2END[5]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(S2END[6]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(S2END[7]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(S2MID[0]),
    .X(net99));
 sky130_fd_sc_hd__buf_2 input100 (.A(S2MID[1]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(S2MID[2]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(S2MID[3]),
    .X(net102));
 sky130_fd_sc_hd__dlymetal6s2s_1 input103 (.A(S2MID[4]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(S2MID[5]),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 input105 (.A(S2MID[6]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(S2MID[7]),
    .X(net106));
 sky130_fd_sc_hd__buf_2 input107 (.A(S4END[0]),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(S4END[1]),
    .X(net108));
 sky130_fd_sc_hd__buf_2 input109 (.A(S4END[2]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(S4END[3]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(SS4END[0]),
    .X(net111));
 sky130_fd_sc_hd__buf_2 input112 (.A(SS4END[1]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(SS4END[2]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(SS4END[3]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(W1END[0]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 input116 (.A(W1END[1]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(W1END[2]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(W1END[3]),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 input119 (.A(W2END[0]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input120 (.A(W2END[1]),
    .X(net120));
 sky130_fd_sc_hd__buf_2 input121 (.A(W2END[2]),
    .X(net121));
 sky130_fd_sc_hd__buf_2 input122 (.A(W2END[3]),
    .X(net122));
 sky130_fd_sc_hd__buf_2 input123 (.A(W2END[4]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(W2END[5]),
    .X(net124));
 sky130_fd_sc_hd__dlymetal6s2s_1 input125 (.A(W2END[6]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(W2END[7]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(W2MID[0]),
    .X(net127));
 sky130_fd_sc_hd__dlymetal6s2s_1 input128 (.A(W2MID[1]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(W2MID[2]),
    .X(net129));
 sky130_fd_sc_hd__dlymetal6s2s_1 input130 (.A(W2MID[3]),
    .X(net130));
 sky130_fd_sc_hd__buf_2 input131 (.A(W2MID[4]),
    .X(net131));
 sky130_fd_sc_hd__dlymetal6s2s_1 input132 (.A(W2MID[5]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(W2MID[6]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input134 (.A(W2MID[7]),
    .X(net134));
 sky130_fd_sc_hd__buf_2 input135 (.A(W6END[0]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 input136 (.A(W6END[1]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(WW4END[0]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 input138 (.A(WW4END[1]),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(WW4END[2]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input140 (.A(WW4END[3]),
    .X(net140));
 sky130_fd_sc_hd__buf_8 output141 (.A(net141),
    .X(Co));
 sky130_fd_sc_hd__clkbuf_4 output142 (.A(net142),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__buf_4 output143 (.A(net143),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__buf_8 output144 (.A(\Inst_LUT4AB_switch_matrix.E1BEG2 ),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__buf_4 output145 (.A(\Inst_LUT4AB_switch_matrix.E1BEG3 ),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__buf_8 output146 (.A(net146),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__buf_4 output147 (.A(net147),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__buf_6 output148 (.A(net148),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__buf_8 output150 (.A(net150),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__buf_6 output151 (.A(net151),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__buf_6 output152 (.A(net152),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__buf_6 output153 (.A(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__buf_6 output163 (.A(\Inst_LUT4AB_switch_matrix.E6BEG0 ),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__buf_8 output164 (.A(\Inst_LUT4AB_switch_matrix.E6BEG1 ),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__buf_6 output178 (.A(\Inst_LUT4AB_switch_matrix.EE4BEG1 ),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__buf_6 output179 (.A(net179),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__buf_8 output180 (.A(\Inst_LUT4AB_switch_matrix.EE4BEG3 ),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net226),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net232),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net241),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_4 output242 (.A(net242),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__buf_4 output243 (.A(\Inst_LUT4AB_switch_matrix.N1BEG1 ),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__buf_4 output244 (.A(net244),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_8 output245 (.A(net245),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_4 output246 (.A(net246),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_6 output247 (.A(net247),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_8 output248 (.A(net248),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_6 output249 (.A(net249),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_8 output250 (.A(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_6 output251 (.A(net251),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_4 output252 (.A(net252),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_6 output253 (.A(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_4 output265 (.A(net265),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_6 output266 (.A(\Inst_LUT4AB_switch_matrix.N4BEG1 ),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_6 output267 (.A(\Inst_LUT4AB_switch_matrix.N4BEG2 ),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_8 output268 (.A(net268),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__buf_6 output282 (.A(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_8 output283 (.A(net283),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_8 output284 (.A(\Inst_LUT4AB_switch_matrix.NN4BEG3 ),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_8 output294 (.A(\Inst_LUT4AB_switch_matrix.S1BEG0 ),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_4 output295 (.A(\Inst_LUT4AB_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__buf_8 output296 (.A(\Inst_LUT4AB_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_8 output297 (.A(\Inst_LUT4AB_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_8 output298 (.A(net298),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_6 output299 (.A(net299),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_8 output300 (.A(net300),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_6 output301 (.A(net301),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_8 output302 (.A(net302),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__buf_6 output303 (.A(net303),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__buf_6 output304 (.A(net443),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__buf_6 output305 (.A(net305),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__buf_6 output317 (.A(net317),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__buf_4 output319 (.A(net319),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__buf_2 output333 (.A(net333),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__buf_6 output334 (.A(\Inst_LUT4AB_switch_matrix.SS4BEG1 ),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__buf_4 output335 (.A(net335),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__buf_4 output336 (.A(net336),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__buf_2 output344 (.A(net344),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net345),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__buf_1 output346 (.A(net346),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_4 output347 (.A(net347),
    .X(W1BEG[0]));
 sky130_fd_sc_hd__buf_4 output348 (.A(\Inst_LUT4AB_switch_matrix.W1BEG1 ),
    .X(W1BEG[1]));
 sky130_fd_sc_hd__buf_8 output349 (.A(\Inst_LUT4AB_switch_matrix.W1BEG2 ),
    .X(W1BEG[2]));
 sky130_fd_sc_hd__buf_8 output350 (.A(net350),
    .X(W1BEG[3]));
 sky130_fd_sc_hd__buf_4 output351 (.A(net351),
    .X(W2BEG[0]));
 sky130_fd_sc_hd__buf_8 output352 (.A(net352),
    .X(W2BEG[1]));
 sky130_fd_sc_hd__buf_4 output353 (.A(net353),
    .X(W2BEG[2]));
 sky130_fd_sc_hd__buf_8 output354 (.A(net354),
    .X(W2BEG[3]));
 sky130_fd_sc_hd__buf_8 output355 (.A(net355),
    .X(W2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output356 (.A(net356),
    .X(W2BEG[5]));
 sky130_fd_sc_hd__buf_8 output357 (.A(net357),
    .X(W2BEG[6]));
 sky130_fd_sc_hd__buf_6 output358 (.A(net358),
    .X(W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(W2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .X(W2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .X(W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output366 (.A(net366),
    .X(W2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output367 (.A(net367),
    .X(W6BEG[0]));
 sky130_fd_sc_hd__buf_6 output368 (.A(\Inst_LUT4AB_switch_matrix.W6BEG0 ),
    .X(W6BEG[10]));
 sky130_fd_sc_hd__buf_6 output369 (.A(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .X(W6BEG[11]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .X(W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(W6BEG[2]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .X(W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .X(W6BEG[5]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net375),
    .X(W6BEG[6]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .X(W6BEG[7]));
 sky130_fd_sc_hd__buf_2 output377 (.A(net377),
    .X(W6BEG[8]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net378),
    .X(W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(WW4BEG[0]));
 sky130_fd_sc_hd__buf_2 output380 (.A(net380),
    .X(WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net381),
    .X(WW4BEG[11]));
 sky130_fd_sc_hd__buf_6 output382 (.A(\Inst_LUT4AB_switch_matrix.WW4BEG0 ),
    .X(WW4BEG[12]));
 sky130_fd_sc_hd__buf_8 output383 (.A(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .X(WW4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .X(WW4BEG[14]));
 sky130_fd_sc_hd__buf_8 output385 (.A(\Inst_LUT4AB_switch_matrix.WW4BEG3 ),
    .X(WW4BEG[15]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .X(WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output387 (.A(net387),
    .X(WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output388 (.A(net388),
    .X(WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output389 (.A(net389),
    .X(WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net390),
    .X(WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output391 (.A(net391),
    .X(WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .X(WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output393 (.A(net393),
    .X(WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output394 (.A(net394),
    .X(WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_UserCLK (.A(UserCLK),
    .X(UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_UserCLK_regs (.A(UserCLK_regs),
    .X(clknet_0_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_0__leaf_UserCLK_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_1__leaf_UserCLK_regs));
 sky130_fd_sc_hd__mux2_4 clone8 (.A0(_0337_),
    .A1(_0338_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .X(net402));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer9 (.A(\Inst_LUT4AB_switch_matrix.M_AH ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(net403),
    .X(net404));
 sky130_fd_sc_hd__buf_6 rebuffer11 (.A(\Inst_LUT4AB_switch_matrix.M_AH ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net405),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(\Inst_LUT4AB_switch_matrix.M_AH ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net407),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_1 clone20 (.A(C),
    .X(net414));
 sky130_fd_sc_hd__dlymetal6s2s_1 clone21 (.A(net637),
    .X(net415));
 sky130_fd_sc_hd__buf_8 rebuffer22 (.A(net617),
    .X(net416));
 sky130_fd_sc_hd__buf_6 rebuffer23 (.A(net617),
    .X(net417));
 sky130_fd_sc_hd__buf_6 rebuffer33 (.A(net486),
    .X(net427));
 sky130_fd_sc_hd__buf_6 rebuffer34 (.A(net427),
    .X(net428));
 sky130_fd_sc_hd__buf_8 clone36 (.A(net521),
    .X(net430));
 sky130_fd_sc_hd__buf_6 rebuffer37 (.A(\Inst_LUT4AB_switch_matrix.M_EF ),
    .X(net431));
 sky130_fd_sc_hd__buf_6 rebuffer38 (.A(H),
    .X(net432));
 sky130_fd_sc_hd__buf_8 clone39 (.A(net657),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 clone40 (.A(A),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_2 rebuffer41 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 rebuffer42 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_2 rebuffer43 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 rebuffer44 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_2 rebuffer45 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_2 rebuffer46 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_2 rebuffer47 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_2 rebuffer48 (.A(net447),
    .X(net442));
 sky130_fd_sc_hd__buf_6 rebuffer49 (.A(net481),
    .X(net443));
 sky130_fd_sc_hd__buf_6 clone50 (.A(net639),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 clone51 (.A(D),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 clone52 (.A(net649),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_2 rebuffer53 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_2 rebuffer54 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_2 rebuffer55 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 rebuffer56 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 rebuffer57 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_2 rebuffer58 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 rebuffer59 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_2 rebuffer60 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_2 rebuffer61 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_2 rebuffer62 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer63 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer64 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer65 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer66 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_2 rebuffer67 (.A(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 clone68 (.A(net634),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_1 clone69 (.A(net624),
    .X(net463));
 sky130_fd_sc_hd__buf_6 clone70 (.A(net645),
    .X(net464));
 sky130_fd_sc_hd__dlymetal6s2s_1 clone83 (.A(net637),
    .X(net477));
 sky130_fd_sc_hd__buf_6 clone84 (.A(net636),
    .X(net478));
 sky130_fd_sc_hd__buf_6 rebuffer85 (.A(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_2 rebuffer86 (.A(\Inst_LUT4AB_switch_matrix.M_AB ),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_2 rebuffer87 (.A(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .X(net481));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer88 (.A(net430),
    .X(net482));
 sky130_fd_sc_hd__buf_6 rebuffer89 (.A(net430),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer90 (.A(net635),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer91 (.A(H),
    .X(net485));
 sky130_fd_sc_hd__buf_6 rebuffer92 (.A(H),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer93 (.A(net512),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer94 (.A(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .X(net488));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer95 (.A(net488),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer119 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer120 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer121 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer122 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer123 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer124 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer125 (.A(_0310_),
    .X(net519));
 sky130_fd_sc_hd__buf_6 rebuffer126 (.A(_0310_),
    .X(net520));
 sky130_fd_sc_hd__buf_6 rebuffer127 (.A(\Inst_LUT4AB_switch_matrix.M_AB ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer128 (.A(_0335_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer129 (.A(net402),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer130 (.A(net402),
    .X(net524));
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_417 ();
endmodule
