magic
tech sky130A
magscale 1 2
timestamp 1746770531
<< viali >>
rect 4997 8585 5031 8619
rect 5733 8585 5767 8619
rect 6101 8585 6135 8619
rect 6837 8585 6871 8619
rect 7941 8585 7975 8619
rect 8309 8585 8343 8619
rect 9321 8585 9355 8619
rect 10425 8585 10459 8619
rect 11161 8585 11195 8619
rect 12265 8585 12299 8619
rect 12633 8585 12667 8619
rect 13737 8585 13771 8619
rect 14473 8585 14507 8619
rect 14841 8585 14875 8619
rect 15209 8585 15243 8619
rect 24961 8585 24995 8619
rect 25421 8585 25455 8619
rect 26157 8585 26191 8619
rect 26525 8585 26559 8619
rect 27813 8585 27847 8619
rect 28181 8585 28215 8619
rect 28549 8585 28583 8619
rect 29653 8585 29687 8619
rect 31493 8585 31527 8619
rect 31861 8585 31895 8619
rect 4813 8449 4847 8483
rect 5181 8449 5215 8483
rect 5549 8449 5583 8483
rect 5917 8449 5951 8483
rect 6653 8449 6687 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 7757 8449 7791 8483
rect 8125 8449 8159 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 10609 8449 10643 8483
rect 10989 8449 11023 8483
rect 11345 8449 11379 8483
rect 12081 8449 12115 8483
rect 12449 8449 12483 8483
rect 12817 8449 12851 8483
rect 13185 8449 13219 8483
rect 13553 8449 13587 8483
rect 13921 8449 13955 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 15393 8449 15427 8483
rect 15761 8449 15795 8483
rect 25145 8449 25179 8483
rect 25237 8449 25271 8483
rect 25605 8449 25639 8483
rect 25973 8449 26007 8483
rect 26341 8449 26375 8483
rect 26985 8449 27019 8483
rect 27353 8449 27387 8483
rect 27997 8449 28031 8483
rect 28365 8449 28399 8483
rect 28733 8449 28767 8483
rect 29101 8449 29135 8483
rect 29837 8449 29871 8483
rect 31309 8449 31343 8483
rect 31677 8449 31711 8483
rect 32321 8449 32355 8483
rect 32689 8449 32723 8483
rect 5365 8313 5399 8347
rect 7113 8313 7147 8347
rect 7481 8313 7515 8347
rect 8585 8313 8619 8347
rect 9689 8313 9723 8347
rect 10793 8313 10827 8347
rect 13001 8313 13035 8347
rect 13369 8313 13403 8347
rect 15853 8313 15887 8347
rect 25789 8313 25823 8347
rect 27169 8313 27203 8347
rect 27537 8313 27571 8347
rect 28917 8313 28951 8347
rect 32505 8313 32539 8347
rect 32873 8313 32907 8347
rect 10057 8245 10091 8279
rect 11897 8245 11931 8279
rect 15577 8245 15611 8279
rect 5733 8041 5767 8075
rect 6101 8041 6135 8075
rect 6469 8041 6503 8075
rect 6837 8041 6871 8075
rect 7205 8041 7239 8075
rect 7573 8041 7607 8075
rect 7849 8041 7883 8075
rect 8309 8041 8343 8075
rect 8677 8041 8711 8075
rect 9321 8041 9355 8075
rect 9689 8041 9723 8075
rect 10057 8041 10091 8075
rect 10425 8041 10459 8075
rect 10793 8041 10827 8075
rect 11161 8041 11195 8075
rect 11529 8041 11563 8075
rect 11989 8041 12023 8075
rect 12265 8041 12299 8075
rect 12633 8041 12667 8075
rect 13001 8041 13035 8075
rect 13369 8041 13403 8075
rect 13737 8041 13771 8075
rect 14473 8041 14507 8075
rect 26157 8041 26191 8075
rect 26525 8041 26559 8075
rect 26801 8041 26835 8075
rect 27169 8041 27203 8075
rect 27537 8041 27571 8075
rect 27997 8041 28031 8075
rect 28273 8041 28307 8075
rect 28641 8041 28675 8075
rect 31769 8041 31803 8075
rect 32137 8041 32171 8075
rect 5549 7837 5583 7871
rect 5917 7837 5951 7871
rect 6285 7837 6319 7871
rect 6653 7837 6687 7871
rect 7021 7837 7055 7871
rect 7389 7837 7423 7871
rect 8033 7837 8067 7871
rect 8125 7837 8159 7871
rect 8493 7837 8527 7871
rect 9505 7837 9539 7871
rect 9873 7837 9907 7871
rect 10241 7837 10275 7871
rect 10609 7837 10643 7871
rect 10977 7837 11011 7871
rect 11345 7837 11379 7871
rect 11713 7837 11747 7871
rect 11805 7837 11839 7871
rect 12449 7837 12483 7871
rect 12817 7837 12851 7871
rect 13185 7837 13219 7871
rect 13553 7837 13587 7871
rect 13921 7837 13955 7871
rect 14657 7837 14691 7871
rect 25973 7837 26007 7871
rect 26341 7837 26375 7871
rect 26985 7837 27019 7871
rect 27353 7837 27387 7871
rect 27721 7837 27755 7871
rect 27813 7837 27847 7871
rect 28457 7837 28491 7871
rect 28825 7837 28859 7871
rect 29193 7837 29227 7871
rect 31585 7837 31619 7871
rect 31953 7837 31987 7871
rect 32321 7837 32355 7871
rect 32689 7837 32723 7871
rect 29009 7701 29043 7735
rect 32505 7701 32539 7735
rect 32873 7701 32907 7735
rect 2513 7497 2547 7531
rect 2789 7497 2823 7531
rect 3341 7497 3375 7531
rect 7389 7497 7423 7531
rect 9413 7497 9447 7531
rect 9873 7497 9907 7531
rect 11345 7497 11379 7531
rect 11989 7497 12023 7531
rect 12265 7497 12299 7531
rect 12541 7497 12575 7531
rect 12817 7497 12851 7531
rect 16405 7497 16439 7531
rect 17049 7497 17083 7531
rect 17417 7497 17451 7531
rect 18521 7497 18555 7531
rect 18797 7497 18831 7531
rect 19533 7497 19567 7531
rect 19809 7497 19843 7531
rect 20729 7497 20763 7531
rect 21097 7497 21131 7531
rect 21373 7497 21407 7531
rect 27813 7497 27847 7531
rect 28549 7497 28583 7531
rect 28917 7497 28951 7531
rect 29193 7497 29227 7531
rect 29745 7497 29779 7531
rect 30665 7497 30699 7531
rect 32505 7497 32539 7531
rect 2145 7361 2179 7395
rect 2513 7361 2547 7395
rect 2605 7361 2639 7395
rect 2881 7361 2915 7395
rect 3157 7361 3191 7395
rect 7205 7361 7239 7395
rect 9229 7361 9263 7395
rect 10057 7361 10091 7395
rect 11161 7361 11195 7395
rect 11897 7361 11931 7395
rect 12181 7361 12215 7395
rect 12449 7361 12483 7395
rect 12725 7361 12759 7395
rect 13001 7361 13035 7395
rect 16497 7361 16531 7395
rect 16773 7361 16807 7395
rect 17141 7361 17175 7395
rect 17233 7361 17267 7395
rect 18245 7361 18279 7395
rect 18337 7361 18371 7395
rect 18613 7361 18647 7395
rect 18889 7361 18923 7395
rect 19257 7361 19291 7395
rect 19349 7361 19383 7395
rect 19625 7361 19659 7395
rect 19993 7361 20027 7395
rect 20453 7361 20487 7395
rect 20821 7361 20855 7395
rect 20913 7361 20947 7395
rect 21189 7361 21223 7395
rect 27997 7361 28031 7395
rect 28365 7361 28399 7395
rect 28825 7361 28859 7395
rect 29101 7361 29135 7395
rect 29377 7361 29411 7395
rect 29929 7361 29963 7395
rect 30205 7361 30239 7395
rect 30849 7361 30883 7395
rect 32321 7361 32355 7395
rect 32689 7361 32723 7395
rect 2329 7225 2363 7259
rect 3065 7225 3099 7259
rect 11713 7225 11747 7259
rect 16957 7225 16991 7259
rect 18153 7225 18187 7259
rect 20177 7225 20211 7259
rect 20637 7225 20671 7259
rect 28641 7225 28675 7259
rect 30021 7225 30055 7259
rect 19165 7157 19199 7191
rect 21465 7157 21499 7191
rect 32873 7157 32907 7191
rect 3985 6953 4019 6987
rect 12081 6953 12115 6987
rect 3157 6749 3191 6783
rect 3433 6749 3467 6783
rect 3801 6749 3835 6783
rect 4077 6749 4111 6783
rect 7205 6749 7239 6783
rect 12265 6749 12299 6783
rect 12541 6749 12575 6783
rect 24133 6749 24167 6783
rect 24593 6749 24627 6783
rect 24869 6749 24903 6783
rect 25145 6749 25179 6783
rect 25605 6749 25639 6783
rect 25973 6749 26007 6783
rect 26341 6749 26375 6783
rect 26709 6749 26743 6783
rect 26985 6749 27019 6783
rect 29285 6749 29319 6783
rect 32321 6749 32355 6783
rect 32689 6749 32723 6783
rect 3341 6613 3375 6647
rect 3617 6613 3651 6647
rect 4261 6613 4295 6647
rect 7389 6613 7423 6647
rect 12357 6613 12391 6647
rect 23949 6613 23983 6647
rect 24409 6613 24443 6647
rect 24685 6613 24719 6647
rect 24961 6613 24995 6647
rect 25421 6613 25455 6647
rect 25789 6613 25823 6647
rect 26157 6613 26191 6647
rect 26525 6613 26559 6647
rect 26801 6613 26835 6647
rect 29101 6613 29135 6647
rect 32505 6613 32539 6647
rect 32873 6613 32907 6647
rect 3985 6409 4019 6443
rect 4997 6409 5031 6443
rect 6745 6409 6779 6443
rect 6929 6409 6963 6443
rect 7205 6409 7239 6443
rect 7481 6409 7515 6443
rect 7573 6409 7607 6443
rect 8125 6409 8159 6443
rect 8401 6409 8435 6443
rect 13737 6409 13771 6443
rect 15117 6409 15151 6443
rect 22661 6409 22695 6443
rect 32873 6409 32907 6443
rect 13277 6341 13311 6375
rect 15485 6341 15519 6375
rect 3985 6273 4019 6307
rect 4077 6273 4111 6307
rect 4537 6273 4571 6307
rect 4813 6273 4847 6307
rect 5089 6273 5123 6307
rect 6561 6273 6595 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 7757 6273 7791 6307
rect 8309 6273 8343 6307
rect 8585 6273 8619 6307
rect 13093 6273 13127 6307
rect 13553 6273 13587 6307
rect 13829 6273 13863 6307
rect 14105 6273 14139 6307
rect 14381 6273 14415 6307
rect 14657 6273 14691 6307
rect 14933 6273 14967 6307
rect 15209 6273 15243 6307
rect 15669 6273 15703 6307
rect 21649 6273 21683 6307
rect 22025 6273 22059 6307
rect 22293 6273 22327 6307
rect 22569 6273 22603 6307
rect 22845 6273 22879 6307
rect 23121 6273 23155 6307
rect 23397 6273 23431 6307
rect 32321 6273 32355 6307
rect 32689 6273 32723 6307
rect 8033 6205 8067 6239
rect 12909 6205 12943 6239
rect 13461 6205 13495 6239
rect 15853 6205 15887 6239
rect 4261 6137 4295 6171
rect 5273 6137 5307 6171
rect 15393 6137 15427 6171
rect 22109 6137 22143 6171
rect 22385 6137 22419 6171
rect 22937 6137 22971 6171
rect 4721 6069 4755 6103
rect 12817 6069 12851 6103
rect 13001 6069 13035 6103
rect 13185 6069 13219 6103
rect 13369 6069 13403 6103
rect 14013 6069 14047 6103
rect 14289 6069 14323 6103
rect 14565 6069 14599 6103
rect 14841 6069 14875 6103
rect 15669 6069 15703 6103
rect 21465 6069 21499 6103
rect 21833 6069 21867 6103
rect 23213 6069 23247 6103
rect 32505 6069 32539 6103
rect 7481 5865 7515 5899
rect 17325 5797 17359 5831
rect 32873 5797 32907 5831
rect 7297 5661 7331 5695
rect 15577 5661 15611 5695
rect 15669 5661 15703 5695
rect 16681 5661 16715 5695
rect 17049 5661 17083 5695
rect 17141 5661 17175 5695
rect 17417 5661 17451 5695
rect 17693 5661 17727 5695
rect 32321 5661 32355 5695
rect 32689 5661 32723 5695
rect 16957 5593 16991 5627
rect 15485 5525 15519 5559
rect 15853 5525 15887 5559
rect 16865 5525 16899 5559
rect 17601 5525 17635 5559
rect 32505 5525 32539 5559
rect 32873 5321 32907 5355
rect 17233 5253 17267 5287
rect 17049 5185 17083 5219
rect 17325 5185 17359 5219
rect 17601 5185 17635 5219
rect 17877 5185 17911 5219
rect 18153 5185 18187 5219
rect 18429 5185 18463 5219
rect 18889 5185 18923 5219
rect 32321 5185 32355 5219
rect 32689 5185 32723 5219
rect 16865 5117 16899 5151
rect 18705 5117 18739 5151
rect 17141 5049 17175 5083
rect 17785 5049 17819 5083
rect 18613 5049 18647 5083
rect 16773 4981 16807 5015
rect 16957 4981 16991 5015
rect 17509 4981 17543 5015
rect 18061 4981 18095 5015
rect 18337 4981 18371 5015
rect 32505 4981 32539 5015
rect 11897 4777 11931 4811
rect 28825 4777 28859 4811
rect 32873 4709 32907 4743
rect 12081 4573 12115 4607
rect 14105 4573 14139 4607
rect 28733 4573 28767 4607
rect 29009 4573 29043 4607
rect 32321 4573 32355 4607
rect 32689 4573 32723 4607
rect 14289 4437 14323 4471
rect 28641 4437 28675 4471
rect 32505 4437 32539 4471
rect 12909 4233 12943 4267
rect 7573 4097 7607 4131
rect 11713 4097 11747 4131
rect 11989 4097 12023 4131
rect 12265 4097 12299 4131
rect 12541 4097 12575 4131
rect 12817 4097 12851 4131
rect 13093 4097 13127 4131
rect 32321 4097 32355 4131
rect 32689 4097 32723 4131
rect 11529 3961 11563 3995
rect 12081 3961 12115 3995
rect 12633 3961 12667 3995
rect 32873 3961 32907 3995
rect 7757 3893 7791 3927
rect 11805 3893 11839 3927
rect 12357 3893 12391 3927
rect 32505 3893 32539 3927
rect 10517 3689 10551 3723
rect 12081 3689 12115 3723
rect 14473 3689 14507 3723
rect 15393 3689 15427 3723
rect 18061 3689 18095 3723
rect 19809 3689 19843 3723
rect 20637 3689 20671 3723
rect 21097 3689 21131 3723
rect 23213 3689 23247 3723
rect 27261 3689 27295 3723
rect 28917 3689 28951 3723
rect 11345 3621 11379 3655
rect 17785 3621 17819 3655
rect 19441 3621 19475 3655
rect 20177 3621 20211 3655
rect 29653 3621 29687 3655
rect 32873 3621 32907 3655
rect 10333 3485 10367 3519
rect 11161 3485 11195 3519
rect 12265 3485 12299 3519
rect 14289 3485 14323 3519
rect 15485 3485 15519 3519
rect 15577 3485 15611 3519
rect 17601 3485 17635 3519
rect 17877 3485 17911 3519
rect 19257 3485 19291 3519
rect 19901 3485 19935 3519
rect 19993 3485 20027 3519
rect 20453 3485 20487 3519
rect 20913 3485 20947 3519
rect 21465 3485 21499 3519
rect 21557 3485 21591 3519
rect 22937 3485 22971 3519
rect 23029 3485 23063 3519
rect 27077 3485 27111 3519
rect 29101 3485 29135 3519
rect 29837 3485 29871 3519
rect 32321 3485 32355 3519
rect 32689 3485 32723 3519
rect 15761 3349 15795 3383
rect 21373 3349 21407 3383
rect 21741 3349 21775 3383
rect 22845 3349 22879 3383
rect 32505 3349 32539 3383
rect 32873 3145 32907 3179
rect 31677 3009 31711 3043
rect 32321 3009 32355 3043
rect 32689 3009 32723 3043
rect 31861 2805 31895 2839
rect 32505 2805 32539 2839
rect 32873 2533 32907 2567
rect 30941 2397 30975 2431
rect 31309 2397 31343 2431
rect 31677 2397 31711 2431
rect 32321 2397 32355 2431
rect 32689 2397 32723 2431
rect 31125 2261 31159 2295
rect 31493 2261 31527 2295
rect 31861 2261 31895 2295
rect 32505 2261 32539 2295
<< metal1 >>
rect 7558 11092 7564 11144
rect 7616 11132 7622 11144
rect 18046 11132 18052 11144
rect 7616 11104 18052 11132
rect 7616 11092 7622 11104
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7064 11036 18000 11064
rect 7064 11024 7070 11036
rect 17972 11008 18000 11036
rect 17954 10956 17960 11008
rect 18012 10956 18018 11008
rect 9582 10820 9588 10872
rect 9640 10860 9646 10872
rect 18690 10860 18696 10872
rect 9640 10832 18696 10860
rect 9640 10820 9646 10832
rect 18690 10820 18696 10832
rect 18748 10820 18754 10872
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 16114 10656 16120 10668
rect 10744 10628 16120 10656
rect 10744 10616 10750 10628
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 15746 10588 15752 10600
rect 14424 10560 15752 10588
rect 14424 10548 14430 10560
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 17770 10520 17776 10532
rect 12032 10492 17776 10520
rect 12032 10480 12038 10492
rect 17770 10480 17776 10492
rect 17828 10480 17834 10532
rect 13262 10140 13268 10192
rect 13320 10180 13326 10192
rect 19794 10180 19800 10192
rect 13320 10152 19800 10180
rect 13320 10140 13326 10152
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 16666 9936 16672 9988
rect 16724 9976 16730 9988
rect 20162 9976 20168 9988
rect 16724 9948 20168 9976
rect 16724 9936 16730 9948
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 13630 9732 13636 9784
rect 13688 9772 13694 9784
rect 19242 9772 19248 9784
rect 13688 9744 19248 9772
rect 13688 9732 13694 9744
rect 19242 9732 19248 9744
rect 19300 9732 19306 9784
rect 18414 9596 18420 9648
rect 18472 9636 18478 9648
rect 20714 9636 20720 9648
rect 18472 9608 20720 9636
rect 18472 9596 18478 9608
rect 20714 9596 20720 9608
rect 20772 9596 20778 9648
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 26694 9568 26700 9580
rect 15712 9540 26700 9568
rect 15712 9528 15718 9540
rect 26694 9528 26700 9540
rect 26752 9528 26758 9580
rect 13446 9460 13452 9512
rect 13504 9500 13510 9512
rect 24394 9500 24400 9512
rect 13504 9472 24400 9500
rect 13504 9460 13510 9472
rect 24394 9460 24400 9472
rect 24452 9460 24458 9512
rect 8662 9392 8668 9444
rect 8720 9432 8726 9444
rect 9306 9432 9312 9444
rect 8720 9404 9312 9432
rect 8720 9392 8726 9404
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 31662 9432 31668 9444
rect 19576 9404 31668 9432
rect 19576 9392 19582 9404
rect 31662 9392 31668 9404
rect 31720 9392 31726 9444
rect 1302 9324 1308 9376
rect 1360 9364 1366 9376
rect 19702 9364 19708 9376
rect 1360 9336 19708 9364
rect 1360 9324 1366 9336
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 1026 9256 1032 9308
rect 1084 9296 1090 9308
rect 19610 9296 19616 9308
rect 1084 9268 19616 9296
rect 1084 9256 1090 9268
rect 19610 9256 19616 9268
rect 19668 9256 19674 9308
rect 19794 9256 19800 9308
rect 19852 9296 19858 9308
rect 32306 9296 32312 9308
rect 19852 9268 32312 9296
rect 19852 9256 19858 9268
rect 32306 9256 32312 9268
rect 32364 9256 32370 9308
rect 13814 9188 13820 9240
rect 13872 9228 13878 9240
rect 24670 9228 24676 9240
rect 13872 9200 24676 9228
rect 13872 9188 13878 9200
rect 24670 9188 24676 9200
rect 24728 9188 24734 9240
rect 21082 9120 21088 9172
rect 21140 9160 21146 9172
rect 21726 9160 21732 9172
rect 21140 9132 21732 9160
rect 21140 9120 21146 9132
rect 21726 9120 21732 9132
rect 21784 9120 21790 9172
rect 290 8984 296 9036
rect 348 9024 354 9036
rect 20438 9024 20444 9036
rect 348 8996 20444 9024
rect 348 8984 354 8996
rect 20438 8984 20444 8996
rect 20496 8984 20502 9036
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 12526 8956 12532 8968
rect 10376 8928 12532 8956
rect 10376 8916 10382 8928
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 18046 8956 18052 8968
rect 12952 8928 18052 8956
rect 12952 8916 12958 8928
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 22738 8916 22744 8968
rect 22796 8956 22802 8968
rect 25590 8956 25596 8968
rect 22796 8928 25596 8956
rect 22796 8916 22802 8928
rect 25590 8916 25596 8928
rect 25648 8916 25654 8968
rect 27522 8916 27528 8968
rect 27580 8956 27586 8968
rect 28534 8956 28540 8968
rect 27580 8928 28540 8956
rect 27580 8916 27586 8928
rect 28534 8916 28540 8928
rect 28592 8916 28598 8968
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7926 8888 7932 8900
rect 7248 8860 7932 8888
rect 7248 8848 7254 8860
rect 7926 8848 7932 8860
rect 7984 8848 7990 8900
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 10778 8888 10784 8900
rect 10192 8860 10784 8888
rect 10192 8848 10198 8860
rect 10778 8848 10784 8860
rect 10836 8848 10842 8900
rect 10870 8848 10876 8900
rect 10928 8888 10934 8900
rect 12158 8888 12164 8900
rect 10928 8860 12164 8888
rect 10928 8848 10934 8860
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 12986 8888 12992 8900
rect 12400 8860 12992 8888
rect 12400 8848 12406 8860
rect 12986 8848 12992 8860
rect 13044 8848 13050 8900
rect 20898 8888 20904 8900
rect 14476 8860 20904 8888
rect 6454 8780 6460 8832
rect 6512 8820 6518 8832
rect 8110 8820 8116 8832
rect 6512 8792 8116 8820
rect 6512 8780 6518 8792
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 11146 8820 11152 8832
rect 10560 8792 11152 8820
rect 10560 8780 10566 8792
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 12710 8780 12716 8832
rect 12768 8820 12774 8832
rect 14476 8820 14504 8860
rect 20898 8848 20904 8860
rect 20956 8848 20962 8900
rect 21358 8848 21364 8900
rect 21416 8888 21422 8900
rect 32674 8888 32680 8900
rect 21416 8860 32680 8888
rect 21416 8848 21422 8860
rect 32674 8848 32680 8860
rect 32732 8848 32738 8900
rect 12768 8792 14504 8820
rect 12768 8780 12774 8792
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 25038 8820 25044 8832
rect 14608 8792 25044 8820
rect 14608 8780 14614 8792
rect 25038 8780 25044 8792
rect 25096 8780 25102 8832
rect 27154 8780 27160 8832
rect 27212 8820 27218 8832
rect 27522 8820 27528 8832
rect 27212 8792 27528 8820
rect 27212 8780 27218 8792
rect 27522 8780 27528 8792
rect 27580 8780 27586 8832
rect 1104 8730 33324 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 33324 8730
rect 1104 8656 33324 8678
rect 4985 8619 5043 8625
rect 4985 8585 4997 8619
rect 5031 8616 5043 8619
rect 5626 8616 5632 8628
rect 5031 8588 5632 8616
rect 5031 8585 5043 8588
rect 4985 8579 5043 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 6730 8616 6736 8628
rect 6135 8588 6736 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 5736 8548 5764 8579
rect 6730 8576 6736 8588
rect 6788 8576 6794 8628
rect 6825 8619 6883 8625
rect 6825 8585 6837 8619
rect 6871 8616 6883 8619
rect 7466 8616 7472 8628
rect 6871 8588 7472 8616
rect 6871 8585 6883 8588
rect 6825 8579 6883 8585
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 7742 8576 7748 8628
rect 7800 8576 7806 8628
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8846 8616 8852 8628
rect 8343 8588 8852 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 6362 8548 6368 8560
rect 5736 8520 6368 8548
rect 6362 8508 6368 8520
rect 6420 8508 6426 8560
rect 7760 8548 7788 8576
rect 7116 8520 7788 8548
rect 7944 8548 7972 8579
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 10042 8616 10048 8628
rect 9355 8588 10048 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10502 8616 10508 8628
rect 10459 8588 10508 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 11054 8616 11060 8628
rect 10796 8588 11060 8616
rect 8570 8548 8576 8560
rect 7944 8520 8576 8548
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 5166 8440 5172 8492
rect 5224 8440 5230 8492
rect 5258 8440 5264 8492
rect 5316 8480 5322 8492
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 5316 8452 5549 8480
rect 5316 8440 5322 8452
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5537 8443 5595 8449
rect 5644 8452 5917 8480
rect 5442 8372 5448 8424
rect 5500 8412 5506 8424
rect 5644 8412 5672 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 5500 8384 5672 8412
rect 5500 8372 5506 8384
rect 4154 8304 4160 8356
rect 4212 8344 4218 8356
rect 5353 8347 5411 8353
rect 4212 8316 5304 8344
rect 4212 8304 4218 8316
rect 5276 8276 5304 8316
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 5994 8344 6000 8356
rect 5399 8316 6000 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 5994 8304 6000 8316
rect 6052 8304 6058 8356
rect 6656 8344 6684 8443
rect 7116 8353 7144 8520
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 10318 8548 10324 8560
rect 8772 8520 10324 8548
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 7466 8480 7472 8492
rect 7331 8452 7472 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 7926 8480 7932 8492
rect 7791 8452 7932 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 7558 8412 7564 8424
rect 7432 8384 7564 8412
rect 7432 8372 7438 8384
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 7668 8412 7696 8443
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 8110 8440 8116 8492
rect 8168 8440 8174 8492
rect 8772 8489 8800 8520
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 10796 8548 10824 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11882 8616 11888 8628
rect 11195 8588 11888 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12342 8616 12348 8628
rect 12299 8588 12348 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 12621 8619 12679 8625
rect 12621 8585 12633 8619
rect 12667 8616 12679 8619
rect 13354 8616 13360 8628
rect 12667 8588 13360 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 14090 8616 14096 8628
rect 13771 8588 14096 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 14458 8576 14464 8628
rect 14516 8576 14522 8628
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 14700 8588 14841 8616
rect 14700 8576 14706 8588
rect 14829 8585 14841 8588
rect 14875 8585 14887 8619
rect 14829 8579 14887 8585
rect 14918 8576 14924 8628
rect 14976 8616 14982 8628
rect 15197 8619 15255 8625
rect 15197 8616 15209 8619
rect 14976 8588 15209 8616
rect 14976 8576 14982 8588
rect 15197 8585 15209 8588
rect 15243 8585 15255 8619
rect 15197 8579 15255 8585
rect 18340 8588 22094 8616
rect 12710 8548 12716 8560
rect 10520 8520 10824 8548
rect 12084 8520 12716 8548
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9766 8480 9772 8492
rect 9539 8452 9772 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10520 8480 10548 8520
rect 10275 8452 10548 8480
rect 10597 8483 10655 8489
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 10778 8480 10784 8492
rect 10643 8452 10784 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 9876 8412 9904 8443
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 10977 8483 11035 8489
rect 10977 8449 10989 8483
rect 11023 8480 11035 8483
rect 11238 8480 11244 8492
rect 11023 8452 11244 8480
rect 11023 8449 11035 8452
rect 10977 8443 11035 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 11606 8480 11612 8492
rect 11379 8452 11612 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 12084 8489 12112 8520
rect 12710 8508 12716 8520
rect 12768 8508 12774 8560
rect 18340 8548 18368 8588
rect 14660 8520 18368 8548
rect 22066 8548 22094 8588
rect 24946 8576 24952 8628
rect 25004 8576 25010 8628
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 25409 8619 25467 8625
rect 25409 8616 25421 8619
rect 25188 8588 25421 8616
rect 25188 8576 25194 8588
rect 25409 8585 25421 8588
rect 25455 8585 25467 8619
rect 25409 8579 25467 8585
rect 25498 8576 25504 8628
rect 25556 8616 25562 8628
rect 26145 8619 26203 8625
rect 26145 8616 26157 8619
rect 25556 8588 26157 8616
rect 25556 8576 25562 8588
rect 26145 8585 26157 8588
rect 26191 8585 26203 8619
rect 26145 8579 26203 8585
rect 26513 8619 26571 8625
rect 26513 8585 26525 8619
rect 26559 8585 26571 8619
rect 26513 8579 26571 8585
rect 22066 8520 25544 8548
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12805 8483 12863 8489
rect 12483 8452 12756 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 10318 8412 10324 8424
rect 7668 8384 7788 8412
rect 9876 8384 10324 8412
rect 7760 8356 7788 8384
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 6104 8316 6684 8344
rect 7101 8347 7159 8353
rect 6104 8276 6132 8316
rect 7101 8313 7113 8347
rect 7147 8313 7159 8347
rect 7101 8307 7159 8313
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8344 7527 8347
rect 7515 8316 7604 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 5276 8248 6132 8276
rect 7576 8276 7604 8316
rect 7742 8304 7748 8356
rect 7800 8304 7806 8356
rect 8202 8344 8208 8356
rect 7852 8316 8208 8344
rect 7852 8276 7880 8316
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8573 8347 8631 8353
rect 8573 8313 8585 8347
rect 8619 8344 8631 8347
rect 8662 8344 8668 8356
rect 8619 8316 8668 8344
rect 8619 8313 8631 8316
rect 8573 8307 8631 8313
rect 8662 8304 8668 8316
rect 8720 8304 8726 8356
rect 9677 8347 9735 8353
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 10410 8344 10416 8356
rect 9723 8316 10416 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 10781 8347 10839 8353
rect 10781 8313 10793 8347
rect 10827 8344 10839 8347
rect 11514 8344 11520 8356
rect 10827 8316 11520 8344
rect 10827 8313 10839 8316
rect 10781 8307 10839 8313
rect 11514 8304 11520 8316
rect 11572 8304 11578 8356
rect 7576 8248 7880 8276
rect 10042 8236 10048 8288
rect 10100 8236 10106 8288
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11422 8276 11428 8288
rect 11204 8248 11428 8276
rect 11204 8236 11210 8248
rect 11422 8236 11428 8248
rect 11480 8236 11486 8288
rect 11885 8279 11943 8285
rect 11885 8245 11897 8279
rect 11931 8276 11943 8279
rect 12618 8276 12624 8288
rect 11931 8248 12624 8276
rect 11931 8245 11943 8248
rect 11885 8239 11943 8245
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 12728 8276 12756 8452
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 12894 8480 12900 8492
rect 12851 8452 12900 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13446 8480 13452 8492
rect 13219 8452 13452 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8480 13599 8483
rect 13814 8480 13820 8492
rect 13587 8452 13820 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 14550 8480 14556 8492
rect 13955 8452 14556 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14660 8489 14688 8520
rect 25516 8492 25544 8520
rect 25682 8508 25688 8560
rect 25740 8548 25746 8560
rect 26528 8548 26556 8579
rect 26786 8576 26792 8628
rect 26844 8616 26850 8628
rect 27801 8619 27859 8625
rect 27801 8616 27813 8619
rect 26844 8588 27813 8616
rect 26844 8576 26850 8588
rect 27801 8585 27813 8588
rect 27847 8585 27859 8619
rect 27801 8579 27859 8585
rect 28169 8619 28227 8625
rect 28169 8585 28181 8619
rect 28215 8585 28227 8619
rect 28169 8579 28227 8585
rect 25740 8520 26556 8548
rect 26988 8520 27476 8548
rect 25740 8508 25746 8520
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14976 8452 15025 8480
rect 14976 8440 14982 8452
rect 15013 8449 15025 8452
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8480 15439 8483
rect 15654 8480 15660 8492
rect 15427 8452 15660 8480
rect 15427 8449 15439 8452
rect 15381 8443 15439 8449
rect 15654 8440 15660 8452
rect 15712 8440 15718 8492
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8480 15807 8483
rect 24486 8480 24492 8492
rect 15795 8452 24492 8480
rect 15795 8449 15807 8452
rect 15749 8443 15807 8449
rect 24486 8440 24492 8452
rect 24544 8440 24550 8492
rect 25130 8440 25136 8492
rect 25188 8440 25194 8492
rect 25222 8440 25228 8492
rect 25280 8440 25286 8492
rect 25498 8440 25504 8492
rect 25556 8440 25562 8492
rect 25593 8483 25651 8489
rect 25593 8449 25605 8483
rect 25639 8449 25651 8483
rect 25593 8443 25651 8449
rect 13722 8412 13728 8424
rect 13280 8384 13728 8412
rect 12989 8347 13047 8353
rect 12989 8313 13001 8347
rect 13035 8344 13047 8347
rect 13280 8344 13308 8384
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 22646 8372 22652 8424
rect 22704 8412 22710 8424
rect 25608 8412 25636 8443
rect 25774 8440 25780 8492
rect 25832 8480 25838 8492
rect 25961 8483 26019 8489
rect 25961 8480 25973 8483
rect 25832 8452 25973 8480
rect 25832 8440 25838 8452
rect 25961 8449 25973 8452
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 26329 8483 26387 8489
rect 26329 8449 26341 8483
rect 26375 8480 26387 8483
rect 26418 8480 26424 8492
rect 26375 8452 26424 8480
rect 26375 8449 26387 8452
rect 26329 8443 26387 8449
rect 26418 8440 26424 8452
rect 26476 8440 26482 8492
rect 26988 8489 27016 8520
rect 26973 8483 27031 8489
rect 26973 8449 26985 8483
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27338 8440 27344 8492
rect 27396 8440 27402 8492
rect 27448 8480 27476 8520
rect 27522 8508 27528 8560
rect 27580 8548 27586 8560
rect 28184 8548 28212 8579
rect 28534 8576 28540 8628
rect 28592 8576 28598 8628
rect 28626 8576 28632 8628
rect 28684 8616 28690 8628
rect 29641 8619 29699 8625
rect 29641 8616 29653 8619
rect 28684 8588 29653 8616
rect 28684 8576 28690 8588
rect 29641 8585 29653 8588
rect 29687 8585 29699 8619
rect 29641 8579 29699 8585
rect 31478 8576 31484 8628
rect 31536 8576 31542 8628
rect 31846 8576 31852 8628
rect 31904 8576 31910 8628
rect 27580 8520 28212 8548
rect 27580 8508 27586 8520
rect 27614 8480 27620 8492
rect 27448 8452 27620 8480
rect 27614 8440 27620 8452
rect 27672 8440 27678 8492
rect 27982 8440 27988 8492
rect 28040 8440 28046 8492
rect 28353 8483 28411 8489
rect 28353 8449 28365 8483
rect 28399 8480 28411 8483
rect 28626 8480 28632 8492
rect 28399 8452 28632 8480
rect 28399 8449 28411 8452
rect 28353 8443 28411 8449
rect 28626 8440 28632 8452
rect 28684 8440 28690 8492
rect 28718 8440 28724 8492
rect 28776 8440 28782 8492
rect 28902 8440 28908 8492
rect 28960 8480 28966 8492
rect 29089 8483 29147 8489
rect 29089 8480 29101 8483
rect 28960 8452 29101 8480
rect 28960 8440 28966 8452
rect 29089 8449 29101 8452
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 29822 8440 29828 8492
rect 29880 8440 29886 8492
rect 31294 8440 31300 8492
rect 31352 8440 31358 8492
rect 31662 8440 31668 8492
rect 31720 8440 31726 8492
rect 32306 8440 32312 8492
rect 32364 8440 32370 8492
rect 32674 8440 32680 8492
rect 32732 8440 32738 8492
rect 22704 8384 25636 8412
rect 22704 8372 22710 8384
rect 26510 8372 26516 8424
rect 26568 8412 26574 8424
rect 26568 8384 27568 8412
rect 26568 8372 26574 8384
rect 13035 8316 13308 8344
rect 13357 8347 13415 8353
rect 13035 8313 13047 8316
rect 12989 8307 13047 8313
rect 13357 8313 13369 8347
rect 13403 8344 13415 8347
rect 13814 8344 13820 8356
rect 13403 8316 13820 8344
rect 13403 8313 13415 8316
rect 13357 8307 13415 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 14826 8304 14832 8356
rect 14884 8344 14890 8356
rect 14884 8316 15332 8344
rect 14884 8304 14890 8316
rect 14550 8276 14556 8288
rect 12728 8248 14556 8276
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 15304 8276 15332 8316
rect 15378 8304 15384 8356
rect 15436 8344 15442 8356
rect 15841 8347 15899 8353
rect 15841 8344 15853 8347
rect 15436 8316 15853 8344
rect 15436 8304 15442 8316
rect 15841 8313 15853 8316
rect 15887 8313 15899 8347
rect 15841 8307 15899 8313
rect 22922 8304 22928 8356
rect 22980 8344 22986 8356
rect 25130 8344 25136 8356
rect 22980 8316 25136 8344
rect 22980 8304 22986 8316
rect 25130 8304 25136 8316
rect 25188 8304 25194 8356
rect 25314 8304 25320 8356
rect 25372 8344 25378 8356
rect 25777 8347 25835 8353
rect 25777 8344 25789 8347
rect 25372 8316 25789 8344
rect 25372 8304 25378 8316
rect 25777 8313 25789 8316
rect 25823 8313 25835 8347
rect 25777 8307 25835 8313
rect 26050 8304 26056 8356
rect 26108 8344 26114 8356
rect 27540 8353 27568 8384
rect 27157 8347 27215 8353
rect 27157 8344 27169 8347
rect 26108 8316 27169 8344
rect 26108 8304 26114 8316
rect 27157 8313 27169 8316
rect 27203 8313 27215 8347
rect 27157 8307 27215 8313
rect 27525 8347 27583 8353
rect 27525 8313 27537 8347
rect 27571 8313 27583 8347
rect 27525 8307 27583 8313
rect 27890 8304 27896 8356
rect 27948 8344 27954 8356
rect 28905 8347 28963 8353
rect 28905 8344 28917 8347
rect 27948 8316 28917 8344
rect 27948 8304 27954 8316
rect 28905 8313 28917 8316
rect 28951 8313 28963 8347
rect 28905 8307 28963 8313
rect 32490 8304 32496 8356
rect 32548 8304 32554 8356
rect 32858 8304 32864 8356
rect 32916 8304 32922 8356
rect 15565 8279 15623 8285
rect 15565 8276 15577 8279
rect 15304 8248 15577 8276
rect 15565 8245 15577 8248
rect 15611 8245 15623 8279
rect 15565 8239 15623 8245
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 19978 8276 19984 8288
rect 16264 8248 19984 8276
rect 16264 8236 16270 8248
rect 19978 8236 19984 8248
rect 20036 8236 20042 8288
rect 24762 8236 24768 8288
rect 24820 8276 24826 8288
rect 31662 8276 31668 8288
rect 24820 8248 31668 8276
rect 24820 8236 24826 8248
rect 31662 8236 31668 8248
rect 31720 8236 31726 8288
rect 1104 8186 33304 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 33304 8186
rect 1104 8112 33304 8134
rect 5721 8075 5779 8081
rect 5721 8041 5733 8075
rect 5767 8072 5779 8075
rect 5810 8072 5816 8084
rect 5767 8044 5816 8072
rect 5767 8041 5779 8044
rect 5721 8035 5779 8041
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 6089 8075 6147 8081
rect 6089 8041 6101 8075
rect 6135 8072 6147 8075
rect 6178 8072 6184 8084
rect 6135 8044 6184 8072
rect 6135 8041 6147 8044
rect 6089 8035 6147 8041
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 6546 8072 6552 8084
rect 6503 8044 6552 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6825 8075 6883 8081
rect 6825 8041 6837 8075
rect 6871 8072 6883 8075
rect 6914 8072 6920 8084
rect 6871 8044 6920 8072
rect 6871 8041 6883 8044
rect 6825 8035 6883 8041
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7282 8072 7288 8084
rect 7239 8044 7288 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7561 8075 7619 8081
rect 7561 8041 7573 8075
rect 7607 8072 7619 8075
rect 7650 8072 7656 8084
rect 7607 8044 7656 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 7834 8032 7840 8084
rect 7892 8032 7898 8084
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8386 8072 8392 8084
rect 8343 8044 8392 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8665 8075 8723 8081
rect 8665 8041 8677 8075
rect 8711 8072 8723 8075
rect 8754 8072 8760 8084
rect 8711 8044 8760 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 9309 8075 9367 8081
rect 9309 8041 9321 8075
rect 9355 8072 9367 8075
rect 9490 8072 9496 8084
rect 9355 8044 9496 8072
rect 9355 8041 9367 8044
rect 9309 8035 9367 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 9677 8075 9735 8081
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 9858 8072 9864 8084
rect 9723 8044 9864 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10226 8072 10232 8084
rect 10091 8044 10232 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 10413 8075 10471 8081
rect 10413 8041 10425 8075
rect 10459 8072 10471 8075
rect 10594 8072 10600 8084
rect 10459 8044 10600 8072
rect 10459 8041 10471 8044
rect 10413 8035 10471 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 10781 8075 10839 8081
rect 10781 8041 10793 8075
rect 10827 8072 10839 8075
rect 10962 8072 10968 8084
rect 10827 8044 10968 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11149 8075 11207 8081
rect 11149 8041 11161 8075
rect 11195 8072 11207 8075
rect 11330 8072 11336 8084
rect 11195 8044 11336 8072
rect 11195 8041 11207 8044
rect 11149 8035 11207 8041
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 11698 8072 11704 8084
rect 11563 8044 11704 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 11977 8075 12035 8081
rect 11977 8041 11989 8075
rect 12023 8072 12035 8075
rect 12066 8072 12072 8084
rect 12023 8044 12072 8072
rect 12023 8041 12035 8044
rect 11977 8035 12035 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12250 8032 12256 8084
rect 12308 8032 12314 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12492 8044 12633 8072
rect 12492 8032 12498 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12860 8044 13001 8072
rect 12860 8032 12866 8044
rect 12989 8041 13001 8044
rect 13035 8041 13047 8075
rect 12989 8035 13047 8041
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 13357 8075 13415 8081
rect 13357 8072 13369 8075
rect 13228 8044 13369 8072
rect 13228 8032 13234 8044
rect 13357 8041 13369 8044
rect 13403 8041 13415 8075
rect 13357 8035 13415 8041
rect 13538 8032 13544 8084
rect 13596 8072 13602 8084
rect 13725 8075 13783 8081
rect 13725 8072 13737 8075
rect 13596 8044 13737 8072
rect 13596 8032 13602 8044
rect 13725 8041 13737 8044
rect 13771 8041 13783 8075
rect 13725 8035 13783 8041
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14461 8075 14519 8081
rect 14461 8072 14473 8075
rect 14332 8044 14473 8072
rect 14332 8032 14338 8044
rect 14461 8041 14473 8044
rect 14507 8041 14519 8075
rect 22922 8072 22928 8084
rect 14461 8035 14519 8041
rect 17788 8044 22928 8072
rect 2130 7964 2136 8016
rect 2188 8004 2194 8016
rect 8478 8004 8484 8016
rect 2188 7976 8484 8004
rect 2188 7964 2194 7976
rect 8478 7964 8484 7976
rect 8536 7964 8542 8016
rect 11422 8004 11428 8016
rect 9876 7976 11428 8004
rect 7466 7896 7472 7948
rect 7524 7936 7530 7948
rect 7524 7908 8156 7936
rect 7524 7896 7530 7908
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 2832 7840 5549 7868
rect 2832 7828 2838 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5902 7828 5908 7880
rect 5960 7828 5966 7880
rect 6270 7828 6276 7880
rect 6328 7828 6334 7880
rect 6638 7828 6644 7880
rect 6696 7828 6702 7880
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 8128 7877 8156 7908
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6788 7840 7021 7868
rect 6788 7828 6794 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 4338 7760 4344 7812
rect 4396 7800 4402 7812
rect 7392 7800 7420 7831
rect 4396 7772 7420 7800
rect 8036 7800 8064 7831
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 9876 7877 9904 7976
rect 11422 7964 11428 7976
rect 11480 7964 11486 8016
rect 11882 8004 11888 8016
rect 11624 7976 11888 8004
rect 11514 7936 11520 7948
rect 10612 7908 11520 7936
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 8386 7800 8392 7812
rect 8036 7772 8392 7800
rect 4396 7760 4402 7772
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 9508 7800 9536 7831
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 10612 7877 10640 7908
rect 11514 7896 11520 7908
rect 11572 7896 11578 7948
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 10962 7828 10968 7880
rect 11020 7828 11026 7880
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7868 11391 7871
rect 11624 7868 11652 7976
rect 11882 7964 11888 7976
rect 11940 7964 11946 8016
rect 17788 8004 17816 8044
rect 22922 8032 22928 8044
rect 22980 8032 22986 8084
rect 25866 8032 25872 8084
rect 25924 8072 25930 8084
rect 26145 8075 26203 8081
rect 26145 8072 26157 8075
rect 25924 8044 26157 8072
rect 25924 8032 25930 8044
rect 26145 8041 26157 8044
rect 26191 8041 26203 8075
rect 26145 8035 26203 8041
rect 26326 8032 26332 8084
rect 26384 8072 26390 8084
rect 26513 8075 26571 8081
rect 26513 8072 26525 8075
rect 26384 8044 26525 8072
rect 26384 8032 26390 8044
rect 26513 8041 26525 8044
rect 26559 8041 26571 8075
rect 26513 8035 26571 8041
rect 26602 8032 26608 8084
rect 26660 8072 26666 8084
rect 26789 8075 26847 8081
rect 26789 8072 26801 8075
rect 26660 8044 26801 8072
rect 26660 8032 26666 8044
rect 26789 8041 26801 8044
rect 26835 8041 26847 8075
rect 26789 8035 26847 8041
rect 26878 8032 26884 8084
rect 26936 8072 26942 8084
rect 27157 8075 27215 8081
rect 27157 8072 27169 8075
rect 26936 8044 27169 8072
rect 26936 8032 26942 8044
rect 27157 8041 27169 8044
rect 27203 8041 27215 8075
rect 27157 8035 27215 8041
rect 27430 8032 27436 8084
rect 27488 8072 27494 8084
rect 27525 8075 27583 8081
rect 27525 8072 27537 8075
rect 27488 8044 27537 8072
rect 27488 8032 27494 8044
rect 27525 8041 27537 8044
rect 27571 8041 27583 8075
rect 27525 8035 27583 8041
rect 27706 8032 27712 8084
rect 27764 8072 27770 8084
rect 27985 8075 28043 8081
rect 27985 8072 27997 8075
rect 27764 8044 27997 8072
rect 27764 8032 27770 8044
rect 27985 8041 27997 8044
rect 28031 8041 28043 8075
rect 27985 8035 28043 8041
rect 28074 8032 28080 8084
rect 28132 8072 28138 8084
rect 28261 8075 28319 8081
rect 28261 8072 28273 8075
rect 28132 8044 28273 8072
rect 28132 8032 28138 8044
rect 28261 8041 28273 8044
rect 28307 8041 28319 8075
rect 28261 8035 28319 8041
rect 28350 8032 28356 8084
rect 28408 8072 28414 8084
rect 28629 8075 28687 8081
rect 28629 8072 28641 8075
rect 28408 8044 28641 8072
rect 28408 8032 28414 8044
rect 28629 8041 28641 8044
rect 28675 8041 28687 8075
rect 28629 8035 28687 8041
rect 31754 8032 31760 8084
rect 31812 8032 31818 8084
rect 32125 8075 32183 8081
rect 32125 8041 32137 8075
rect 32171 8072 32183 8075
rect 33410 8072 33416 8084
rect 32171 8044 33416 8072
rect 32171 8041 32183 8044
rect 32125 8035 32183 8041
rect 33410 8032 33416 8044
rect 33468 8032 33474 8084
rect 13556 7976 17816 8004
rect 11379 7840 11652 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 11698 7828 11704 7880
rect 11756 7828 11762 7880
rect 11790 7828 11796 7880
rect 11848 7828 11854 7880
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7837 12495 7871
rect 12437 7831 12495 7837
rect 10042 7800 10048 7812
rect 9508 7772 10048 7800
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 12452 7800 12480 7831
rect 12802 7828 12808 7880
rect 12860 7828 12866 7880
rect 13170 7828 13176 7880
rect 13228 7828 13234 7880
rect 13556 7877 13584 7976
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 17920 7976 31754 8004
rect 17920 7964 17926 7976
rect 18506 7896 18512 7948
rect 18564 7936 18570 7948
rect 31726 7936 31754 7976
rect 32398 7936 32404 7948
rect 18564 7908 31616 7936
rect 31726 7908 32404 7936
rect 18564 7896 18570 7908
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7837 13967 7871
rect 13909 7831 13967 7837
rect 13354 7800 13360 7812
rect 12452 7772 13360 7800
rect 13354 7760 13360 7772
rect 13412 7760 13418 7812
rect 13924 7800 13952 7831
rect 14642 7828 14648 7880
rect 14700 7828 14706 7880
rect 25314 7828 25320 7880
rect 25372 7868 25378 7880
rect 25961 7871 26019 7877
rect 25961 7868 25973 7871
rect 25372 7840 25973 7868
rect 25372 7828 25378 7840
rect 25961 7837 25973 7840
rect 26007 7837 26019 7871
rect 25961 7831 26019 7837
rect 26329 7871 26387 7877
rect 26329 7837 26341 7871
rect 26375 7837 26387 7871
rect 26329 7831 26387 7837
rect 26973 7871 27031 7877
rect 26973 7837 26985 7871
rect 27019 7837 27031 7871
rect 26973 7831 27031 7837
rect 27341 7871 27399 7877
rect 27341 7837 27353 7871
rect 27387 7868 27399 7871
rect 27614 7868 27620 7880
rect 27387 7840 27620 7868
rect 27387 7837 27399 7840
rect 27341 7831 27399 7837
rect 20346 7800 20352 7812
rect 13924 7772 20352 7800
rect 20346 7760 20352 7772
rect 20404 7760 20410 7812
rect 24854 7760 24860 7812
rect 24912 7800 24918 7812
rect 26344 7800 26372 7831
rect 24912 7772 26372 7800
rect 26988 7800 27016 7831
rect 27614 7828 27620 7840
rect 27672 7828 27678 7880
rect 27706 7828 27712 7880
rect 27764 7828 27770 7880
rect 27798 7828 27804 7880
rect 27856 7828 27862 7880
rect 28445 7871 28503 7877
rect 28445 7837 28457 7871
rect 28491 7837 28503 7871
rect 28445 7831 28503 7837
rect 28350 7800 28356 7812
rect 26988 7772 28356 7800
rect 24912 7760 24918 7772
rect 28350 7760 28356 7772
rect 28408 7760 28414 7812
rect 28460 7800 28488 7831
rect 28810 7828 28816 7880
rect 28868 7828 28874 7880
rect 29181 7871 29239 7877
rect 29181 7837 29193 7871
rect 29227 7868 29239 7871
rect 30650 7868 30656 7880
rect 29227 7840 30656 7868
rect 29227 7837 29239 7840
rect 29181 7831 29239 7837
rect 30650 7828 30656 7840
rect 30708 7828 30714 7880
rect 31588 7877 31616 7908
rect 32398 7896 32404 7908
rect 32456 7896 32462 7948
rect 31573 7871 31631 7877
rect 31573 7837 31585 7871
rect 31619 7837 31631 7871
rect 31573 7831 31631 7837
rect 31662 7828 31668 7880
rect 31720 7868 31726 7880
rect 31941 7871 31999 7877
rect 31941 7868 31953 7871
rect 31720 7840 31953 7868
rect 31720 7828 31726 7840
rect 31941 7837 31953 7840
rect 31987 7837 31999 7871
rect 31941 7831 31999 7837
rect 32306 7828 32312 7880
rect 32364 7828 32370 7880
rect 32674 7828 32680 7880
rect 32732 7828 32738 7880
rect 29086 7800 29092 7812
rect 28460 7772 29092 7800
rect 29086 7760 29092 7772
rect 29144 7760 29150 7812
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 10594 7732 10600 7744
rect 2556 7704 10600 7732
rect 2556 7692 2562 7704
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 12526 7732 12532 7744
rect 11020 7704 12532 7732
rect 11020 7692 11026 7704
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 20254 7732 20260 7744
rect 16908 7704 20260 7732
rect 16908 7692 16914 7704
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 22186 7692 22192 7744
rect 22244 7732 22250 7744
rect 26694 7732 26700 7744
rect 22244 7704 26700 7732
rect 22244 7692 22250 7704
rect 26694 7692 26700 7704
rect 26752 7692 26758 7744
rect 28442 7692 28448 7744
rect 28500 7732 28506 7744
rect 28997 7735 29055 7741
rect 28997 7732 29009 7735
rect 28500 7704 29009 7732
rect 28500 7692 28506 7704
rect 28997 7701 29009 7704
rect 29043 7701 29055 7735
rect 28997 7695 29055 7701
rect 32490 7692 32496 7744
rect 32548 7692 32554 7744
rect 32861 7735 32919 7741
rect 32861 7701 32873 7735
rect 32907 7732 32919 7735
rect 33594 7732 33600 7744
rect 32907 7704 33600 7732
rect 32907 7701 32919 7704
rect 32861 7695 32919 7701
rect 33594 7692 33600 7704
rect 33652 7692 33658 7744
rect 1104 7642 33324 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 33324 7642
rect 1104 7568 33324 7590
rect 2498 7488 2504 7540
rect 2556 7488 2562 7540
rect 2774 7488 2780 7540
rect 2832 7488 2838 7540
rect 3329 7531 3387 7537
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 5902 7528 5908 7540
rect 3375 7500 5908 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7377 7531 7435 7537
rect 7377 7528 7389 7531
rect 7156 7500 7389 7528
rect 7156 7488 7162 7500
rect 7377 7497 7389 7500
rect 7423 7497 7435 7531
rect 7377 7491 7435 7497
rect 9398 7488 9404 7540
rect 9456 7488 9462 7540
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 9732 7500 9873 7528
rect 9732 7488 9738 7500
rect 9861 7497 9873 7500
rect 9907 7497 9919 7531
rect 11146 7528 11152 7540
rect 9861 7491 9919 7497
rect 10980 7500 11152 7528
rect 10980 7460 11008 7500
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 11333 7531 11391 7537
rect 11333 7497 11345 7531
rect 11379 7528 11391 7531
rect 11790 7528 11796 7540
rect 11379 7500 11796 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 11977 7531 12035 7537
rect 11977 7528 11989 7531
rect 11940 7500 11989 7528
rect 11940 7488 11946 7500
rect 11977 7497 11989 7500
rect 12023 7497 12035 7531
rect 12253 7531 12311 7537
rect 12253 7528 12265 7531
rect 11977 7491 12035 7497
rect 12084 7500 12265 7528
rect 2884 7432 11008 7460
rect 2130 7352 2136 7404
rect 2188 7352 2194 7404
rect 2884 7401 2912 7432
rect 11054 7420 11060 7472
rect 11112 7460 11118 7472
rect 12084 7460 12112 7500
rect 12253 7497 12265 7500
rect 12299 7497 12311 7531
rect 12253 7491 12311 7497
rect 12526 7488 12532 7540
rect 12584 7488 12590 7540
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 12805 7531 12863 7537
rect 12805 7528 12817 7531
rect 12768 7500 12817 7528
rect 12768 7488 12774 7500
rect 12805 7497 12817 7500
rect 12851 7497 12863 7531
rect 12805 7491 12863 7497
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 16298 7528 16304 7540
rect 13412 7500 16304 7528
rect 13412 7488 13418 7500
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 16390 7488 16396 7540
rect 16448 7488 16454 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16632 7500 17049 7528
rect 16632 7488 16638 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 17405 7531 17463 7537
rect 17405 7497 17417 7531
rect 17451 7528 17463 7531
rect 17862 7528 17868 7540
rect 17451 7500 17868 7528
rect 17451 7497 17463 7500
rect 17405 7491 17463 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18506 7488 18512 7540
rect 18564 7488 18570 7540
rect 18785 7531 18843 7537
rect 18785 7497 18797 7531
rect 18831 7497 18843 7531
rect 18785 7491 18843 7497
rect 16666 7460 16672 7472
rect 11112 7432 12112 7460
rect 12268 7432 12572 7460
rect 11112 7420 11118 7432
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2547 7364 2605 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 4028 7364 7205 7392
rect 4028 7352 4034 7364
rect 7193 7361 7205 7364
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 9214 7352 9220 7404
rect 9272 7352 9278 7404
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7392 10103 7395
rect 10962 7392 10968 7404
rect 10091 7364 10968 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11146 7352 11152 7404
rect 11204 7352 11210 7404
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 12169 7395 12227 7401
rect 12169 7361 12181 7395
rect 12215 7392 12227 7395
rect 12268 7392 12296 7432
rect 12544 7404 12572 7432
rect 12728 7432 16672 7460
rect 12215 7364 12296 7392
rect 12437 7395 12495 7401
rect 12215 7361 12227 7364
rect 12169 7355 12227 7361
rect 12437 7361 12449 7395
rect 12483 7361 12495 7395
rect 12437 7355 12495 7361
rect 4798 7324 4804 7336
rect 2746 7296 4804 7324
rect 2317 7259 2375 7265
rect 2317 7225 2329 7259
rect 2363 7256 2375 7259
rect 2746 7256 2774 7296
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 2363 7228 2774 7256
rect 3053 7259 3111 7265
rect 2363 7225 2375 7228
rect 2317 7219 2375 7225
rect 3053 7225 3065 7259
rect 3099 7256 3111 7259
rect 5166 7256 5172 7268
rect 3099 7228 5172 7256
rect 3099 7225 3111 7228
rect 3053 7219 3111 7225
rect 5166 7216 5172 7228
rect 5224 7216 5230 7268
rect 10226 7216 10232 7268
rect 10284 7256 10290 7268
rect 11054 7256 11060 7268
rect 10284 7228 11060 7256
rect 10284 7216 10290 7228
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 11238 7216 11244 7268
rect 11296 7256 11302 7268
rect 11701 7259 11759 7265
rect 11701 7256 11713 7259
rect 11296 7228 11713 7256
rect 11296 7216 11302 7228
rect 11701 7225 11713 7228
rect 11747 7225 11759 7259
rect 11900 7256 11928 7355
rect 12452 7324 12480 7355
rect 12526 7352 12532 7404
rect 12584 7352 12590 7404
rect 12728 7401 12756 7432
rect 16666 7420 16672 7432
rect 16724 7420 16730 7472
rect 18800 7460 18828 7491
rect 19518 7488 19524 7540
rect 19576 7488 19582 7540
rect 19794 7488 19800 7540
rect 19852 7488 19858 7540
rect 20714 7488 20720 7540
rect 20772 7488 20778 7540
rect 21085 7531 21143 7537
rect 21085 7497 21097 7531
rect 21131 7528 21143 7531
rect 21266 7528 21272 7540
rect 21131 7500 21272 7528
rect 21131 7497 21143 7500
rect 21085 7491 21143 7497
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 21361 7531 21419 7537
rect 21361 7497 21373 7531
rect 21407 7497 21419 7531
rect 21361 7491 21419 7497
rect 21376 7460 21404 7491
rect 21542 7488 21548 7540
rect 21600 7528 21606 7540
rect 25222 7528 25228 7540
rect 21600 7500 25228 7528
rect 21600 7488 21606 7500
rect 25222 7488 25228 7500
rect 25280 7488 25286 7540
rect 27798 7488 27804 7540
rect 27856 7488 27862 7540
rect 28537 7531 28595 7537
rect 28537 7497 28549 7531
rect 28583 7528 28595 7531
rect 28718 7528 28724 7540
rect 28583 7500 28724 7528
rect 28583 7497 28595 7500
rect 28537 7491 28595 7497
rect 28718 7488 28724 7500
rect 28776 7488 28782 7540
rect 28902 7488 28908 7540
rect 28960 7488 28966 7540
rect 29086 7488 29092 7540
rect 29144 7528 29150 7540
rect 29181 7531 29239 7537
rect 29181 7528 29193 7531
rect 29144 7500 29193 7528
rect 29144 7488 29150 7500
rect 29181 7497 29193 7500
rect 29227 7497 29239 7531
rect 29181 7491 29239 7497
rect 29733 7531 29791 7537
rect 29733 7497 29745 7531
rect 29779 7528 29791 7531
rect 29822 7528 29828 7540
rect 29779 7500 29828 7528
rect 29779 7497 29791 7500
rect 29733 7491 29791 7497
rect 29822 7488 29828 7500
rect 29880 7488 29886 7540
rect 30650 7488 30656 7540
rect 30708 7488 30714 7540
rect 32493 7531 32551 7537
rect 32493 7497 32505 7531
rect 32539 7528 32551 7531
rect 32582 7528 32588 7540
rect 32539 7500 32588 7528
rect 32539 7497 32551 7500
rect 32493 7491 32551 7497
rect 32582 7488 32588 7500
rect 32640 7488 32646 7540
rect 32766 7460 32772 7472
rect 18800 7432 21312 7460
rect 21376 7432 28948 7460
rect 12713 7395 12771 7401
rect 12713 7361 12725 7395
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7392 13047 7395
rect 16206 7392 16212 7404
rect 13035 7364 16212 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7392 16543 7395
rect 16761 7395 16819 7401
rect 16761 7392 16773 7395
rect 16531 7364 16773 7392
rect 16531 7361 16543 7364
rect 16485 7355 16543 7361
rect 16761 7361 16773 7364
rect 16807 7361 16819 7395
rect 16761 7355 16819 7361
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 17175 7364 17233 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7392 18291 7395
rect 18325 7395 18383 7401
rect 18325 7392 18337 7395
rect 18279 7364 18337 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 18325 7361 18337 7364
rect 18371 7361 18383 7395
rect 18325 7355 18383 7361
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 18656 7364 18889 7392
rect 18656 7352 18662 7364
rect 18877 7361 18889 7364
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 19245 7395 19303 7401
rect 19245 7361 19257 7395
rect 19291 7392 19303 7395
rect 19337 7395 19395 7401
rect 19337 7392 19349 7395
rect 19291 7364 19349 7392
rect 19291 7361 19303 7364
rect 19245 7355 19303 7361
rect 19337 7361 19349 7364
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 19610 7352 19616 7404
rect 19668 7352 19674 7404
rect 19702 7352 19708 7404
rect 19760 7392 19766 7404
rect 19981 7395 20039 7401
rect 19981 7392 19993 7395
rect 19760 7364 19993 7392
rect 19760 7352 19766 7364
rect 19981 7361 19993 7364
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 20438 7352 20444 7404
rect 20496 7352 20502 7404
rect 20809 7395 20867 7401
rect 20809 7361 20821 7395
rect 20855 7392 20867 7395
rect 20901 7395 20959 7401
rect 20901 7392 20913 7395
rect 20855 7364 20913 7392
rect 20855 7361 20867 7364
rect 20809 7355 20867 7361
rect 20901 7361 20913 7364
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 21174 7352 21180 7404
rect 21232 7352 21238 7404
rect 21284 7392 21312 7432
rect 24762 7392 24768 7404
rect 21284 7364 24768 7392
rect 24762 7352 24768 7364
rect 24820 7352 24826 7404
rect 24946 7352 24952 7404
rect 25004 7392 25010 7404
rect 27985 7395 28043 7401
rect 27985 7392 27997 7395
rect 25004 7364 27997 7392
rect 25004 7352 25010 7364
rect 27985 7361 27997 7364
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 28074 7352 28080 7404
rect 28132 7392 28138 7404
rect 28353 7395 28411 7401
rect 28353 7392 28365 7395
rect 28132 7364 28365 7392
rect 28132 7352 28138 7364
rect 28353 7361 28365 7364
rect 28399 7361 28411 7395
rect 28353 7355 28411 7361
rect 28442 7352 28448 7404
rect 28500 7392 28506 7404
rect 28813 7395 28871 7401
rect 28813 7392 28825 7395
rect 28500 7364 28825 7392
rect 28500 7352 28506 7364
rect 28813 7361 28825 7364
rect 28859 7361 28871 7395
rect 28813 7355 28871 7361
rect 12452 7296 12756 7324
rect 12434 7256 12440 7268
rect 11900 7228 12440 7256
rect 11701 7219 11759 7225
rect 12434 7216 12440 7228
rect 12492 7216 12498 7268
rect 12728 7256 12756 7296
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 19794 7324 19800 7336
rect 12860 7296 19800 7324
rect 12860 7284 12866 7296
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 26786 7324 26792 7336
rect 20180 7296 26792 7324
rect 16850 7256 16856 7268
rect 12728 7228 16856 7256
rect 16850 7216 16856 7228
rect 16908 7216 16914 7268
rect 16945 7259 17003 7265
rect 16945 7225 16957 7259
rect 16991 7256 17003 7259
rect 17954 7256 17960 7268
rect 16991 7228 17960 7256
rect 16991 7225 17003 7228
rect 16945 7219 17003 7225
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 18138 7216 18144 7268
rect 18196 7216 18202 7268
rect 20180 7265 20208 7296
rect 26786 7284 26792 7296
rect 26844 7284 26850 7336
rect 28920 7324 28948 7432
rect 29932 7432 32772 7460
rect 29086 7352 29092 7404
rect 29144 7352 29150 7404
rect 29362 7352 29368 7404
rect 29420 7352 29426 7404
rect 29932 7401 29960 7432
rect 32766 7420 32772 7432
rect 32824 7420 32830 7472
rect 29917 7395 29975 7401
rect 29917 7361 29929 7395
rect 29963 7361 29975 7395
rect 29917 7355 29975 7361
rect 30193 7395 30251 7401
rect 30193 7361 30205 7395
rect 30239 7361 30251 7395
rect 30193 7355 30251 7361
rect 30837 7395 30895 7401
rect 30837 7361 30849 7395
rect 30883 7392 30895 7395
rect 31202 7392 31208 7404
rect 30883 7364 31208 7392
rect 30883 7361 30895 7364
rect 30837 7355 30895 7361
rect 28736 7296 28948 7324
rect 20165 7259 20223 7265
rect 20165 7225 20177 7259
rect 20211 7225 20223 7259
rect 20165 7219 20223 7225
rect 20625 7259 20683 7265
rect 20625 7225 20637 7259
rect 20671 7256 20683 7259
rect 26878 7256 26884 7268
rect 20671 7228 26884 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 26878 7216 26884 7228
rect 26936 7216 26942 7268
rect 27706 7216 27712 7268
rect 27764 7256 27770 7268
rect 28629 7259 28687 7265
rect 28629 7256 28641 7259
rect 27764 7228 28641 7256
rect 27764 7216 27770 7228
rect 28629 7225 28641 7228
rect 28675 7225 28687 7259
rect 28629 7219 28687 7225
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 10870 7188 10876 7200
rect 3200 7160 10876 7188
rect 3200 7148 3206 7160
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 12342 7188 12348 7200
rect 11020 7160 12348 7188
rect 11020 7148 11026 7160
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 13262 7188 13268 7200
rect 12584 7160 13268 7188
rect 12584 7148 12590 7160
rect 13262 7148 13268 7160
rect 13320 7148 13326 7200
rect 17770 7148 17776 7200
rect 17828 7188 17834 7200
rect 19153 7191 19211 7197
rect 19153 7188 19165 7191
rect 17828 7160 19165 7188
rect 17828 7148 17834 7160
rect 19153 7157 19165 7160
rect 19199 7157 19211 7191
rect 19153 7151 19211 7157
rect 21174 7148 21180 7200
rect 21232 7188 21238 7200
rect 21453 7191 21511 7197
rect 21453 7188 21465 7191
rect 21232 7160 21465 7188
rect 21232 7148 21238 7160
rect 21453 7157 21465 7160
rect 21499 7157 21511 7191
rect 28736 7188 28764 7296
rect 29638 7284 29644 7336
rect 29696 7324 29702 7336
rect 30208 7324 30236 7355
rect 31202 7352 31208 7364
rect 31260 7352 31266 7404
rect 32309 7395 32367 7401
rect 32309 7392 32321 7395
rect 31726 7364 32321 7392
rect 29696 7296 30236 7324
rect 29696 7284 29702 7296
rect 28810 7216 28816 7268
rect 28868 7256 28874 7268
rect 30009 7259 30067 7265
rect 30009 7256 30021 7259
rect 28868 7228 30021 7256
rect 28868 7216 28874 7228
rect 30009 7225 30021 7228
rect 30055 7225 30067 7259
rect 31726 7256 31754 7364
rect 32309 7361 32321 7364
rect 32355 7361 32367 7395
rect 32309 7355 32367 7361
rect 32398 7352 32404 7404
rect 32456 7392 32462 7404
rect 32677 7395 32735 7401
rect 32677 7392 32689 7395
rect 32456 7364 32689 7392
rect 32456 7352 32462 7364
rect 32677 7361 32689 7364
rect 32723 7361 32735 7395
rect 32677 7355 32735 7361
rect 32674 7256 32680 7268
rect 30009 7219 30067 7225
rect 30116 7228 31754 7256
rect 32232 7228 32680 7256
rect 30116 7188 30144 7228
rect 28736 7160 30144 7188
rect 21453 7151 21511 7157
rect 30190 7148 30196 7200
rect 30248 7188 30254 7200
rect 32232 7188 32260 7228
rect 32674 7216 32680 7228
rect 32732 7216 32738 7268
rect 30248 7160 32260 7188
rect 30248 7148 30254 7160
rect 32858 7148 32864 7200
rect 32916 7148 32922 7200
rect 1104 7098 33304 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 33304 7098
rect 1104 7024 33304 7046
rect 3970 6944 3976 6996
rect 4028 6944 4034 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 11756 6956 12081 6984
rect 11756 6944 11762 6956
rect 12069 6953 12081 6956
rect 12115 6953 12127 6987
rect 12069 6947 12127 6953
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 15562 6984 15568 6996
rect 12492 6956 15568 6984
rect 12492 6944 12498 6956
rect 15562 6944 15568 6956
rect 15620 6944 15626 6996
rect 24578 6944 24584 6996
rect 24636 6984 24642 6996
rect 24636 6956 24992 6984
rect 24636 6944 24642 6956
rect 4430 6916 4436 6928
rect 3712 6888 4436 6916
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 3326 6780 3332 6792
rect 3191 6752 3332 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3712 6780 3740 6888
rect 4430 6876 4436 6888
rect 4488 6876 4494 6928
rect 11146 6876 11152 6928
rect 11204 6916 11210 6928
rect 19058 6916 19064 6928
rect 11204 6888 19064 6916
rect 11204 6876 11210 6888
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 23106 6876 23112 6928
rect 23164 6916 23170 6928
rect 23164 6888 24900 6916
rect 23164 6876 23170 6888
rect 6822 6848 6828 6860
rect 3804 6820 6828 6848
rect 3804 6789 3832 6820
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 9950 6848 9956 6860
rect 7116 6820 9956 6848
rect 3467 6752 3740 6780
rect 3789 6783 3847 6789
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6780 4123 6783
rect 6914 6780 6920 6792
rect 4111 6752 6920 6780
rect 4111 6749 4123 6752
rect 4065 6743 4123 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 4338 6712 4344 6724
rect 3344 6684 4344 6712
rect 3344 6653 3372 6684
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 4430 6672 4436 6724
rect 4488 6712 4494 6724
rect 7116 6712 7144 6820
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 12894 6848 12900 6860
rect 12406 6820 12900 6848
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12406 6780 12434 6820
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 17034 6848 17040 6860
rect 13044 6820 17040 6848
rect 13044 6808 13050 6820
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 23290 6808 23296 6860
rect 23348 6848 23354 6860
rect 23348 6820 24624 6848
rect 23348 6808 23354 6820
rect 12299 6752 12434 6780
rect 12529 6783 12587 6789
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 13630 6780 13636 6792
rect 12575 6752 13636 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 4488 6684 7144 6712
rect 7208 6712 7236 6743
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 14550 6740 14556 6792
rect 14608 6780 14614 6792
rect 21910 6780 21916 6792
rect 14608 6752 21916 6780
rect 14608 6740 14614 6752
rect 21910 6740 21916 6752
rect 21968 6740 21974 6792
rect 23474 6740 23480 6792
rect 23532 6780 23538 6792
rect 24596 6789 24624 6820
rect 24872 6789 24900 6888
rect 24964 6848 24992 6956
rect 26878 6944 26884 6996
rect 26936 6984 26942 6996
rect 32306 6984 32312 6996
rect 26936 6956 32312 6984
rect 26936 6944 26942 6956
rect 32306 6944 32312 6956
rect 32364 6944 32370 6996
rect 26786 6876 26792 6928
rect 26844 6916 26850 6928
rect 30190 6916 30196 6928
rect 26844 6888 30196 6916
rect 26844 6876 26850 6888
rect 30190 6876 30196 6888
rect 30248 6876 30254 6928
rect 24964 6820 26004 6848
rect 24121 6783 24179 6789
rect 24121 6780 24133 6783
rect 23532 6752 24133 6780
rect 23532 6740 23538 6752
rect 24121 6749 24133 6752
rect 24167 6749 24179 6783
rect 24121 6743 24179 6749
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6749 24639 6783
rect 24581 6743 24639 6749
rect 24857 6783 24915 6789
rect 24857 6749 24869 6783
rect 24903 6749 24915 6783
rect 24857 6743 24915 6749
rect 25130 6740 25136 6792
rect 25188 6740 25194 6792
rect 25590 6740 25596 6792
rect 25648 6740 25654 6792
rect 25976 6789 26004 6820
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6749 26019 6783
rect 25961 6743 26019 6749
rect 26326 6740 26332 6792
rect 26384 6740 26390 6792
rect 26694 6740 26700 6792
rect 26752 6740 26758 6792
rect 26970 6740 26976 6792
rect 27028 6740 27034 6792
rect 29270 6740 29276 6792
rect 29328 6740 29334 6792
rect 30650 6740 30656 6792
rect 30708 6780 30714 6792
rect 32309 6783 32367 6789
rect 32309 6780 32321 6783
rect 30708 6752 32321 6780
rect 30708 6740 30714 6752
rect 32309 6749 32321 6752
rect 32355 6749 32367 6783
rect 32309 6743 32367 6749
rect 32398 6740 32404 6792
rect 32456 6780 32462 6792
rect 32677 6783 32735 6789
rect 32677 6780 32689 6783
rect 32456 6752 32689 6780
rect 32456 6740 32462 6752
rect 32677 6749 32689 6752
rect 32723 6749 32735 6783
rect 32677 6743 32735 6749
rect 14826 6712 14832 6724
rect 7208 6684 14832 6712
rect 4488 6672 4494 6684
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 14918 6672 14924 6724
rect 14976 6712 14982 6724
rect 33410 6712 33416 6724
rect 14976 6684 26188 6712
rect 14976 6672 14982 6684
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6613 3387 6647
rect 3329 6607 3387 6613
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 4154 6644 4160 6656
rect 3651 6616 4160 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4249 6647 4307 6653
rect 4249 6613 4261 6647
rect 4295 6644 4307 6647
rect 6730 6644 6736 6656
rect 4295 6616 6736 6644
rect 4295 6613 4307 6616
rect 4249 6607 4307 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 7377 6647 7435 6653
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 9214 6644 9220 6656
rect 7423 6616 9220 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 11664 6616 12357 6644
rect 11664 6604 11670 6616
rect 12345 6613 12357 6616
rect 12391 6613 12403 6647
rect 12345 6607 12403 6613
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 17586 6644 17592 6656
rect 13228 6616 17592 6644
rect 13228 6604 13234 6616
rect 17586 6604 17592 6616
rect 17644 6604 17650 6656
rect 20346 6604 20352 6656
rect 20404 6644 20410 6656
rect 23937 6647 23995 6653
rect 23937 6644 23949 6647
rect 20404 6616 23949 6644
rect 20404 6604 20410 6616
rect 23937 6613 23949 6616
rect 23983 6613 23995 6647
rect 23937 6607 23995 6613
rect 24394 6604 24400 6656
rect 24452 6604 24458 6656
rect 24670 6604 24676 6656
rect 24728 6604 24734 6656
rect 24949 6647 25007 6653
rect 24949 6613 24961 6647
rect 24995 6644 25007 6647
rect 25038 6644 25044 6656
rect 24995 6616 25044 6644
rect 24995 6613 25007 6616
rect 24949 6607 25007 6613
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 25406 6604 25412 6656
rect 25464 6604 25470 6656
rect 25498 6604 25504 6656
rect 25556 6644 25562 6656
rect 26160 6653 26188 6684
rect 32508 6684 33416 6712
rect 25777 6647 25835 6653
rect 25777 6644 25789 6647
rect 25556 6616 25789 6644
rect 25556 6604 25562 6616
rect 25777 6613 25789 6616
rect 25823 6613 25835 6647
rect 25777 6607 25835 6613
rect 26145 6647 26203 6653
rect 26145 6613 26157 6647
rect 26191 6613 26203 6647
rect 26145 6607 26203 6613
rect 26418 6604 26424 6656
rect 26476 6644 26482 6656
rect 26513 6647 26571 6653
rect 26513 6644 26525 6647
rect 26476 6616 26525 6644
rect 26476 6604 26482 6616
rect 26513 6613 26525 6616
rect 26559 6613 26571 6647
rect 26513 6607 26571 6613
rect 26602 6604 26608 6656
rect 26660 6644 26666 6656
rect 26789 6647 26847 6653
rect 26789 6644 26801 6647
rect 26660 6616 26801 6644
rect 26660 6604 26666 6616
rect 26789 6613 26801 6616
rect 26835 6613 26847 6647
rect 26789 6607 26847 6613
rect 28626 6604 28632 6656
rect 28684 6644 28690 6656
rect 32508 6653 32536 6684
rect 33410 6672 33416 6684
rect 33468 6672 33474 6724
rect 29089 6647 29147 6653
rect 29089 6644 29101 6647
rect 28684 6616 29101 6644
rect 28684 6604 28690 6616
rect 29089 6613 29101 6616
rect 29135 6613 29147 6647
rect 29089 6607 29147 6613
rect 32493 6647 32551 6653
rect 32493 6613 32505 6647
rect 32539 6613 32551 6647
rect 32493 6607 32551 6613
rect 32858 6604 32864 6656
rect 32916 6604 32922 6656
rect 1104 6554 33324 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 33324 6554
rect 1104 6480 33324 6502
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4890 6440 4896 6452
rect 4019 6412 4896 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5258 6440 5264 6452
rect 5031 6412 5264 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6512 6412 6745 6440
rect 6512 6400 6518 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 6917 6443 6975 6449
rect 6917 6409 6929 6443
rect 6963 6440 6975 6443
rect 7098 6440 7104 6452
rect 6963 6412 7104 6440
rect 6963 6409 6975 6412
rect 6917 6403 6975 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 7190 6400 7196 6452
rect 7248 6400 7254 6452
rect 7466 6400 7472 6452
rect 7524 6400 7530 6452
rect 7558 6400 7564 6452
rect 7616 6400 7622 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 7800 6412 8125 6440
rect 7800 6400 7806 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 8113 6403 8171 6409
rect 8386 6400 8392 6452
rect 8444 6400 8450 6452
rect 13722 6400 13728 6452
rect 13780 6400 13786 6452
rect 14458 6400 14464 6452
rect 14516 6440 14522 6452
rect 15105 6443 15163 6449
rect 15105 6440 15117 6443
rect 14516 6412 15117 6440
rect 14516 6400 14522 6412
rect 15105 6409 15117 6412
rect 15151 6409 15163 6443
rect 15105 6403 15163 6409
rect 15194 6400 15200 6452
rect 15252 6440 15258 6452
rect 17494 6440 17500 6452
rect 15252 6412 17500 6440
rect 15252 6400 15258 6412
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 17586 6400 17592 6452
rect 17644 6440 17650 6452
rect 22649 6443 22707 6449
rect 22649 6440 22661 6443
rect 17644 6412 22661 6440
rect 17644 6400 17650 6412
rect 22649 6409 22661 6412
rect 22695 6409 22707 6443
rect 24210 6440 24216 6452
rect 22649 6403 22707 6409
rect 22848 6412 24216 6440
rect 12986 6372 12992 6384
rect 6472 6344 12992 6372
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6304 4031 6307
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 4019 6276 4077 6304
rect 4019 6273 4031 6276
rect 3973 6267 4031 6273
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4522 6264 4528 6316
rect 4580 6264 4586 6316
rect 4798 6264 4804 6316
rect 4856 6264 4862 6316
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 6472 6304 6500 6344
rect 12986 6332 12992 6344
rect 13044 6332 13050 6384
rect 13265 6375 13323 6381
rect 13265 6341 13277 6375
rect 13311 6372 13323 6375
rect 15473 6375 15531 6381
rect 15473 6372 15485 6375
rect 13311 6344 13676 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 5123 6276 6500 6304
rect 6549 6307 6607 6313
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 7009 6307 7067 6313
rect 6595 6276 6960 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 6638 6236 6644 6248
rect 4264 6208 6644 6236
rect 4264 6177 4292 6208
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 4249 6171 4307 6177
rect 4249 6137 4261 6171
rect 4295 6137 4307 6171
rect 4249 6131 4307 6137
rect 5261 6171 5319 6177
rect 5261 6137 5273 6171
rect 5307 6168 5319 6171
rect 5442 6168 5448 6180
rect 5307 6140 5448 6168
rect 5307 6137 5319 6140
rect 5261 6131 5319 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 4709 6103 4767 6109
rect 4709 6069 4721 6103
rect 4755 6100 4767 6103
rect 6270 6100 6276 6112
rect 4755 6072 6276 6100
rect 4755 6069 4767 6072
rect 4709 6063 4767 6069
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 6932 6100 6960 6276
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7190 6304 7196 6316
rect 7055 6276 7196 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7300 6168 7328 6267
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 9582 6304 9588 6316
rect 8619 6276 9588 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6236 8079 6239
rect 8312 6236 8340 6267
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6304 13139 6307
rect 13541 6307 13599 6313
rect 13541 6304 13553 6307
rect 13127 6276 13553 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 13541 6273 13553 6276
rect 13587 6273 13599 6307
rect 13648 6304 13676 6344
rect 14660 6344 15485 6372
rect 13817 6307 13875 6313
rect 13817 6304 13829 6307
rect 13648 6276 13829 6304
rect 13541 6267 13599 6273
rect 13817 6273 13829 6276
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13964 6276 14105 6304
rect 13964 6264 13970 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 12158 6236 12164 6248
rect 8067 6208 12164 6236
rect 8067 6205 8079 6208
rect 8021 6199 8079 6205
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 12897 6239 12955 6245
rect 12897 6205 12909 6239
rect 12943 6236 12955 6239
rect 13449 6239 13507 6245
rect 12943 6208 13400 6236
rect 12943 6205 12955 6208
rect 12897 6199 12955 6205
rect 8294 6168 8300 6180
rect 7300 6140 8300 6168
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 13372 6168 13400 6208
rect 13449 6205 13461 6239
rect 13495 6236 13507 6239
rect 14384 6236 14412 6267
rect 14550 6264 14556 6316
rect 14608 6304 14614 6316
rect 14660 6313 14688 6344
rect 15473 6341 15485 6344
rect 15519 6341 15531 6375
rect 15473 6335 15531 6341
rect 16574 6332 16580 6384
rect 16632 6372 16638 6384
rect 17218 6372 17224 6384
rect 16632 6344 17224 6372
rect 16632 6332 16638 6344
rect 17218 6332 17224 6344
rect 17276 6332 17282 6384
rect 21652 6344 22508 6372
rect 21652 6313 21680 6344
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 14608 6276 14657 6304
rect 14608 6264 14614 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14645 6267 14703 6273
rect 14844 6276 14933 6304
rect 13495 6208 14412 6236
rect 14844 6236 14872 6276
rect 14921 6273 14933 6276
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6304 15255 6307
rect 15657 6307 15715 6313
rect 15657 6304 15669 6307
rect 15243 6276 15669 6304
rect 15243 6273 15255 6276
rect 15197 6267 15255 6273
rect 15657 6273 15669 6276
rect 15703 6273 15715 6307
rect 15657 6267 15715 6273
rect 21637 6307 21695 6313
rect 21637 6273 21649 6307
rect 21683 6273 21695 6307
rect 21637 6267 21695 6273
rect 21910 6264 21916 6316
rect 21968 6264 21974 6316
rect 22002 6264 22008 6316
rect 22060 6313 22066 6316
rect 22060 6267 22071 6313
rect 22060 6264 22066 6267
rect 22278 6264 22284 6316
rect 22336 6264 22342 6316
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 14844 6208 15853 6236
rect 13495 6205 13507 6208
rect 13449 6199 13507 6205
rect 13372 6140 13584 6168
rect 11974 6100 11980 6112
rect 6932 6072 11980 6100
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12802 6060 12808 6112
rect 12860 6060 12866 6112
rect 12986 6060 12992 6112
rect 13044 6060 13050 6112
rect 13170 6060 13176 6112
rect 13228 6060 13234 6112
rect 13354 6060 13360 6112
rect 13412 6060 13418 6112
rect 13556 6100 13584 6140
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 14844 6168 14872 6208
rect 15841 6205 15853 6208
rect 15887 6205 15899 6239
rect 15841 6199 15899 6205
rect 16298 6196 16304 6248
rect 16356 6236 16362 6248
rect 21928 6236 21956 6264
rect 16356 6208 21864 6236
rect 21928 6208 22416 6236
rect 16356 6196 16362 6208
rect 13688 6140 14872 6168
rect 15381 6171 15439 6177
rect 13688 6128 13694 6140
rect 15381 6137 15393 6171
rect 15427 6168 15439 6171
rect 16022 6168 16028 6180
rect 15427 6140 16028 6168
rect 15427 6137 15439 6140
rect 15381 6131 15439 6137
rect 16022 6128 16028 6140
rect 16080 6128 16086 6180
rect 19794 6128 19800 6180
rect 19852 6168 19858 6180
rect 21836 6168 21864 6208
rect 22388 6177 22416 6208
rect 22097 6171 22155 6177
rect 22097 6168 22109 6171
rect 19852 6140 21588 6168
rect 21836 6140 22109 6168
rect 19852 6128 19858 6140
rect 13906 6100 13912 6112
rect 13556 6072 13912 6100
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 13998 6060 14004 6112
rect 14056 6060 14062 6112
rect 14277 6103 14335 6109
rect 14277 6069 14289 6103
rect 14323 6100 14335 6103
rect 14366 6100 14372 6112
rect 14323 6072 14372 6100
rect 14323 6069 14335 6072
rect 14277 6063 14335 6069
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 14553 6103 14611 6109
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 14734 6100 14740 6112
rect 14599 6072 14740 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 14734 6060 14740 6072
rect 14792 6060 14798 6112
rect 14829 6103 14887 6109
rect 14829 6069 14841 6103
rect 14875 6100 14887 6103
rect 14918 6100 14924 6112
rect 14875 6072 14924 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 15654 6060 15660 6112
rect 15712 6060 15718 6112
rect 17954 6060 17960 6112
rect 18012 6100 18018 6112
rect 19426 6100 19432 6112
rect 18012 6072 19432 6100
rect 18012 6060 18018 6072
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 20898 6060 20904 6112
rect 20956 6100 20962 6112
rect 21453 6103 21511 6109
rect 21453 6100 21465 6103
rect 20956 6072 21465 6100
rect 20956 6060 20962 6072
rect 21453 6069 21465 6072
rect 21499 6069 21511 6103
rect 21560 6100 21588 6140
rect 22097 6137 22109 6140
rect 22143 6137 22155 6171
rect 22097 6131 22155 6137
rect 22373 6171 22431 6177
rect 22373 6137 22385 6171
rect 22419 6137 22431 6171
rect 22373 6131 22431 6137
rect 21821 6103 21879 6109
rect 21821 6100 21833 6103
rect 21560 6072 21833 6100
rect 21453 6063 21511 6069
rect 21821 6069 21833 6072
rect 21867 6069 21879 6103
rect 22480 6100 22508 6344
rect 22848 6313 22876 6412
rect 24210 6400 24216 6412
rect 24268 6400 24274 6452
rect 24486 6400 24492 6452
rect 24544 6440 24550 6452
rect 26418 6440 26424 6452
rect 24544 6412 26424 6440
rect 24544 6400 24550 6412
rect 26418 6400 26424 6412
rect 26476 6400 26482 6452
rect 32858 6400 32864 6452
rect 32916 6400 32922 6452
rect 23842 6372 23848 6384
rect 23124 6344 23848 6372
rect 23124 6313 23152 6344
rect 23842 6332 23848 6344
rect 23900 6332 23906 6384
rect 22557 6307 22615 6313
rect 22557 6273 22569 6307
rect 22603 6273 22615 6307
rect 22557 6267 22615 6273
rect 22833 6307 22891 6313
rect 22833 6273 22845 6307
rect 22879 6273 22891 6307
rect 22833 6267 22891 6273
rect 23109 6307 23167 6313
rect 23109 6273 23121 6307
rect 23155 6273 23167 6307
rect 23109 6267 23167 6273
rect 23385 6307 23443 6313
rect 23385 6273 23397 6307
rect 23431 6304 23443 6307
rect 23658 6304 23664 6316
rect 23431 6276 23664 6304
rect 23431 6273 23443 6276
rect 23385 6267 23443 6273
rect 22572 6236 22600 6267
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 32306 6264 32312 6316
rect 32364 6264 32370 6316
rect 32677 6307 32735 6313
rect 32677 6273 32689 6307
rect 32723 6273 32735 6307
rect 32677 6267 32735 6273
rect 24026 6236 24032 6248
rect 22572 6208 24032 6236
rect 24026 6196 24032 6208
rect 24084 6196 24090 6248
rect 30466 6196 30472 6248
rect 30524 6236 30530 6248
rect 32692 6236 32720 6267
rect 30524 6208 32720 6236
rect 30524 6196 30530 6208
rect 22922 6128 22928 6180
rect 22980 6128 22986 6180
rect 24302 6168 24308 6180
rect 23124 6140 24308 6168
rect 23124 6100 23152 6140
rect 24302 6128 24308 6140
rect 24360 6128 24366 6180
rect 22480 6072 23152 6100
rect 21821 6063 21879 6069
rect 23198 6060 23204 6112
rect 23256 6060 23262 6112
rect 32490 6060 32496 6112
rect 32548 6060 32554 6112
rect 1104 6010 33304 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 33304 6010
rect 1104 5936 33304 5958
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 7374 5896 7380 5908
rect 4856 5868 7380 5896
rect 4856 5856 4862 5868
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7469 5899 7527 5905
rect 7469 5865 7481 5899
rect 7515 5896 7527 5899
rect 8478 5896 8484 5908
rect 7515 5868 8484 5896
rect 7515 5865 7527 5868
rect 7469 5859 7527 5865
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 12710 5896 12716 5908
rect 8588 5868 12716 5896
rect 4522 5788 4528 5840
rect 4580 5828 4586 5840
rect 8588 5828 8616 5868
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 17954 5896 17960 5908
rect 12952 5868 17960 5896
rect 12952 5856 12958 5868
rect 17954 5856 17960 5868
rect 18012 5856 18018 5908
rect 18046 5856 18052 5908
rect 18104 5896 18110 5908
rect 23198 5896 23204 5908
rect 18104 5868 23204 5896
rect 18104 5856 18110 5868
rect 23198 5856 23204 5868
rect 23256 5856 23262 5908
rect 32306 5896 32312 5908
rect 31726 5868 32312 5896
rect 4580 5800 8616 5828
rect 4580 5788 4586 5800
rect 10962 5788 10968 5840
rect 11020 5828 11026 5840
rect 13354 5828 13360 5840
rect 11020 5800 13360 5828
rect 11020 5788 11026 5800
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 16482 5828 16488 5840
rect 14568 5800 16488 5828
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 6972 5732 12434 5760
rect 6972 5720 6978 5732
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 7064 5664 7297 5692
rect 7064 5652 7070 5664
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 12406 5692 12434 5732
rect 14568 5692 14596 5800
rect 16482 5788 16488 5800
rect 16540 5788 16546 5840
rect 17313 5831 17371 5837
rect 17313 5797 17325 5831
rect 17359 5828 17371 5831
rect 19702 5828 19708 5840
rect 17359 5800 19708 5828
rect 17359 5797 17371 5800
rect 17313 5791 17371 5797
rect 19702 5788 19708 5800
rect 19760 5788 19766 5840
rect 20346 5788 20352 5840
rect 20404 5828 20410 5840
rect 31726 5828 31754 5868
rect 32306 5856 32312 5868
rect 32364 5856 32370 5908
rect 20404 5800 31754 5828
rect 20404 5788 20410 5800
rect 32858 5788 32864 5840
rect 32916 5788 32922 5840
rect 14642 5720 14648 5772
rect 14700 5760 14706 5772
rect 25406 5760 25412 5772
rect 14700 5732 25412 5760
rect 14700 5720 14706 5732
rect 25406 5720 25412 5732
rect 25464 5720 25470 5772
rect 32398 5760 32404 5772
rect 27356 5732 32404 5760
rect 12406 5664 14596 5692
rect 15565 5695 15623 5701
rect 7285 5655 7343 5661
rect 15565 5661 15577 5695
rect 15611 5692 15623 5695
rect 15657 5695 15715 5701
rect 15657 5692 15669 5695
rect 15611 5664 15669 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 15657 5661 15669 5664
rect 15703 5661 15715 5695
rect 16574 5692 16580 5704
rect 15657 5655 15715 5661
rect 16408 5664 16580 5692
rect 3418 5584 3424 5636
rect 3476 5624 3482 5636
rect 10686 5624 10692 5636
rect 3476 5596 10692 5624
rect 3476 5584 3482 5596
rect 10686 5584 10692 5596
rect 10744 5584 10750 5636
rect 12710 5584 12716 5636
rect 12768 5624 12774 5636
rect 16408 5624 16436 5664
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 16666 5652 16672 5704
rect 16724 5652 16730 5704
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5692 17095 5695
rect 17129 5695 17187 5701
rect 17129 5692 17141 5695
rect 17083 5664 17141 5692
rect 17083 5661 17095 5664
rect 17037 5655 17095 5661
rect 17129 5661 17141 5664
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 17402 5652 17408 5704
rect 17460 5692 17466 5704
rect 17681 5695 17739 5701
rect 17681 5692 17693 5695
rect 17460 5664 17693 5692
rect 17460 5652 17466 5664
rect 17681 5661 17693 5664
rect 17727 5661 17739 5695
rect 17681 5655 17739 5661
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 27356 5692 27384 5732
rect 32398 5720 32404 5732
rect 32456 5720 32462 5772
rect 20680 5664 27384 5692
rect 20680 5652 20686 5664
rect 27430 5652 27436 5704
rect 27488 5692 27494 5704
rect 32309 5695 32367 5701
rect 32309 5692 32321 5695
rect 27488 5664 32321 5692
rect 27488 5652 27494 5664
rect 32309 5661 32321 5664
rect 32355 5661 32367 5695
rect 32309 5655 32367 5661
rect 32677 5695 32735 5701
rect 32677 5661 32689 5695
rect 32723 5661 32735 5695
rect 32677 5655 32735 5661
rect 12768 5596 16436 5624
rect 12768 5584 12774 5596
rect 16482 5584 16488 5636
rect 16540 5624 16546 5636
rect 16945 5627 17003 5633
rect 16945 5624 16957 5627
rect 16540 5596 16957 5624
rect 16540 5584 16546 5596
rect 16945 5593 16957 5596
rect 16991 5593 17003 5627
rect 19794 5624 19800 5636
rect 16945 5587 17003 5593
rect 17604 5596 19800 5624
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14550 5556 14556 5568
rect 13872 5528 14556 5556
rect 13872 5516 13878 5528
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 15470 5516 15476 5568
rect 15528 5516 15534 5568
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16574 5556 16580 5568
rect 15887 5528 16580 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 16850 5516 16856 5568
rect 16908 5516 16914 5568
rect 17604 5565 17632 5596
rect 19794 5584 19800 5596
rect 19852 5584 19858 5636
rect 30558 5584 30564 5636
rect 30616 5624 30622 5636
rect 32692 5624 32720 5655
rect 30616 5596 32720 5624
rect 30616 5584 30622 5596
rect 17589 5559 17647 5565
rect 17589 5525 17601 5559
rect 17635 5525 17647 5559
rect 17589 5519 17647 5525
rect 32493 5559 32551 5565
rect 32493 5525 32505 5559
rect 32539 5556 32551 5559
rect 33410 5556 33416 5568
rect 32539 5528 33416 5556
rect 32539 5525 32551 5528
rect 32493 5519 32551 5525
rect 33410 5516 33416 5528
rect 33468 5516 33474 5568
rect 1104 5466 33324 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 33324 5466
rect 1104 5392 33324 5414
rect 12066 5312 12072 5364
rect 12124 5352 12130 5364
rect 15746 5352 15752 5364
rect 12124 5324 15752 5352
rect 12124 5312 12130 5324
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 15838 5312 15844 5364
rect 15896 5352 15902 5364
rect 17402 5352 17408 5364
rect 15896 5324 17408 5352
rect 15896 5312 15902 5324
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 17644 5324 18276 5352
rect 17644 5312 17650 5324
rect 17221 5287 17279 5293
rect 17221 5253 17233 5287
rect 17267 5284 17279 5287
rect 17267 5256 17908 5284
rect 17267 5253 17279 5256
rect 17221 5247 17279 5253
rect 17880 5225 17908 5256
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5216 17095 5219
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 17083 5188 17325 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17313 5185 17325 5188
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 17589 5219 17647 5225
rect 17589 5185 17601 5219
rect 17635 5185 17647 5219
rect 17589 5179 17647 5185
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 16758 5148 16764 5160
rect 4764 5120 16764 5148
rect 4764 5108 4770 5120
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5148 16911 5151
rect 17604 5148 17632 5179
rect 18138 5176 18144 5228
rect 18196 5176 18202 5228
rect 18248 5216 18276 5324
rect 32858 5312 32864 5364
rect 32916 5312 32922 5364
rect 22066 5256 32720 5284
rect 18417 5219 18475 5225
rect 18417 5216 18429 5219
rect 18248 5188 18429 5216
rect 18417 5185 18429 5188
rect 18463 5216 18475 5219
rect 18877 5219 18935 5225
rect 18877 5216 18889 5219
rect 18463 5188 18889 5216
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 18877 5185 18889 5188
rect 18923 5185 18935 5219
rect 18877 5179 18935 5185
rect 19702 5176 19708 5228
rect 19760 5216 19766 5228
rect 22066 5216 22094 5256
rect 19760 5188 22094 5216
rect 19760 5176 19766 5188
rect 32306 5176 32312 5228
rect 32364 5176 32370 5228
rect 32692 5225 32720 5256
rect 32677 5219 32735 5225
rect 32677 5185 32689 5219
rect 32723 5185 32735 5219
rect 32677 5179 32735 5185
rect 16899 5120 17632 5148
rect 18156 5148 18184 5176
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18156 5120 18705 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18782 5108 18788 5160
rect 18840 5148 18846 5160
rect 30650 5148 30656 5160
rect 18840 5120 30656 5148
rect 18840 5108 18846 5120
rect 30650 5108 30656 5120
rect 30708 5108 30714 5160
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 14642 5080 14648 5092
rect 4120 5052 14648 5080
rect 4120 5040 4126 5052
rect 14642 5040 14648 5052
rect 14700 5040 14706 5092
rect 14918 5040 14924 5092
rect 14976 5080 14982 5092
rect 17129 5083 17187 5089
rect 17129 5080 17141 5083
rect 14976 5052 17141 5080
rect 14976 5040 14982 5052
rect 17129 5049 17141 5052
rect 17175 5049 17187 5083
rect 17129 5043 17187 5049
rect 17773 5083 17831 5089
rect 17773 5049 17785 5083
rect 17819 5080 17831 5083
rect 18506 5080 18512 5092
rect 17819 5052 18512 5080
rect 17819 5049 17831 5052
rect 17773 5043 17831 5049
rect 18506 5040 18512 5052
rect 18564 5040 18570 5092
rect 18601 5083 18659 5089
rect 18601 5049 18613 5083
rect 18647 5080 18659 5083
rect 28902 5080 28908 5092
rect 18647 5052 28908 5080
rect 18647 5049 18659 5052
rect 18601 5043 18659 5049
rect 28902 5040 28908 5052
rect 28960 5040 28966 5092
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 16761 5015 16819 5021
rect 16761 5012 16773 5015
rect 14608 4984 16773 5012
rect 14608 4972 14614 4984
rect 16761 4981 16773 4984
rect 16807 4981 16819 5015
rect 16761 4975 16819 4981
rect 16942 4972 16948 5024
rect 17000 4972 17006 5024
rect 17494 4972 17500 5024
rect 17552 4972 17558 5024
rect 18046 4972 18052 5024
rect 18104 4972 18110 5024
rect 18322 4972 18328 5024
rect 18380 4972 18386 5024
rect 26786 4972 26792 5024
rect 26844 5012 26850 5024
rect 31754 5012 31760 5024
rect 26844 4984 31760 5012
rect 26844 4972 26850 4984
rect 31754 4972 31760 4984
rect 31812 4972 31818 5024
rect 32490 4972 32496 5024
rect 32548 4972 32554 5024
rect 1104 4922 33304 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 33304 4922
rect 1104 4848 33304 4870
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 11885 4811 11943 4817
rect 11885 4808 11897 4811
rect 11572 4780 11897 4808
rect 11572 4768 11578 4780
rect 11885 4777 11897 4780
rect 11931 4777 11943 4811
rect 11885 4771 11943 4777
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 17954 4808 17960 4820
rect 14700 4780 17960 4808
rect 14700 4768 14706 4780
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 18322 4768 18328 4820
rect 18380 4808 18386 4820
rect 26878 4808 26884 4820
rect 18380 4780 26884 4808
rect 18380 4768 18386 4780
rect 26878 4768 26884 4780
rect 26936 4768 26942 4820
rect 27614 4768 27620 4820
rect 27672 4808 27678 4820
rect 28813 4811 28871 4817
rect 28813 4808 28825 4811
rect 27672 4780 28825 4808
rect 27672 4768 27678 4780
rect 28813 4777 28825 4780
rect 28859 4777 28871 4811
rect 28813 4771 28871 4777
rect 2774 4700 2780 4752
rect 2832 4740 2838 4752
rect 17862 4740 17868 4752
rect 2832 4712 17868 4740
rect 2832 4700 2838 4712
rect 17862 4700 17868 4712
rect 17920 4700 17926 4752
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 31662 4740 31668 4752
rect 18104 4712 31668 4740
rect 18104 4700 18110 4712
rect 31662 4700 31668 4712
rect 31720 4700 31726 4752
rect 32858 4700 32864 4752
rect 32916 4700 32922 4752
rect 16574 4632 16580 4684
rect 16632 4672 16638 4684
rect 16632 4644 31754 4672
rect 16632 4632 16638 4644
rect 12066 4564 12072 4616
rect 12124 4564 12130 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 12406 4576 14105 4604
rect 7834 4496 7840 4548
rect 7892 4536 7898 4548
rect 12406 4536 12434 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 28721 4607 28779 4613
rect 16448 4576 22094 4604
rect 16448 4564 16454 4576
rect 7892 4508 12434 4536
rect 7892 4496 7898 4508
rect 15746 4496 15752 4548
rect 15804 4536 15810 4548
rect 20530 4536 20536 4548
rect 15804 4508 20536 4536
rect 15804 4496 15810 4508
rect 20530 4496 20536 4508
rect 20588 4496 20594 4548
rect 22066 4536 22094 4576
rect 28721 4573 28733 4607
rect 28767 4604 28779 4607
rect 28997 4607 29055 4613
rect 28997 4604 29009 4607
rect 28767 4576 29009 4604
rect 28767 4573 28779 4576
rect 28721 4567 28779 4573
rect 28997 4573 29009 4576
rect 29043 4573 29055 4607
rect 31726 4604 31754 4644
rect 32309 4607 32367 4613
rect 32309 4604 32321 4607
rect 31726 4576 32321 4604
rect 28997 4567 29055 4573
rect 32309 4573 32321 4576
rect 32355 4573 32367 4607
rect 32309 4567 32367 4573
rect 32677 4607 32735 4613
rect 32677 4573 32689 4607
rect 32723 4573 32735 4607
rect 32677 4567 32735 4573
rect 32692 4536 32720 4567
rect 22066 4508 32720 4536
rect 14277 4471 14335 4477
rect 14277 4437 14289 4471
rect 14323 4468 14335 4471
rect 17126 4468 17132 4480
rect 14323 4440 17132 4468
rect 14323 4437 14335 4440
rect 14277 4431 14335 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 18690 4428 18696 4480
rect 18748 4468 18754 4480
rect 28629 4471 28687 4477
rect 28629 4468 28641 4471
rect 18748 4440 28641 4468
rect 18748 4428 18754 4440
rect 28629 4437 28641 4440
rect 28675 4437 28687 4471
rect 28629 4431 28687 4437
rect 28902 4428 28908 4480
rect 28960 4468 28966 4480
rect 32398 4468 32404 4480
rect 28960 4440 32404 4468
rect 28960 4428 28966 4440
rect 32398 4428 32404 4440
rect 32456 4428 32462 4480
rect 32493 4471 32551 4477
rect 32493 4437 32505 4471
rect 32539 4468 32551 4471
rect 33410 4468 33416 4480
rect 32539 4440 33416 4468
rect 32539 4437 32551 4440
rect 32493 4431 32551 4437
rect 33410 4428 33416 4440
rect 33468 4428 33474 4480
rect 1104 4378 33324 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 33324 4378
rect 1104 4304 33324 4326
rect 12342 4224 12348 4276
rect 12400 4264 12406 4276
rect 12897 4267 12955 4273
rect 12897 4264 12909 4267
rect 12400 4236 12909 4264
rect 12400 4224 12406 4236
rect 12897 4233 12909 4236
rect 12943 4233 12955 4267
rect 13078 4264 13084 4276
rect 12897 4227 12955 4233
rect 13004 4236 13084 4264
rect 3418 4088 3424 4140
rect 3476 4128 3482 4140
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 3476 4100 7573 4128
rect 3476 4088 3482 4100
rect 7561 4097 7573 4100
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10100 4100 11652 4128
rect 10100 4088 10106 4100
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 10376 3964 11529 3992
rect 10376 3952 10382 3964
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 11624 3992 11652 4100
rect 11698 4088 11704 4140
rect 11756 4088 11762 4140
rect 11974 4088 11980 4140
rect 12032 4088 12038 4140
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12529 4131 12587 4137
rect 12299 4100 12434 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 11848 4032 12112 4060
rect 11848 4020 11854 4032
rect 12084 4001 12112 4032
rect 12069 3995 12127 4001
rect 11624 3964 11928 3992
rect 11517 3955 11575 3961
rect 7742 3884 7748 3936
rect 7800 3884 7806 3936
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 9824 3896 11805 3924
rect 9824 3884 9830 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 11900 3924 11928 3964
rect 12069 3961 12081 3995
rect 12115 3961 12127 3995
rect 12406 3992 12434 4100
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4128 12863 4131
rect 13004 4128 13032 4236
rect 13078 4224 13084 4236
rect 13136 4224 13142 4276
rect 17494 4224 17500 4276
rect 17552 4264 17558 4276
rect 26786 4264 26792 4276
rect 17552 4236 26792 4264
rect 17552 4224 17558 4236
rect 26786 4224 26792 4236
rect 26844 4224 26850 4276
rect 26878 4224 26884 4276
rect 26936 4264 26942 4276
rect 26936 4236 32720 4264
rect 26936 4224 26942 4236
rect 14826 4156 14832 4208
rect 14884 4196 14890 4208
rect 15378 4196 15384 4208
rect 14884 4168 15384 4196
rect 14884 4156 14890 4168
rect 15378 4156 15384 4168
rect 15436 4156 15442 4208
rect 12851 4100 13032 4128
rect 13081 4131 13139 4137
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 16482 4128 16488 4140
rect 13127 4100 16488 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 12544 4060 12572 4091
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 31662 4088 31668 4140
rect 31720 4128 31726 4140
rect 32692 4137 32720 4236
rect 32309 4131 32367 4137
rect 32309 4128 32321 4131
rect 31720 4100 32321 4128
rect 31720 4088 31726 4100
rect 32309 4097 32321 4100
rect 32355 4097 32367 4131
rect 32309 4091 32367 4097
rect 32677 4131 32735 4137
rect 32677 4097 32689 4131
rect 32723 4097 32735 4131
rect 32677 4091 32735 4097
rect 16390 4060 16396 4072
rect 12544 4032 16396 4060
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 22646 4060 22652 4072
rect 17276 4032 22652 4060
rect 17276 4020 17282 4032
rect 22646 4020 22652 4032
rect 22704 4020 22710 4072
rect 12406 3964 12572 3992
rect 12069 3955 12127 3961
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 11900 3896 12357 3924
rect 11793 3887 11851 3893
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12544 3924 12572 3964
rect 12618 3952 12624 4004
rect 12676 3952 12682 4004
rect 32858 3952 32864 4004
rect 32916 3952 32922 4004
rect 19334 3924 19340 3936
rect 12544 3896 19340 3924
rect 12345 3887 12403 3893
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 21082 3884 21088 3936
rect 21140 3924 21146 3936
rect 25314 3924 25320 3936
rect 21140 3896 25320 3924
rect 21140 3884 21146 3896
rect 25314 3884 25320 3896
rect 25372 3884 25378 3936
rect 32490 3884 32496 3936
rect 32548 3884 32554 3936
rect 1104 3834 33304 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 33304 3834
rect 1104 3760 33304 3782
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 8386 3720 8392 3732
rect 7340 3692 8392 3720
rect 7340 3680 7346 3692
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 10502 3680 10508 3732
rect 10560 3680 10566 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 12069 3723 12127 3729
rect 12069 3720 12081 3723
rect 11112 3692 12081 3720
rect 11112 3680 11118 3692
rect 12069 3689 12081 3692
rect 12115 3689 12127 3723
rect 12069 3683 12127 3689
rect 14461 3723 14519 3729
rect 14461 3689 14473 3723
rect 14507 3720 14519 3723
rect 15102 3720 15108 3732
rect 14507 3692 15108 3720
rect 14507 3689 14519 3692
rect 14461 3683 14519 3689
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 15378 3680 15384 3732
rect 15436 3680 15442 3732
rect 18049 3723 18107 3729
rect 15488 3692 18000 3720
rect 11333 3655 11391 3661
rect 11333 3621 11345 3655
rect 11379 3621 11391 3655
rect 11333 3615 11391 3621
rect 11348 3584 11376 3615
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 15488 3652 15516 3692
rect 11756 3624 15516 3652
rect 11756 3612 11762 3624
rect 15562 3612 15568 3664
rect 15620 3652 15626 3664
rect 15620 3624 17356 3652
rect 15620 3612 15626 3624
rect 17218 3584 17224 3596
rect 11348 3556 17224 3584
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 17328 3584 17356 3624
rect 17770 3612 17776 3664
rect 17828 3612 17834 3664
rect 17972 3652 18000 3692
rect 18049 3689 18061 3723
rect 18095 3720 18107 3723
rect 18782 3720 18788 3732
rect 18095 3692 18788 3720
rect 18095 3689 18107 3692
rect 18049 3683 18107 3689
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 19610 3680 19616 3732
rect 19668 3720 19674 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19668 3692 19809 3720
rect 19668 3680 19674 3692
rect 19797 3689 19809 3692
rect 19843 3689 19855 3723
rect 20346 3720 20352 3732
rect 19797 3683 19855 3689
rect 20088 3692 20352 3720
rect 18414 3652 18420 3664
rect 17972 3624 18420 3652
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 19429 3655 19487 3661
rect 19429 3621 19441 3655
rect 19475 3652 19487 3655
rect 20088 3652 20116 3692
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20622 3680 20628 3732
rect 20680 3680 20686 3732
rect 21082 3680 21088 3732
rect 21140 3680 21146 3732
rect 23201 3723 23259 3729
rect 23201 3689 23213 3723
rect 23247 3720 23259 3723
rect 24854 3720 24860 3732
rect 23247 3692 24860 3720
rect 23247 3689 23259 3692
rect 23201 3683 23259 3689
rect 24854 3680 24860 3692
rect 24912 3680 24918 3732
rect 27249 3723 27307 3729
rect 27249 3689 27261 3723
rect 27295 3720 27307 3723
rect 27338 3720 27344 3732
rect 27295 3692 27344 3720
rect 27295 3689 27307 3692
rect 27249 3683 27307 3689
rect 27338 3680 27344 3692
rect 27396 3680 27402 3732
rect 28350 3680 28356 3732
rect 28408 3720 28414 3732
rect 28905 3723 28963 3729
rect 28905 3720 28917 3723
rect 28408 3692 28917 3720
rect 28408 3680 28414 3692
rect 28905 3689 28917 3692
rect 28951 3689 28963 3723
rect 28905 3683 28963 3689
rect 19475 3624 20116 3652
rect 20165 3655 20223 3661
rect 19475 3621 19487 3624
rect 19429 3615 19487 3621
rect 20165 3621 20177 3655
rect 20211 3652 20223 3655
rect 27430 3652 27436 3664
rect 20211 3624 27436 3652
rect 20211 3621 20223 3624
rect 20165 3615 20223 3621
rect 27430 3612 27436 3624
rect 27488 3612 27494 3664
rect 27982 3612 27988 3664
rect 28040 3652 28046 3664
rect 29641 3655 29699 3661
rect 29641 3652 29653 3655
rect 28040 3624 29653 3652
rect 28040 3612 28046 3624
rect 29641 3621 29653 3624
rect 29687 3621 29699 3655
rect 29641 3615 29699 3621
rect 32858 3612 32864 3664
rect 32916 3612 32922 3664
rect 17328 3556 29132 3584
rect 1486 3476 1492 3528
rect 1544 3516 1550 3528
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 1544 3488 10333 3516
rect 1544 3476 1550 3488
rect 10321 3485 10333 3488
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 14182 3516 14188 3528
rect 12299 3488 14188 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 4614 3408 4620 3460
rect 4672 3448 4678 3460
rect 11164 3448 11192 3479
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3516 15531 3519
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 15519 3488 15577 3516
rect 15519 3485 15531 3488
rect 15473 3479 15531 3485
rect 15565 3485 15577 3488
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 16816 3488 17601 3516
rect 16816 3476 16822 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 17862 3476 17868 3528
rect 17920 3476 17926 3528
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 18012 3488 19257 3516
rect 18012 3476 18018 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19889 3519 19947 3525
rect 19889 3485 19901 3519
rect 19935 3516 19947 3519
rect 19981 3519 20039 3525
rect 19981 3516 19993 3519
rect 19935 3488 19993 3516
rect 19935 3485 19947 3488
rect 19889 3479 19947 3485
rect 19981 3485 19993 3488
rect 20027 3485 20039 3519
rect 19981 3479 20039 3485
rect 20438 3476 20444 3528
rect 20496 3476 20502 3528
rect 20901 3519 20959 3525
rect 20901 3485 20913 3519
rect 20947 3485 20959 3519
rect 20901 3479 20959 3485
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3516 21511 3519
rect 21545 3519 21603 3525
rect 21545 3516 21557 3519
rect 21499 3488 21557 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 21545 3485 21557 3488
rect 21591 3485 21603 3519
rect 21545 3479 21603 3485
rect 22925 3519 22983 3525
rect 22925 3485 22937 3519
rect 22971 3516 22983 3519
rect 23017 3519 23075 3525
rect 23017 3516 23029 3519
rect 22971 3488 23029 3516
rect 22971 3485 22983 3488
rect 22925 3479 22983 3485
rect 23017 3485 23029 3488
rect 23063 3485 23075 3519
rect 23017 3479 23075 3485
rect 4672 3420 11192 3448
rect 4672 3408 4678 3420
rect 16666 3408 16672 3460
rect 16724 3448 16730 3460
rect 20916 3448 20944 3479
rect 24854 3476 24860 3528
rect 24912 3516 24918 3528
rect 29104 3525 29132 3556
rect 27065 3519 27123 3525
rect 27065 3516 27077 3519
rect 24912 3488 27077 3516
rect 24912 3476 24918 3488
rect 27065 3485 27077 3488
rect 27111 3485 27123 3519
rect 27065 3479 27123 3485
rect 29089 3519 29147 3525
rect 29089 3485 29101 3519
rect 29135 3485 29147 3519
rect 29089 3479 29147 3485
rect 29825 3519 29883 3525
rect 29825 3485 29837 3519
rect 29871 3485 29883 3519
rect 29825 3479 29883 3485
rect 27522 3448 27528 3460
rect 16724 3420 20944 3448
rect 22066 3420 27528 3448
rect 16724 3408 16730 3420
rect 15746 3340 15752 3392
rect 15804 3340 15810 3392
rect 21358 3340 21364 3392
rect 21416 3340 21422 3392
rect 21729 3383 21787 3389
rect 21729 3349 21741 3383
rect 21775 3380 21787 3383
rect 22066 3380 22094 3420
rect 27522 3408 27528 3420
rect 27580 3408 27586 3460
rect 27614 3408 27620 3460
rect 27672 3448 27678 3460
rect 29840 3448 29868 3479
rect 30650 3476 30656 3528
rect 30708 3516 30714 3528
rect 32309 3519 32367 3525
rect 32309 3516 32321 3519
rect 30708 3488 32321 3516
rect 30708 3476 30714 3488
rect 32309 3485 32321 3488
rect 32355 3485 32367 3519
rect 32309 3479 32367 3485
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 32677 3519 32735 3525
rect 32677 3516 32689 3519
rect 32456 3488 32689 3516
rect 32456 3476 32462 3488
rect 32677 3485 32689 3488
rect 32723 3485 32735 3519
rect 32677 3479 32735 3485
rect 27672 3420 29868 3448
rect 27672 3408 27678 3420
rect 21775 3352 22094 3380
rect 21775 3349 21787 3352
rect 21729 3343 21787 3349
rect 22830 3340 22836 3392
rect 22888 3340 22894 3392
rect 32493 3383 32551 3389
rect 32493 3349 32505 3383
rect 32539 3380 32551 3383
rect 33410 3380 33416 3392
rect 32539 3352 33416 3380
rect 32539 3349 32551 3352
rect 32493 3343 32551 3349
rect 33410 3340 33416 3352
rect 33468 3340 33474 3392
rect 1104 3290 33324 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 33324 3290
rect 1104 3216 33324 3238
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 22830 3176 22836 3188
rect 12492 3148 22836 3176
rect 12492 3136 12498 3148
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 32858 3136 32864 3188
rect 32916 3136 32922 3188
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 14274 3108 14280 3120
rect 6236 3080 14280 3108
rect 6236 3068 6242 3080
rect 14274 3068 14280 3080
rect 14332 3068 14338 3120
rect 18506 3068 18512 3120
rect 18564 3108 18570 3120
rect 31846 3108 31852 3120
rect 18564 3080 31852 3108
rect 18564 3068 18570 3080
rect 31846 3068 31852 3080
rect 31904 3068 31910 3120
rect 32030 3068 32036 3120
rect 32088 3108 32094 3120
rect 32088 3080 32720 3108
rect 32088 3068 32094 3080
rect 14458 3000 14464 3052
rect 14516 3040 14522 3052
rect 32692 3049 32720 3080
rect 31665 3043 31723 3049
rect 31665 3040 31677 3043
rect 14516 3012 31677 3040
rect 14516 3000 14522 3012
rect 31665 3009 31677 3012
rect 31711 3009 31723 3043
rect 31665 3003 31723 3009
rect 32309 3043 32367 3049
rect 32309 3009 32321 3043
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 32677 3043 32735 3049
rect 32677 3009 32689 3043
rect 32723 3009 32735 3043
rect 32677 3003 32735 3009
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 21542 2972 21548 2984
rect 7800 2944 21548 2972
rect 7800 2932 7806 2944
rect 21542 2932 21548 2944
rect 21600 2932 21606 2984
rect 30650 2972 30656 2984
rect 22066 2944 30656 2972
rect 14366 2864 14372 2916
rect 14424 2904 14430 2916
rect 22066 2904 22094 2944
rect 30650 2932 30656 2944
rect 30708 2932 30714 2984
rect 14424 2876 22094 2904
rect 14424 2864 14430 2876
rect 30374 2864 30380 2916
rect 30432 2904 30438 2916
rect 32324 2904 32352 3003
rect 30432 2876 32352 2904
rect 30432 2864 30438 2876
rect 15746 2796 15752 2848
rect 15804 2836 15810 2848
rect 30558 2836 30564 2848
rect 15804 2808 30564 2836
rect 15804 2796 15810 2808
rect 30558 2796 30564 2808
rect 30616 2796 30622 2848
rect 31846 2796 31852 2848
rect 31904 2796 31910 2848
rect 32490 2796 32496 2848
rect 32548 2796 32554 2848
rect 1104 2746 33304 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 33304 2746
rect 1104 2672 33304 2694
rect 16022 2592 16028 2644
rect 16080 2632 16086 2644
rect 31294 2632 31300 2644
rect 16080 2604 31300 2632
rect 16080 2592 16086 2604
rect 31294 2592 31300 2604
rect 31352 2592 31358 2644
rect 16850 2524 16856 2576
rect 16908 2564 16914 2576
rect 16908 2536 31156 2564
rect 16908 2524 16914 2536
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 31128 2496 31156 2536
rect 32858 2524 32864 2576
rect 32916 2524 32922 2576
rect 14792 2468 31064 2496
rect 31128 2468 32720 2496
rect 14792 2456 14798 2468
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 13780 2400 30941 2428
rect 13780 2388 13786 2400
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 3510 2320 3516 2372
rect 3568 2360 3574 2372
rect 20438 2360 20444 2372
rect 3568 2332 20444 2360
rect 3568 2320 3574 2332
rect 20438 2320 20444 2332
rect 20496 2320 20502 2372
rect 31036 2360 31064 2468
rect 31294 2388 31300 2440
rect 31352 2388 31358 2440
rect 31665 2431 31723 2437
rect 31665 2397 31677 2431
rect 31711 2397 31723 2431
rect 31665 2391 31723 2397
rect 31680 2360 31708 2391
rect 31754 2388 31760 2440
rect 31812 2428 31818 2440
rect 32692 2437 32720 2468
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31812 2400 32321 2428
rect 31812 2388 31818 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 32677 2431 32735 2437
rect 32677 2397 32689 2431
rect 32723 2397 32735 2431
rect 32677 2391 32735 2397
rect 31036 2332 31708 2360
rect 20254 2252 20260 2304
rect 20312 2292 20318 2304
rect 29270 2292 29276 2304
rect 20312 2264 29276 2292
rect 20312 2252 20318 2264
rect 29270 2252 29276 2264
rect 29328 2252 29334 2304
rect 31110 2252 31116 2304
rect 31168 2252 31174 2304
rect 31478 2252 31484 2304
rect 31536 2252 31542 2304
rect 31846 2252 31852 2304
rect 31904 2252 31910 2304
rect 32493 2295 32551 2301
rect 32493 2261 32505 2295
rect 32539 2292 32551 2295
rect 33410 2292 33416 2304
rect 32539 2264 33416 2292
rect 32539 2261 32551 2264
rect 32493 2255 32551 2261
rect 33410 2252 33416 2264
rect 33468 2252 33474 2304
rect 1104 2202 33324 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 33324 2202
rect 1104 2128 33324 2150
rect 10870 2048 10876 2100
rect 10928 2088 10934 2100
rect 21358 2088 21364 2100
rect 10928 2060 21364 2088
rect 10928 2048 10934 2060
rect 21358 2048 21364 2060
rect 21416 2048 21422 2100
rect 14090 8 14096 60
rect 14148 48 14154 60
rect 24854 48 24860 60
rect 14148 20 24860 48
rect 14148 8 14154 20
rect 24854 8 24860 20
rect 24912 8 24918 60
<< via1 >>
rect 7564 11092 7616 11144
rect 18052 11092 18104 11144
rect 7012 11024 7064 11076
rect 17960 10956 18012 11008
rect 9588 10820 9640 10872
rect 18696 10820 18748 10872
rect 10692 10616 10744 10668
rect 16120 10616 16172 10668
rect 14372 10548 14424 10600
rect 15752 10548 15804 10600
rect 11980 10480 12032 10532
rect 17776 10480 17828 10532
rect 13268 10140 13320 10192
rect 19800 10140 19852 10192
rect 16672 9936 16724 9988
rect 20168 9936 20220 9988
rect 13636 9732 13688 9784
rect 19248 9732 19300 9784
rect 18420 9596 18472 9648
rect 20720 9596 20772 9648
rect 15660 9528 15712 9580
rect 26700 9528 26752 9580
rect 13452 9460 13504 9512
rect 24400 9460 24452 9512
rect 8668 9392 8720 9444
rect 9312 9392 9364 9444
rect 19524 9392 19576 9444
rect 31668 9392 31720 9444
rect 1308 9324 1360 9376
rect 19708 9324 19760 9376
rect 1032 9256 1084 9308
rect 19616 9256 19668 9308
rect 19800 9256 19852 9308
rect 32312 9256 32364 9308
rect 13820 9188 13872 9240
rect 24676 9188 24728 9240
rect 21088 9120 21140 9172
rect 21732 9120 21784 9172
rect 296 8984 348 9036
rect 20444 8984 20496 9036
rect 10324 8916 10376 8968
rect 12532 8916 12584 8968
rect 12900 8916 12952 8968
rect 18052 8916 18104 8968
rect 22744 8916 22796 8968
rect 25596 8916 25648 8968
rect 27528 8916 27580 8968
rect 28540 8916 28592 8968
rect 7196 8848 7248 8900
rect 7932 8848 7984 8900
rect 10140 8848 10192 8900
rect 10784 8848 10836 8900
rect 10876 8848 10928 8900
rect 12164 8848 12216 8900
rect 12348 8848 12400 8900
rect 12992 8848 13044 8900
rect 6460 8780 6512 8832
rect 8116 8780 8168 8832
rect 10508 8780 10560 8832
rect 11152 8780 11204 8832
rect 12716 8780 12768 8832
rect 20904 8848 20956 8900
rect 21364 8848 21416 8900
rect 32680 8848 32732 8900
rect 14556 8780 14608 8832
rect 25044 8780 25096 8832
rect 27160 8780 27212 8832
rect 27528 8780 27580 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 5632 8576 5684 8628
rect 6736 8576 6788 8628
rect 7472 8576 7524 8628
rect 7748 8576 7800 8628
rect 6368 8508 6420 8560
rect 8852 8576 8904 8628
rect 10048 8576 10100 8628
rect 10508 8576 10560 8628
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 5264 8440 5316 8492
rect 5448 8372 5500 8424
rect 4160 8304 4212 8356
rect 6000 8304 6052 8356
rect 8576 8508 8628 8560
rect 7472 8440 7524 8492
rect 7380 8372 7432 8424
rect 7564 8372 7616 8424
rect 7932 8440 7984 8492
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 10324 8508 10376 8560
rect 11060 8576 11112 8628
rect 11888 8576 11940 8628
rect 12348 8576 12400 8628
rect 13360 8576 13412 8628
rect 14096 8576 14148 8628
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 14648 8576 14700 8628
rect 14924 8576 14976 8628
rect 9772 8440 9824 8492
rect 10784 8440 10836 8492
rect 11244 8440 11296 8492
rect 11612 8440 11664 8492
rect 12716 8508 12768 8560
rect 24952 8619 25004 8628
rect 24952 8585 24961 8619
rect 24961 8585 24995 8619
rect 24995 8585 25004 8619
rect 24952 8576 25004 8585
rect 25136 8576 25188 8628
rect 25504 8576 25556 8628
rect 10324 8372 10376 8424
rect 7748 8304 7800 8356
rect 8208 8304 8260 8356
rect 8668 8304 8720 8356
rect 10416 8304 10468 8356
rect 11520 8304 11572 8356
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 11152 8236 11204 8288
rect 11428 8236 11480 8288
rect 12624 8236 12676 8288
rect 12900 8440 12952 8492
rect 13452 8440 13504 8492
rect 13820 8440 13872 8492
rect 14556 8440 14608 8492
rect 25688 8508 25740 8560
rect 26792 8576 26844 8628
rect 14924 8440 14976 8492
rect 15660 8440 15712 8492
rect 24492 8440 24544 8492
rect 25136 8483 25188 8492
rect 25136 8449 25145 8483
rect 25145 8449 25179 8483
rect 25179 8449 25188 8483
rect 25136 8440 25188 8449
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 25504 8440 25556 8492
rect 13728 8372 13780 8424
rect 22652 8372 22704 8424
rect 25780 8440 25832 8492
rect 26424 8440 26476 8492
rect 27344 8483 27396 8492
rect 27344 8449 27353 8483
rect 27353 8449 27387 8483
rect 27387 8449 27396 8483
rect 27344 8440 27396 8449
rect 27528 8508 27580 8560
rect 28540 8619 28592 8628
rect 28540 8585 28549 8619
rect 28549 8585 28583 8619
rect 28583 8585 28592 8619
rect 28540 8576 28592 8585
rect 28632 8576 28684 8628
rect 31484 8619 31536 8628
rect 31484 8585 31493 8619
rect 31493 8585 31527 8619
rect 31527 8585 31536 8619
rect 31484 8576 31536 8585
rect 31852 8619 31904 8628
rect 31852 8585 31861 8619
rect 31861 8585 31895 8619
rect 31895 8585 31904 8619
rect 31852 8576 31904 8585
rect 27620 8440 27672 8492
rect 27988 8483 28040 8492
rect 27988 8449 27997 8483
rect 27997 8449 28031 8483
rect 28031 8449 28040 8483
rect 27988 8440 28040 8449
rect 28632 8440 28684 8492
rect 28724 8483 28776 8492
rect 28724 8449 28733 8483
rect 28733 8449 28767 8483
rect 28767 8449 28776 8483
rect 28724 8440 28776 8449
rect 28908 8440 28960 8492
rect 29828 8483 29880 8492
rect 29828 8449 29837 8483
rect 29837 8449 29871 8483
rect 29871 8449 29880 8483
rect 29828 8440 29880 8449
rect 31300 8483 31352 8492
rect 31300 8449 31309 8483
rect 31309 8449 31343 8483
rect 31343 8449 31352 8483
rect 31300 8440 31352 8449
rect 31668 8483 31720 8492
rect 31668 8449 31677 8483
rect 31677 8449 31711 8483
rect 31711 8449 31720 8483
rect 31668 8440 31720 8449
rect 32312 8483 32364 8492
rect 32312 8449 32321 8483
rect 32321 8449 32355 8483
rect 32355 8449 32364 8483
rect 32312 8440 32364 8449
rect 32680 8483 32732 8492
rect 32680 8449 32689 8483
rect 32689 8449 32723 8483
rect 32723 8449 32732 8483
rect 32680 8440 32732 8449
rect 26516 8372 26568 8424
rect 13820 8304 13872 8356
rect 14832 8304 14884 8356
rect 14556 8236 14608 8288
rect 15384 8304 15436 8356
rect 22928 8304 22980 8356
rect 25136 8304 25188 8356
rect 25320 8304 25372 8356
rect 26056 8304 26108 8356
rect 27896 8304 27948 8356
rect 32496 8347 32548 8356
rect 32496 8313 32505 8347
rect 32505 8313 32539 8347
rect 32539 8313 32548 8347
rect 32496 8304 32548 8313
rect 32864 8347 32916 8356
rect 32864 8313 32873 8347
rect 32873 8313 32907 8347
rect 32907 8313 32916 8347
rect 32864 8304 32916 8313
rect 16212 8236 16264 8288
rect 19984 8236 20036 8288
rect 24768 8236 24820 8288
rect 31668 8236 31720 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 5816 8032 5868 8084
rect 6184 8032 6236 8084
rect 6552 8032 6604 8084
rect 6920 8032 6972 8084
rect 7288 8032 7340 8084
rect 7656 8032 7708 8084
rect 7840 8075 7892 8084
rect 7840 8041 7849 8075
rect 7849 8041 7883 8075
rect 7883 8041 7892 8075
rect 7840 8032 7892 8041
rect 8392 8032 8444 8084
rect 8760 8032 8812 8084
rect 9496 8032 9548 8084
rect 9864 8032 9916 8084
rect 10232 8032 10284 8084
rect 10600 8032 10652 8084
rect 10968 8032 11020 8084
rect 11336 8032 11388 8084
rect 11704 8032 11756 8084
rect 12072 8032 12124 8084
rect 12256 8075 12308 8084
rect 12256 8041 12265 8075
rect 12265 8041 12299 8075
rect 12299 8041 12308 8075
rect 12256 8032 12308 8041
rect 12440 8032 12492 8084
rect 12808 8032 12860 8084
rect 13176 8032 13228 8084
rect 13544 8032 13596 8084
rect 14280 8032 14332 8084
rect 2136 7964 2188 8016
rect 8484 7964 8536 8016
rect 7472 7896 7524 7948
rect 2780 7828 2832 7880
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 6736 7828 6788 7880
rect 4344 7760 4396 7812
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 11428 7964 11480 8016
rect 8392 7760 8444 7812
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 11520 7896 11572 7948
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 11888 7964 11940 8016
rect 22928 8032 22980 8084
rect 25872 8032 25924 8084
rect 26332 8032 26384 8084
rect 26608 8032 26660 8084
rect 26884 8032 26936 8084
rect 27436 8032 27488 8084
rect 27712 8032 27764 8084
rect 28080 8032 28132 8084
rect 28356 8032 28408 8084
rect 31760 8075 31812 8084
rect 31760 8041 31769 8075
rect 31769 8041 31803 8075
rect 31803 8041 31812 8075
rect 31760 8032 31812 8041
rect 33416 8032 33468 8084
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 10048 7760 10100 7812
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 17868 7964 17920 8016
rect 18512 7896 18564 7948
rect 13360 7760 13412 7812
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 25320 7828 25372 7880
rect 20352 7760 20404 7812
rect 24860 7760 24912 7812
rect 27620 7828 27672 7880
rect 27712 7871 27764 7880
rect 27712 7837 27721 7871
rect 27721 7837 27755 7871
rect 27755 7837 27764 7871
rect 27712 7828 27764 7837
rect 27804 7871 27856 7880
rect 27804 7837 27813 7871
rect 27813 7837 27847 7871
rect 27847 7837 27856 7871
rect 27804 7828 27856 7837
rect 28356 7760 28408 7812
rect 28816 7871 28868 7880
rect 28816 7837 28825 7871
rect 28825 7837 28859 7871
rect 28859 7837 28868 7871
rect 28816 7828 28868 7837
rect 30656 7828 30708 7880
rect 32404 7896 32456 7948
rect 31668 7828 31720 7880
rect 32312 7871 32364 7880
rect 32312 7837 32321 7871
rect 32321 7837 32355 7871
rect 32355 7837 32364 7871
rect 32312 7828 32364 7837
rect 32680 7871 32732 7880
rect 32680 7837 32689 7871
rect 32689 7837 32723 7871
rect 32723 7837 32732 7871
rect 32680 7828 32732 7837
rect 29092 7760 29144 7812
rect 2504 7692 2556 7744
rect 10600 7692 10652 7744
rect 10968 7692 11020 7744
rect 12532 7692 12584 7744
rect 16856 7692 16908 7744
rect 20260 7692 20312 7744
rect 22192 7692 22244 7744
rect 26700 7692 26752 7744
rect 28448 7692 28500 7744
rect 32496 7735 32548 7744
rect 32496 7701 32505 7735
rect 32505 7701 32539 7735
rect 32539 7701 32548 7735
rect 32496 7692 32548 7701
rect 33600 7692 33652 7744
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 5908 7488 5960 7540
rect 7104 7488 7156 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 9680 7488 9732 7540
rect 11152 7488 11204 7540
rect 11796 7488 11848 7540
rect 11888 7488 11940 7540
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 11060 7420 11112 7472
rect 12532 7531 12584 7540
rect 12532 7497 12541 7531
rect 12541 7497 12575 7531
rect 12575 7497 12584 7531
rect 12532 7488 12584 7497
rect 12716 7488 12768 7540
rect 13360 7488 13412 7540
rect 16304 7488 16356 7540
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 16580 7488 16632 7540
rect 17868 7488 17920 7540
rect 18512 7531 18564 7540
rect 18512 7497 18521 7531
rect 18521 7497 18555 7531
rect 18555 7497 18564 7531
rect 18512 7488 18564 7497
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3976 7352 4028 7404
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 10968 7352 11020 7404
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 4804 7284 4856 7336
rect 5172 7216 5224 7268
rect 10232 7216 10284 7268
rect 11060 7216 11112 7268
rect 11244 7216 11296 7268
rect 12532 7352 12584 7404
rect 16672 7420 16724 7472
rect 19524 7531 19576 7540
rect 19524 7497 19533 7531
rect 19533 7497 19567 7531
rect 19567 7497 19576 7531
rect 19524 7488 19576 7497
rect 19800 7531 19852 7540
rect 19800 7497 19809 7531
rect 19809 7497 19843 7531
rect 19843 7497 19852 7531
rect 19800 7488 19852 7497
rect 20720 7531 20772 7540
rect 20720 7497 20729 7531
rect 20729 7497 20763 7531
rect 20763 7497 20772 7531
rect 20720 7488 20772 7497
rect 21272 7488 21324 7540
rect 21548 7488 21600 7540
rect 25228 7488 25280 7540
rect 27804 7531 27856 7540
rect 27804 7497 27813 7531
rect 27813 7497 27847 7531
rect 27847 7497 27856 7531
rect 27804 7488 27856 7497
rect 28724 7488 28776 7540
rect 28908 7531 28960 7540
rect 28908 7497 28917 7531
rect 28917 7497 28951 7531
rect 28951 7497 28960 7531
rect 28908 7488 28960 7497
rect 29092 7488 29144 7540
rect 29828 7488 29880 7540
rect 30656 7531 30708 7540
rect 30656 7497 30665 7531
rect 30665 7497 30699 7531
rect 30699 7497 30708 7531
rect 30656 7488 30708 7497
rect 32588 7488 32640 7540
rect 16212 7352 16264 7404
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 19616 7395 19668 7404
rect 19616 7361 19625 7395
rect 19625 7361 19659 7395
rect 19659 7361 19668 7395
rect 19616 7352 19668 7361
rect 19708 7352 19760 7404
rect 20444 7395 20496 7404
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 24768 7352 24820 7404
rect 24952 7352 25004 7404
rect 28080 7352 28132 7404
rect 28448 7352 28500 7404
rect 12440 7216 12492 7268
rect 12808 7284 12860 7336
rect 19800 7284 19852 7336
rect 16856 7216 16908 7268
rect 17960 7216 18012 7268
rect 18144 7259 18196 7268
rect 18144 7225 18153 7259
rect 18153 7225 18187 7259
rect 18187 7225 18196 7259
rect 18144 7216 18196 7225
rect 26792 7284 26844 7336
rect 29092 7395 29144 7404
rect 29092 7361 29101 7395
rect 29101 7361 29135 7395
rect 29135 7361 29144 7395
rect 29092 7352 29144 7361
rect 29368 7395 29420 7404
rect 29368 7361 29377 7395
rect 29377 7361 29411 7395
rect 29411 7361 29420 7395
rect 29368 7352 29420 7361
rect 32772 7420 32824 7472
rect 26884 7216 26936 7268
rect 27712 7216 27764 7268
rect 3148 7148 3200 7200
rect 10876 7148 10928 7200
rect 10968 7148 11020 7200
rect 12348 7148 12400 7200
rect 12532 7148 12584 7200
rect 13268 7148 13320 7200
rect 17776 7148 17828 7200
rect 21180 7148 21232 7200
rect 29644 7284 29696 7336
rect 31208 7352 31260 7404
rect 28816 7216 28868 7268
rect 32404 7352 32456 7404
rect 30196 7148 30248 7200
rect 32680 7216 32732 7268
rect 32864 7191 32916 7200
rect 32864 7157 32873 7191
rect 32873 7157 32907 7191
rect 32907 7157 32916 7191
rect 32864 7148 32916 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 3976 6987 4028 6996
rect 3976 6953 3985 6987
rect 3985 6953 4019 6987
rect 4019 6953 4028 6987
rect 3976 6944 4028 6953
rect 11704 6944 11756 6996
rect 12440 6944 12492 6996
rect 15568 6944 15620 6996
rect 24584 6944 24636 6996
rect 3332 6740 3384 6792
rect 4436 6876 4488 6928
rect 11152 6876 11204 6928
rect 19064 6876 19116 6928
rect 23112 6876 23164 6928
rect 6828 6808 6880 6860
rect 6920 6740 6972 6792
rect 4344 6672 4396 6724
rect 4436 6672 4488 6724
rect 9956 6808 10008 6860
rect 12900 6808 12952 6860
rect 12992 6808 13044 6860
rect 17040 6808 17092 6860
rect 23296 6808 23348 6860
rect 13636 6740 13688 6792
rect 14556 6740 14608 6792
rect 21916 6740 21968 6792
rect 23480 6740 23532 6792
rect 26884 6944 26936 6996
rect 32312 6944 32364 6996
rect 26792 6876 26844 6928
rect 30196 6876 30248 6928
rect 25136 6783 25188 6792
rect 25136 6749 25145 6783
rect 25145 6749 25179 6783
rect 25179 6749 25188 6783
rect 25136 6740 25188 6749
rect 25596 6783 25648 6792
rect 25596 6749 25605 6783
rect 25605 6749 25639 6783
rect 25639 6749 25648 6783
rect 25596 6740 25648 6749
rect 26332 6783 26384 6792
rect 26332 6749 26341 6783
rect 26341 6749 26375 6783
rect 26375 6749 26384 6783
rect 26332 6740 26384 6749
rect 26700 6783 26752 6792
rect 26700 6749 26709 6783
rect 26709 6749 26743 6783
rect 26743 6749 26752 6783
rect 26700 6740 26752 6749
rect 26976 6783 27028 6792
rect 26976 6749 26985 6783
rect 26985 6749 27019 6783
rect 27019 6749 27028 6783
rect 26976 6740 27028 6749
rect 29276 6783 29328 6792
rect 29276 6749 29285 6783
rect 29285 6749 29319 6783
rect 29319 6749 29328 6783
rect 29276 6740 29328 6749
rect 30656 6740 30708 6792
rect 32404 6740 32456 6792
rect 14832 6672 14884 6724
rect 14924 6672 14976 6724
rect 4160 6604 4212 6656
rect 6736 6604 6788 6656
rect 9220 6604 9272 6656
rect 11612 6604 11664 6656
rect 13176 6604 13228 6656
rect 17592 6604 17644 6656
rect 20352 6604 20404 6656
rect 24400 6647 24452 6656
rect 24400 6613 24409 6647
rect 24409 6613 24443 6647
rect 24443 6613 24452 6647
rect 24400 6604 24452 6613
rect 24676 6647 24728 6656
rect 24676 6613 24685 6647
rect 24685 6613 24719 6647
rect 24719 6613 24728 6647
rect 24676 6604 24728 6613
rect 25044 6604 25096 6656
rect 25412 6647 25464 6656
rect 25412 6613 25421 6647
rect 25421 6613 25455 6647
rect 25455 6613 25464 6647
rect 25412 6604 25464 6613
rect 25504 6604 25556 6656
rect 26424 6604 26476 6656
rect 26608 6604 26660 6656
rect 28632 6604 28684 6656
rect 33416 6672 33468 6724
rect 32864 6647 32916 6656
rect 32864 6613 32873 6647
rect 32873 6613 32907 6647
rect 32907 6613 32916 6647
rect 32864 6604 32916 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 4896 6400 4948 6452
rect 5264 6400 5316 6452
rect 6460 6400 6512 6452
rect 7104 6400 7156 6452
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 7472 6443 7524 6452
rect 7472 6409 7481 6443
rect 7481 6409 7515 6443
rect 7515 6409 7524 6443
rect 7472 6400 7524 6409
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 7748 6400 7800 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 13728 6443 13780 6452
rect 13728 6409 13737 6443
rect 13737 6409 13771 6443
rect 13771 6409 13780 6443
rect 13728 6400 13780 6409
rect 14464 6400 14516 6452
rect 15200 6400 15252 6452
rect 17500 6400 17552 6452
rect 17592 6400 17644 6452
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 4804 6264 4856 6273
rect 12992 6332 13044 6384
rect 6644 6196 6696 6248
rect 5448 6128 5500 6180
rect 6276 6060 6328 6112
rect 7196 6264 7248 6316
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 9588 6264 9640 6316
rect 13912 6264 13964 6316
rect 12164 6196 12216 6248
rect 8300 6128 8352 6180
rect 14556 6264 14608 6316
rect 16580 6332 16632 6384
rect 17224 6332 17276 6384
rect 21916 6264 21968 6316
rect 22008 6307 22060 6316
rect 22008 6273 22025 6307
rect 22025 6273 22059 6307
rect 22059 6273 22060 6307
rect 22008 6264 22060 6273
rect 22284 6307 22336 6316
rect 22284 6273 22293 6307
rect 22293 6273 22327 6307
rect 22327 6273 22336 6307
rect 22284 6264 22336 6273
rect 11980 6060 12032 6112
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 12992 6103 13044 6112
rect 12992 6069 13001 6103
rect 13001 6069 13035 6103
rect 13035 6069 13044 6103
rect 12992 6060 13044 6069
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 13636 6128 13688 6180
rect 16304 6196 16356 6248
rect 16028 6128 16080 6180
rect 19800 6128 19852 6180
rect 13912 6060 13964 6112
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14004 6060 14056 6069
rect 14372 6060 14424 6112
rect 14740 6060 14792 6112
rect 14924 6060 14976 6112
rect 15660 6103 15712 6112
rect 15660 6069 15669 6103
rect 15669 6069 15703 6103
rect 15703 6069 15712 6103
rect 15660 6060 15712 6069
rect 17960 6060 18012 6112
rect 19432 6060 19484 6112
rect 20904 6060 20956 6112
rect 24216 6400 24268 6452
rect 24492 6400 24544 6452
rect 26424 6400 26476 6452
rect 32864 6443 32916 6452
rect 32864 6409 32873 6443
rect 32873 6409 32907 6443
rect 32907 6409 32916 6443
rect 32864 6400 32916 6409
rect 23848 6332 23900 6384
rect 23664 6264 23716 6316
rect 32312 6307 32364 6316
rect 32312 6273 32321 6307
rect 32321 6273 32355 6307
rect 32355 6273 32364 6307
rect 32312 6264 32364 6273
rect 24032 6196 24084 6248
rect 30472 6196 30524 6248
rect 22928 6171 22980 6180
rect 22928 6137 22937 6171
rect 22937 6137 22971 6171
rect 22971 6137 22980 6171
rect 22928 6128 22980 6137
rect 24308 6128 24360 6180
rect 23204 6103 23256 6112
rect 23204 6069 23213 6103
rect 23213 6069 23247 6103
rect 23247 6069 23256 6103
rect 23204 6060 23256 6069
rect 32496 6103 32548 6112
rect 32496 6069 32505 6103
rect 32505 6069 32539 6103
rect 32539 6069 32548 6103
rect 32496 6060 32548 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 4804 5856 4856 5908
rect 7380 5856 7432 5908
rect 8484 5856 8536 5908
rect 4528 5788 4580 5840
rect 12716 5856 12768 5908
rect 12900 5856 12952 5908
rect 17960 5856 18012 5908
rect 18052 5856 18104 5908
rect 23204 5856 23256 5908
rect 10968 5788 11020 5840
rect 13360 5788 13412 5840
rect 6920 5720 6972 5772
rect 7012 5652 7064 5704
rect 16488 5788 16540 5840
rect 19708 5788 19760 5840
rect 20352 5788 20404 5840
rect 32312 5856 32364 5908
rect 32864 5831 32916 5840
rect 32864 5797 32873 5831
rect 32873 5797 32907 5831
rect 32907 5797 32916 5831
rect 32864 5788 32916 5797
rect 14648 5720 14700 5772
rect 25412 5720 25464 5772
rect 3424 5584 3476 5636
rect 10692 5584 10744 5636
rect 12716 5584 12768 5636
rect 16580 5652 16632 5704
rect 16672 5695 16724 5704
rect 16672 5661 16681 5695
rect 16681 5661 16715 5695
rect 16715 5661 16724 5695
rect 16672 5652 16724 5661
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 20628 5652 20680 5704
rect 32404 5720 32456 5772
rect 27436 5652 27488 5704
rect 16488 5584 16540 5636
rect 13820 5516 13872 5568
rect 14556 5516 14608 5568
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 16580 5516 16632 5568
rect 16856 5559 16908 5568
rect 16856 5525 16865 5559
rect 16865 5525 16899 5559
rect 16899 5525 16908 5559
rect 16856 5516 16908 5525
rect 19800 5584 19852 5636
rect 30564 5584 30616 5636
rect 33416 5516 33468 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 12072 5312 12124 5364
rect 15752 5312 15804 5364
rect 15844 5312 15896 5364
rect 17408 5312 17460 5364
rect 17592 5312 17644 5364
rect 4712 5108 4764 5160
rect 16764 5108 16816 5160
rect 18144 5219 18196 5228
rect 18144 5185 18153 5219
rect 18153 5185 18187 5219
rect 18187 5185 18196 5219
rect 18144 5176 18196 5185
rect 32864 5355 32916 5364
rect 32864 5321 32873 5355
rect 32873 5321 32907 5355
rect 32907 5321 32916 5355
rect 32864 5312 32916 5321
rect 19708 5176 19760 5228
rect 32312 5219 32364 5228
rect 32312 5185 32321 5219
rect 32321 5185 32355 5219
rect 32355 5185 32364 5219
rect 32312 5176 32364 5185
rect 18788 5108 18840 5160
rect 30656 5108 30708 5160
rect 4068 5040 4120 5092
rect 14648 5040 14700 5092
rect 14924 5040 14976 5092
rect 18512 5040 18564 5092
rect 28908 5040 28960 5092
rect 14556 4972 14608 5024
rect 16948 5015 17000 5024
rect 16948 4981 16957 5015
rect 16957 4981 16991 5015
rect 16991 4981 17000 5015
rect 16948 4972 17000 4981
rect 17500 5015 17552 5024
rect 17500 4981 17509 5015
rect 17509 4981 17543 5015
rect 17543 4981 17552 5015
rect 17500 4972 17552 4981
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 18328 5015 18380 5024
rect 18328 4981 18337 5015
rect 18337 4981 18371 5015
rect 18371 4981 18380 5015
rect 18328 4972 18380 4981
rect 26792 4972 26844 5024
rect 31760 4972 31812 5024
rect 32496 5015 32548 5024
rect 32496 4981 32505 5015
rect 32505 4981 32539 5015
rect 32539 4981 32548 5015
rect 32496 4972 32548 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 11520 4768 11572 4820
rect 14648 4768 14700 4820
rect 17960 4768 18012 4820
rect 18328 4768 18380 4820
rect 26884 4768 26936 4820
rect 27620 4768 27672 4820
rect 2780 4700 2832 4752
rect 17868 4700 17920 4752
rect 18052 4700 18104 4752
rect 31668 4700 31720 4752
rect 32864 4743 32916 4752
rect 32864 4709 32873 4743
rect 32873 4709 32907 4743
rect 32907 4709 32916 4743
rect 32864 4700 32916 4709
rect 16580 4632 16632 4684
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 7840 4496 7892 4548
rect 16396 4564 16448 4616
rect 15752 4496 15804 4548
rect 20536 4496 20588 4548
rect 17132 4428 17184 4480
rect 18696 4428 18748 4480
rect 28908 4428 28960 4480
rect 32404 4428 32456 4480
rect 33416 4428 33468 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 12348 4224 12400 4276
rect 3424 4088 3476 4140
rect 10048 4088 10100 4140
rect 10324 3952 10376 4004
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 11796 4020 11848 4072
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 9772 3884 9824 3936
rect 13084 4224 13136 4276
rect 17500 4224 17552 4276
rect 26792 4224 26844 4276
rect 26884 4224 26936 4276
rect 14832 4156 14884 4208
rect 15384 4156 15436 4208
rect 16488 4088 16540 4140
rect 31668 4088 31720 4140
rect 16396 4020 16448 4072
rect 17224 4020 17276 4072
rect 22652 4020 22704 4072
rect 12624 3995 12676 4004
rect 12624 3961 12633 3995
rect 12633 3961 12667 3995
rect 12667 3961 12676 3995
rect 12624 3952 12676 3961
rect 32864 3995 32916 4004
rect 32864 3961 32873 3995
rect 32873 3961 32907 3995
rect 32907 3961 32916 3995
rect 32864 3952 32916 3961
rect 19340 3884 19392 3936
rect 21088 3884 21140 3936
rect 25320 3884 25372 3936
rect 32496 3927 32548 3936
rect 32496 3893 32505 3927
rect 32505 3893 32539 3927
rect 32539 3893 32548 3927
rect 32496 3884 32548 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 7288 3680 7340 3732
rect 8392 3680 8444 3732
rect 10508 3723 10560 3732
rect 10508 3689 10517 3723
rect 10517 3689 10551 3723
rect 10551 3689 10560 3723
rect 10508 3680 10560 3689
rect 11060 3680 11112 3732
rect 15108 3680 15160 3732
rect 15384 3723 15436 3732
rect 15384 3689 15393 3723
rect 15393 3689 15427 3723
rect 15427 3689 15436 3723
rect 15384 3680 15436 3689
rect 11704 3612 11756 3664
rect 15568 3612 15620 3664
rect 17224 3544 17276 3596
rect 17776 3655 17828 3664
rect 17776 3621 17785 3655
rect 17785 3621 17819 3655
rect 17819 3621 17828 3655
rect 17776 3612 17828 3621
rect 18788 3680 18840 3732
rect 19616 3680 19668 3732
rect 18420 3612 18472 3664
rect 20352 3680 20404 3732
rect 20628 3723 20680 3732
rect 20628 3689 20637 3723
rect 20637 3689 20671 3723
rect 20671 3689 20680 3723
rect 20628 3680 20680 3689
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 24860 3680 24912 3732
rect 27344 3680 27396 3732
rect 28356 3680 28408 3732
rect 27436 3612 27488 3664
rect 27988 3612 28040 3664
rect 32864 3655 32916 3664
rect 32864 3621 32873 3655
rect 32873 3621 32907 3655
rect 32907 3621 32916 3655
rect 32864 3612 32916 3621
rect 1492 3476 1544 3528
rect 4620 3408 4672 3460
rect 14188 3476 14240 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 16764 3476 16816 3528
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 17960 3476 18012 3528
rect 20444 3519 20496 3528
rect 20444 3485 20453 3519
rect 20453 3485 20487 3519
rect 20487 3485 20496 3519
rect 20444 3476 20496 3485
rect 16672 3408 16724 3460
rect 24860 3476 24912 3528
rect 15752 3383 15804 3392
rect 15752 3349 15761 3383
rect 15761 3349 15795 3383
rect 15795 3349 15804 3383
rect 15752 3340 15804 3349
rect 21364 3383 21416 3392
rect 21364 3349 21373 3383
rect 21373 3349 21407 3383
rect 21407 3349 21416 3383
rect 21364 3340 21416 3349
rect 27528 3408 27580 3460
rect 27620 3408 27672 3460
rect 30656 3476 30708 3528
rect 32404 3476 32456 3528
rect 22836 3383 22888 3392
rect 22836 3349 22845 3383
rect 22845 3349 22879 3383
rect 22879 3349 22888 3383
rect 22836 3340 22888 3349
rect 33416 3340 33468 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 12440 3136 12492 3188
rect 22836 3136 22888 3188
rect 32864 3179 32916 3188
rect 32864 3145 32873 3179
rect 32873 3145 32907 3179
rect 32907 3145 32916 3179
rect 32864 3136 32916 3145
rect 6184 3068 6236 3120
rect 14280 3068 14332 3120
rect 18512 3068 18564 3120
rect 31852 3068 31904 3120
rect 32036 3068 32088 3120
rect 14464 3000 14516 3052
rect 7748 2932 7800 2984
rect 21548 2932 21600 2984
rect 14372 2864 14424 2916
rect 30656 2932 30708 2984
rect 30380 2864 30432 2916
rect 15752 2796 15804 2848
rect 30564 2796 30616 2848
rect 31852 2839 31904 2848
rect 31852 2805 31861 2839
rect 31861 2805 31895 2839
rect 31895 2805 31904 2839
rect 31852 2796 31904 2805
rect 32496 2839 32548 2848
rect 32496 2805 32505 2839
rect 32505 2805 32539 2839
rect 32539 2805 32548 2839
rect 32496 2796 32548 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 16028 2592 16080 2644
rect 31300 2592 31352 2644
rect 16856 2524 16908 2576
rect 14740 2456 14792 2508
rect 32864 2567 32916 2576
rect 32864 2533 32873 2567
rect 32873 2533 32907 2567
rect 32907 2533 32916 2567
rect 32864 2524 32916 2533
rect 13728 2388 13780 2440
rect 3516 2320 3568 2372
rect 20444 2320 20496 2372
rect 31300 2431 31352 2440
rect 31300 2397 31309 2431
rect 31309 2397 31343 2431
rect 31343 2397 31352 2431
rect 31300 2388 31352 2397
rect 31760 2388 31812 2440
rect 20260 2252 20312 2304
rect 29276 2252 29328 2304
rect 31116 2295 31168 2304
rect 31116 2261 31125 2295
rect 31125 2261 31159 2295
rect 31159 2261 31168 2295
rect 31116 2252 31168 2261
rect 31484 2295 31536 2304
rect 31484 2261 31493 2295
rect 31493 2261 31527 2295
rect 31527 2261 31536 2295
rect 31484 2252 31536 2261
rect 31852 2295 31904 2304
rect 31852 2261 31861 2295
rect 31861 2261 31895 2295
rect 31895 2261 31904 2295
rect 31852 2252 31904 2261
rect 33416 2252 33468 2304
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 10876 2048 10928 2100
rect 21364 2048 21416 2100
rect 14096 8 14148 60
rect 24860 8 24912 60
<< metal2 >>
rect 5630 11096 5686 11152
rect 5814 11096 5870 11152
rect 5998 11096 6054 11152
rect 6182 11096 6238 11152
rect 6366 11096 6422 11152
rect 6550 11096 6606 11152
rect 6734 11096 6790 11152
rect 6918 11096 6974 11152
rect 7102 11096 7158 11152
rect 7286 11096 7342 11152
rect 7470 11096 7526 11152
rect 7564 11144 7616 11150
rect 5078 9616 5134 9625
rect 5078 9551 5134 9560
rect 1308 9376 1360 9382
rect 1308 9318 1360 9324
rect 1032 9308 1084 9314
rect 1032 9250 1084 9256
rect 296 9036 348 9042
rect 296 8978 348 8984
rect 308 7449 336 8978
rect 1044 8265 1072 9250
rect 1030 8256 1086 8265
rect 1030 8191 1086 8200
rect 1320 7721 1348 9318
rect 2870 9208 2926 9217
rect 2870 9143 2926 9152
rect 2884 8809 2912 9143
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 294 7440 350 7449
rect 2148 7410 2176 7958
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7546 2544 7686
rect 2792 7546 2820 7822
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 294 7375 350 7384
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3160 7206 3188 7346
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 3988 7002 4016 7346
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3514 6896 3570 6905
rect 3514 6831 3570 6840
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 2778 6624 2834 6633
rect 3344 6610 3372 6734
rect 3344 6582 3464 6610
rect 2778 6559 2834 6568
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2792 4758 2820 6559
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 3436 5642 3464 6582
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 2870 5536 2926 5545
rect 2870 5471 2926 5480
rect 2884 5250 2912 5471
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2962 5264 3018 5273
rect 2884 5222 2962 5250
rect 2962 5199 3018 5208
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2870 4720 2926 4729
rect 2870 4655 2926 4664
rect 2884 4570 2912 4655
rect 2884 4542 3372 4570
rect 3344 4434 3372 4542
rect 3422 4448 3478 4457
rect 3344 4406 3422 4434
rect 3010 4380 3318 4389
rect 3422 4383 3478 4392
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1504 56 1532 3470
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 3068 56 3188 82
rect 1490 0 1546 56
rect 3054 54 3188 56
rect 3054 0 3110 54
rect 3160 42 3188 54
rect 3436 42 3464 4082
rect 3528 2378 3556 6831
rect 4172 6662 4200 8298
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4356 6730 4384 7754
rect 4816 7342 4844 8434
rect 4804 7336 4856 7342
rect 5092 7313 5120 9551
rect 5354 9344 5410 9353
rect 5354 9279 5410 9288
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 4804 7278 4856 7284
rect 5078 7304 5134 7313
rect 5184 7274 5212 8434
rect 5078 7239 5134 7248
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4448 6730 4476 6870
rect 4894 6760 4950 6769
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4436 6724 4488 6730
rect 4894 6695 4950 6704
rect 4436 6666 4488 6672
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4908 6458 4936 6695
rect 5276 6458 5304 8434
rect 5368 7449 5396 9279
rect 5644 8634 5672 11096
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5354 7440 5410 7449
rect 5354 7375 5410 7384
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 4710 6352 4766 6361
rect 4528 6316 4580 6322
rect 4710 6287 4766 6296
rect 4804 6316 4856 6322
rect 4528 6258 4580 6264
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4080 5098 4108 6151
rect 4540 5846 4568 6258
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 4724 5166 4752 6287
rect 4804 6258 4856 6264
rect 4816 5914 4844 6258
rect 5460 6186 5488 8366
rect 5828 8090 5856 11096
rect 6012 8362 6040 11096
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 6196 8090 6224 11096
rect 6380 8566 6408 11096
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 5920 7546 5948 7822
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 6288 6118 6316 7822
rect 6472 6458 6500 8774
rect 6564 8090 6592 11096
rect 6748 8634 6776 11096
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6932 8090 6960 11096
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6656 6254 6684 7822
rect 6748 6662 6776 7822
rect 6826 6896 6882 6905
rect 6826 6831 6828 6840
rect 6880 6831 6882 6840
rect 6828 6802 6880 6808
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 6932 5778 6960 6734
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 7024 5710 7052 11018
rect 7116 7546 7144 11096
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7208 6458 7236 8842
rect 7300 8090 7328 11096
rect 7378 9480 7434 9489
rect 7378 9415 7434 9424
rect 7392 8537 7420 9415
rect 7484 8634 7512 11096
rect 7654 11096 7710 11152
rect 7838 11096 7894 11152
rect 8022 11096 8078 11152
rect 8206 11096 8262 11152
rect 8298 11112 8354 11121
rect 7564 11086 7616 11092
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7378 8528 7434 8537
rect 7378 8463 7434 8472
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7116 6304 7144 6394
rect 7196 6316 7248 6322
rect 7116 6276 7196 6304
rect 7392 6304 7420 8366
rect 7484 8265 7512 8434
rect 7576 8430 7604 11086
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7470 8256 7526 8265
rect 7470 8191 7526 8200
rect 7668 8090 7696 11096
rect 7852 9602 7880 11096
rect 7760 9574 7880 9602
rect 7760 8634 7788 9574
rect 8036 9466 8064 11096
rect 7852 9438 8064 9466
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7562 7984 7618 7993
rect 7472 7948 7524 7954
rect 7562 7919 7618 7928
rect 7472 7890 7524 7896
rect 7484 6458 7512 7890
rect 7576 6458 7604 7919
rect 7760 6458 7788 8298
rect 7852 8090 7880 9438
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 7944 8498 7972 8842
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 8498 8156 8774
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8220 8362 8248 11096
rect 8390 11096 8446 11152
rect 8574 11096 8630 11152
rect 8758 11096 8814 11152
rect 8942 11096 8998 11152
rect 9126 11096 9182 11152
rect 9310 11096 9366 11152
rect 9494 11096 9550 11152
rect 9678 11096 9734 11152
rect 9862 11096 9918 11152
rect 10046 11096 10102 11152
rect 10230 11096 10286 11152
rect 10414 11096 10470 11152
rect 10598 11096 10654 11152
rect 10782 11096 10838 11152
rect 10966 11096 11022 11152
rect 11150 11096 11206 11152
rect 11334 11096 11390 11152
rect 11518 11096 11574 11152
rect 11702 11096 11758 11152
rect 11886 11096 11942 11152
rect 12070 11096 12126 11152
rect 12254 11096 12310 11152
rect 12438 11096 12494 11152
rect 12622 11096 12678 11152
rect 12806 11096 12862 11152
rect 12990 11096 13046 11152
rect 13174 11096 13230 11152
rect 13358 11096 13414 11152
rect 13542 11096 13598 11152
rect 13726 11096 13782 11152
rect 13910 11096 13966 11152
rect 14094 11096 14150 11152
rect 14278 11096 14334 11152
rect 14462 11096 14518 11152
rect 14646 11096 14702 11152
rect 14830 11096 14886 11152
rect 15014 11096 15070 11152
rect 15198 11096 15254 11152
rect 15382 11096 15438 11152
rect 15566 11096 15622 11152
rect 15750 11096 15806 11152
rect 15934 11096 15990 11152
rect 16118 11096 16174 11152
rect 16302 11096 16358 11152
rect 16486 11096 16542 11152
rect 16670 11096 16726 11152
rect 16854 11096 16910 11152
rect 17038 11096 17094 11152
rect 17222 11096 17278 11152
rect 17406 11096 17462 11152
rect 17590 11096 17646 11152
rect 17774 11096 17830 11152
rect 17958 11096 18014 11152
rect 18052 11144 18104 11150
rect 8298 11047 8354 11056
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7248 6276 7420 6304
rect 7746 6352 7802 6361
rect 7746 6287 7748 6296
rect 7196 6258 7248 6264
rect 7800 6287 7802 6296
rect 7748 6258 7800 6264
rect 8312 6186 8340 11047
rect 8404 8090 8432 11096
rect 8482 9752 8538 9761
rect 8482 9687 8538 9696
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8496 8022 8524 9687
rect 8588 8566 8616 11096
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8680 8362 8708 9386
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8772 8090 8800 11096
rect 8956 8820 8984 11096
rect 9140 9194 9168 11096
rect 9324 9450 9352 11096
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9140 9166 9444 9194
rect 8864 8792 8984 8820
rect 8864 8634 8892 8792
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 6458 8432 7754
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 8496 5914 8524 7822
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9416 7546 9444 9166
rect 9508 8090 9536 11096
rect 9588 10872 9640 10878
rect 9588 10814 9640 10820
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9232 6662 9260 7346
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9600 6322 9628 10814
rect 9692 7546 9720 11096
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 7392 5817 7420 5850
rect 7378 5808 7434 5817
rect 7378 5743 7434 5752
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 8482 5128 8538 5137
rect 4068 5092 4120 5098
rect 8482 5063 8538 5072
rect 4068 5034 4120 5040
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 8496 4729 8524 5063
rect 8482 4720 8538 4729
rect 8482 4655 8538 4664
rect 8666 4720 8722 4729
rect 8666 4655 8722 4664
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7300 3505 7328 3674
rect 7286 3496 7342 3505
rect 4620 3460 4672 3466
rect 7286 3431 7342 3440
rect 4620 3402 4672 3408
rect 3516 2372 3568 2378
rect 3516 2314 3568 2320
rect 4632 56 4660 3402
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 6196 56 6224 3062
rect 7760 2990 7788 3878
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7852 2774 7880 4490
rect 8680 4457 8708 4655
rect 8666 4448 8722 4457
rect 8666 4383 8722 4392
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9784 3942 9812 8434
rect 9876 8090 9904 11096
rect 9954 9888 10010 9897
rect 9954 9823 10010 9832
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9968 6866 9996 9823
rect 10060 8634 10088 11096
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10152 8514 10180 8842
rect 10060 8486 10180 8514
rect 10060 8294 10088 8486
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10244 8090 10272 11096
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10336 8566 10364 8910
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 10060 4146 10088 7754
rect 10244 7274 10272 7822
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10336 4010 10364 8366
rect 10428 8362 10456 11096
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8634 10548 8774
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10506 8528 10562 8537
rect 10506 8463 10562 8472
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 8390 3768 8446 3777
rect 10520 3738 10548 8463
rect 10612 8090 10640 11096
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10598 7984 10654 7993
rect 10598 7919 10654 7928
rect 10612 7750 10640 7919
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10704 5642 10732 10610
rect 10796 8906 10824 11096
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10796 7585 10824 8434
rect 10782 7576 10838 7585
rect 10782 7511 10838 7520
rect 10888 7206 10916 8842
rect 10980 8090 11008 11096
rect 11164 8838 11192 11096
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10980 7750 11008 7822
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 11072 7478 11100 8570
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 7546 11192 8230
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 10980 7206 11008 7346
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 8390 3703 8392 3712
rect 8444 3703 8446 3712
rect 10508 3732 10560 3738
rect 8392 3674 8444 3680
rect 10508 3674 10560 3680
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 9402 2952 9458 2961
rect 9402 2887 9458 2896
rect 7760 2746 7880 2774
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 7760 56 7788 2746
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9416 1442 9444 2887
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 9324 1414 9444 1442
rect 9324 56 9352 1414
rect 10888 56 10916 2042
rect 10980 1193 11008 5782
rect 11072 3738 11100 7210
rect 11164 6934 11192 7346
rect 11256 7274 11284 8434
rect 11348 8090 11376 11096
rect 11426 10024 11482 10033
rect 11426 9959 11482 9968
rect 11440 8294 11468 9959
rect 11532 8362 11560 11096
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11440 4298 11468 7958
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11532 4826 11560 7890
rect 11624 6662 11652 8434
rect 11716 8090 11744 11096
rect 11900 8634 11928 11096
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11888 8016 11940 8022
rect 11888 7958 11940 7964
rect 11992 7970 12020 10474
rect 12084 8090 12112 11096
rect 12162 10160 12218 10169
rect 12162 10095 12218 10104
rect 12176 8906 12204 10095
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12162 8664 12218 8673
rect 12162 8599 12218 8608
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11716 7002 11744 7822
rect 11808 7546 11836 7822
rect 11900 7546 11928 7958
rect 11992 7942 12112 7970
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 12084 7426 12112 7942
rect 11992 7398 12112 7426
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11992 6118 12020 7398
rect 12176 6254 12204 8599
rect 12268 8090 12296 11096
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12360 8634 12388 8842
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12452 8090 12480 11096
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12544 7834 12572 8910
rect 12636 8294 12664 11096
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12728 8566 12756 8774
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12820 8090 12848 11096
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12912 8498 12940 8910
rect 13004 8906 13032 11096
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 12990 8800 13046 8809
rect 12990 8735 13046 8744
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 13004 8378 13032 8735
rect 13004 8350 13124 8378
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12808 7880 12860 7886
rect 12544 7806 12664 7834
rect 12808 7822 12860 7828
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12544 7546 12572 7686
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12440 7268 12492 7274
rect 12440 7210 12492 7216
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 12084 4622 12112 5306
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 11440 4270 11836 4298
rect 12360 4282 12388 7142
rect 12452 7002 12480 7210
rect 12544 7206 12572 7346
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11716 3670 11744 4082
rect 11808 4078 11836 4270
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11992 3505 12020 4082
rect 12636 4010 12664 7806
rect 12714 7576 12770 7585
rect 12714 7511 12716 7520
rect 12768 7511 12770 7520
rect 12716 7482 12768 7488
rect 12820 7342 12848 7822
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12728 5642 12756 5850
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12820 3777 12848 6054
rect 12912 5914 12940 6802
rect 13004 6390 13032 6802
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12806 3768 12862 3777
rect 12806 3703 12862 3712
rect 11978 3496 12034 3505
rect 11978 3431 12034 3440
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 10966 1184 11022 1193
rect 10966 1119 11022 1128
rect 12452 56 12480 3130
rect 13004 2009 13032 6054
rect 13096 4282 13124 8350
rect 13188 8090 13216 11096
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13188 6662 13216 7822
rect 13280 7206 13308 10134
rect 13372 8634 13400 11096
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13464 8498 13492 9454
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13556 8090 13584 11096
rect 13636 9784 13688 9790
rect 13636 9726 13688 9732
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13360 7812 13412 7818
rect 13360 7754 13412 7760
rect 13372 7546 13400 7754
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13648 6798 13676 9726
rect 13740 8430 13768 11096
rect 13820 9240 13872 9246
rect 13820 9182 13872 9188
rect 13832 8498 13860 9182
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13728 8424 13780 8430
rect 13924 8378 13952 11096
rect 14002 10296 14058 10305
rect 14002 10231 14058 10240
rect 14016 8673 14044 10231
rect 14002 8664 14058 8673
rect 14108 8634 14136 11096
rect 14002 8599 14058 8608
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13728 8366 13780 8372
rect 13832 8362 13952 8378
rect 13820 8356 13952 8362
rect 13872 8350 13952 8356
rect 13820 8298 13872 8304
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14292 8090 14320 11096
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14384 7993 14412 10542
rect 14476 8634 14504 11096
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14568 8498 14596 8774
rect 14660 8634 14688 11096
rect 14738 9072 14794 9081
rect 14738 9007 14794 9016
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14370 7984 14426 7993
rect 14370 7919 14426 7928
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14568 6798 14596 8230
rect 14752 7993 14780 9007
rect 14844 8362 14872 11096
rect 15028 8888 15056 11096
rect 15212 9058 15240 11096
rect 15396 10169 15424 11096
rect 15382 10160 15438 10169
rect 15382 10095 15438 10104
rect 15580 10033 15608 11096
rect 15764 10606 15792 11096
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15566 10024 15622 10033
rect 15566 9959 15622 9968
rect 15948 9761 15976 11096
rect 16132 10674 16160 11096
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16316 9897 16344 11096
rect 16302 9888 16358 9897
rect 16302 9823 16358 9832
rect 15934 9752 15990 9761
rect 15934 9687 15990 9696
rect 15566 9616 15622 9625
rect 15566 9551 15622 9560
rect 15660 9580 15712 9586
rect 15212 9030 15424 9058
rect 14936 8860 15056 8888
rect 14936 8634 14964 8860
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14738 7984 14794 7993
rect 14738 7919 14794 7928
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13188 4729 13216 6054
rect 13372 5846 13400 6054
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13174 4720 13230 4729
rect 13174 4655 13230 4664
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12990 2000 13046 2009
rect 12990 1935 13046 1944
rect 13648 1737 13676 6122
rect 13740 2446 13768 6394
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13924 6118 13952 6258
rect 14002 6216 14058 6225
rect 14002 6151 14058 6160
rect 14016 6118 14044 6151
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 4865 13860 5510
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13818 4856 13874 4865
rect 13950 4859 14258 4868
rect 13818 4791 13874 4800
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 14188 3528 14240 3534
rect 14002 3496 14058 3505
rect 14002 3431 14058 3440
rect 14186 3496 14188 3505
rect 14280 3528 14332 3534
rect 14240 3496 14242 3505
rect 14280 3470 14332 3476
rect 14186 3431 14242 3440
rect 14016 3346 14044 3431
rect 14016 3318 14228 3346
rect 14200 2938 14228 3318
rect 14292 3126 14320 3470
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14200 2910 14320 2938
rect 14384 2922 14412 6054
rect 14476 3058 14504 6394
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14568 5574 14596 6258
rect 14660 5778 14688 7822
rect 14936 6730 14964 8434
rect 15396 8362 15424 9030
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15580 7002 15608 9551
rect 15660 9522 15712 9528
rect 15672 8498 15700 9522
rect 16394 9208 16450 9217
rect 16394 9143 16450 9152
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16224 7410 16252 8230
rect 16408 7546 16436 9143
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 14844 6338 14872 6666
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15212 6338 15240 6394
rect 14844 6310 15240 6338
rect 16316 6254 16344 7482
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16394 6216 16450 6225
rect 16028 6180 16080 6186
rect 16394 6151 16450 6160
rect 16028 6122 16080 6128
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14568 3369 14596 4966
rect 14660 4826 14688 5034
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14554 3360 14610 3369
rect 14554 3295 14610 3304
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14292 2802 14320 2910
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 14370 2816 14426 2825
rect 14292 2774 14370 2802
rect 13950 2748 14258 2757
rect 14370 2751 14426 2760
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 14752 2514 14780 6054
rect 14830 5672 14886 5681
rect 14830 5607 14886 5616
rect 14844 4214 14872 5607
rect 14936 5250 14964 6054
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 14936 5222 15056 5250
rect 14924 5092 14976 5098
rect 14924 5034 14976 5040
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14936 4049 14964 5034
rect 15028 4729 15056 5222
rect 15014 4720 15070 4729
rect 15014 4655 15070 4664
rect 15488 4593 15516 5510
rect 15474 4584 15530 4593
rect 15474 4519 15530 4528
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 14922 4040 14978 4049
rect 14922 3975 14978 3984
rect 15106 4040 15162 4049
rect 15106 3975 15162 3984
rect 15120 3738 15148 3975
rect 15396 3738 15424 4150
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 13634 1728 13690 1737
rect 13634 1663 13690 1672
rect 14016 66 14136 82
rect 14016 60 14148 66
rect 14016 56 14096 60
rect 3160 14 3464 42
rect 4618 0 4674 56
rect 6182 0 6238 56
rect 7746 0 7802 56
rect 9310 0 9366 56
rect 10874 0 10930 56
rect 12438 0 12494 56
rect 14002 54 14096 56
rect 14002 0 14058 54
rect 15580 56 15608 3606
rect 15672 1465 15700 6054
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15764 4554 15792 5306
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15764 2854 15792 3334
rect 15856 3097 15884 5306
rect 15842 3088 15898 3097
rect 15842 3023 15898 3032
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 16040 2650 16068 6122
rect 16408 4622 16436 6151
rect 16500 5846 16528 11096
rect 16684 10146 16712 11096
rect 16684 10118 16804 10146
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16578 7848 16634 7857
rect 16578 7783 16634 7792
rect 16592 7546 16620 7783
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16684 7478 16712 9930
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16776 6905 16804 10118
rect 16868 8922 16896 11096
rect 16868 8894 16988 8922
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16868 7274 16896 7686
rect 16856 7268 16908 7274
rect 16856 7210 16908 7216
rect 16762 6896 16818 6905
rect 16762 6831 16818 6840
rect 16960 6769 16988 8894
rect 17052 6866 17080 11096
rect 17130 9208 17186 9217
rect 17130 9143 17186 9152
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 16946 6760 17002 6769
rect 16946 6695 17002 6704
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16592 5710 16620 6326
rect 16580 5704 16632 5710
rect 16672 5704 16724 5710
rect 16580 5646 16632 5652
rect 16670 5672 16672 5681
rect 16724 5672 16726 5681
rect 16488 5636 16540 5642
rect 16670 5607 16726 5616
rect 16488 5578 16540 5584
rect 16500 5137 16528 5578
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16486 5128 16542 5137
rect 16486 5063 16542 5072
rect 16592 4690 16620 5510
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16408 3097 16436 4014
rect 16500 3505 16528 4082
rect 16776 3534 16804 5102
rect 16764 3528 16816 3534
rect 16486 3496 16542 3505
rect 16764 3470 16816 3476
rect 16486 3431 16542 3440
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16394 3088 16450 3097
rect 16394 3023 16450 3032
rect 16684 2961 16712 3402
rect 16670 2952 16726 2961
rect 16670 2887 16726 2896
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 16868 2582 16896 5510
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 16960 2417 16988 4966
rect 17144 4486 17172 9143
rect 17236 6390 17264 11096
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17420 5817 17448 11096
rect 17604 8922 17632 11096
rect 17788 10538 17816 11096
rect 17972 11014 18000 11096
rect 18142 11098 18198 11152
rect 18104 11096 18198 11098
rect 18326 11112 18382 11152
rect 18104 11092 18184 11096
rect 18052 11086 18184 11092
rect 18064 11070 18184 11086
rect 18510 11096 18566 11152
rect 18694 11096 18750 11152
rect 18878 11096 18934 11152
rect 19062 11096 19118 11152
rect 19246 11096 19302 11152
rect 19430 11096 19486 11152
rect 19614 11096 19670 11152
rect 19798 11096 19854 11152
rect 19982 11096 20038 11152
rect 20166 11096 20222 11152
rect 20350 11096 20406 11152
rect 20534 11096 20590 11152
rect 20718 11096 20774 11152
rect 20902 11096 20958 11152
rect 21086 11096 21142 11152
rect 21270 11096 21326 11152
rect 21454 11096 21510 11152
rect 21638 11096 21694 11152
rect 21822 11096 21878 11152
rect 22006 11096 22062 11152
rect 22190 11096 22246 11152
rect 22374 11096 22430 11152
rect 22558 11096 22614 11152
rect 22742 11096 22798 11152
rect 22926 11096 22982 11152
rect 23110 11096 23166 11152
rect 23294 11096 23350 11152
rect 23478 11096 23534 11152
rect 23662 11096 23718 11152
rect 23846 11096 23902 11152
rect 24030 11096 24086 11152
rect 24214 11096 24270 11152
rect 24398 11096 24454 11152
rect 24582 11096 24638 11152
rect 24766 11096 24822 11152
rect 24950 11096 25006 11152
rect 25134 11096 25190 11152
rect 25318 11096 25374 11152
rect 25502 11096 25558 11152
rect 25686 11096 25742 11152
rect 25870 11096 25926 11152
rect 26054 11096 26110 11152
rect 26238 11096 26294 11152
rect 26422 11096 26478 11152
rect 26606 11096 26662 11152
rect 26790 11096 26846 11152
rect 26974 11096 27030 11152
rect 27158 11096 27214 11152
rect 27342 11096 27398 11152
rect 27526 11096 27582 11152
rect 27710 11096 27766 11152
rect 27894 11096 27950 11152
rect 28078 11096 28134 11152
rect 28262 11096 28318 11152
rect 28446 11096 28502 11152
rect 28630 11096 28686 11152
rect 18326 11047 18382 11056
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 18524 10305 18552 11096
rect 18708 10878 18736 11096
rect 18696 10872 18748 10878
rect 18696 10814 18748 10820
rect 18510 10296 18566 10305
rect 18510 10231 18566 10240
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 17774 9480 17830 9489
rect 17774 9415 17830 9424
rect 17512 8894 17632 8922
rect 17512 6458 17540 8894
rect 17788 7206 17816 9415
rect 17958 9344 18014 9353
rect 17958 9279 18014 9288
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17880 7546 17908 7958
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17972 7274 18000 9279
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17604 6458 17632 6598
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17972 5914 18000 6054
rect 18064 5914 18092 8910
rect 18142 7304 18198 7313
rect 18142 7239 18144 7248
rect 18196 7239 18198 7248
rect 18144 7210 18196 7216
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17406 5808 17462 5817
rect 17406 5743 17462 5752
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17420 5370 17448 5646
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17512 4282 17540 4966
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17236 3602 17264 4014
rect 17604 3641 17632 5306
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17868 4752 17920 4758
rect 17868 4694 17920 4700
rect 17776 3664 17828 3670
rect 17590 3632 17646 3641
rect 17224 3596 17276 3602
rect 17590 3567 17646 3576
rect 17774 3632 17776 3641
rect 17828 3632 17830 3641
rect 17774 3567 17830 3576
rect 17224 3538 17276 3544
rect 17880 3534 17908 4694
rect 17972 3534 18000 4762
rect 18064 4758 18092 4966
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 18156 4185 18184 5170
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18340 4826 18368 4966
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18142 4176 18198 4185
rect 18142 4111 18198 4120
rect 18432 3670 18460 9590
rect 18602 7984 18658 7993
rect 18512 7948 18564 7954
rect 18602 7919 18658 7928
rect 18512 7890 18564 7896
rect 18524 7546 18552 7890
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18616 7410 18644 7919
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18892 6361 18920 11096
rect 19076 6934 19104 11096
rect 19260 9790 19288 11096
rect 19248 9784 19300 9790
rect 19248 9726 19300 9732
rect 19338 7576 19394 7585
rect 19338 7511 19394 7520
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 18878 6352 18934 6361
rect 18878 6287 18934 6296
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18524 3126 18552 5034
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18512 3120 18564 3126
rect 18512 3062 18564 3068
rect 16946 2408 17002 2417
rect 16946 2343 17002 2352
rect 17130 2000 17186 2009
rect 17130 1935 17186 1944
rect 15658 1456 15714 1465
rect 15658 1391 15714 1400
rect 17144 56 17172 1935
rect 18708 56 18736 4422
rect 18800 3738 18828 5102
rect 19352 3942 19380 7511
rect 19444 6118 19472 11096
rect 19628 9625 19656 11096
rect 19812 10198 19840 11096
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19614 9616 19670 9625
rect 19614 9551 19670 9560
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19536 7546 19564 9386
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19616 9308 19668 9314
rect 19616 9250 19668 9256
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19628 7410 19656 9250
rect 19720 7410 19748 9318
rect 19800 9308 19852 9314
rect 19800 9250 19852 9256
rect 19812 7546 19840 9250
rect 19996 8294 20024 11096
rect 20180 9994 20208 11096
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20364 8072 20392 11096
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20272 8044 20392 8072
rect 20272 7750 20300 8044
rect 20352 7812 20404 7818
rect 20352 7754 20404 7760
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19812 6186 19840 7278
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 20364 6662 20392 7754
rect 20456 7410 20484 8978
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 19800 6180 19852 6186
rect 19800 6122 19852 6128
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 19708 5840 19760 5846
rect 19708 5782 19760 5788
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 19614 5264 19670 5273
rect 19720 5234 19748 5782
rect 19800 5636 19852 5642
rect 19800 5578 19852 5584
rect 19614 5199 19670 5208
rect 19708 5228 19760 5234
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19628 3738 19656 5199
rect 19708 5170 19760 5176
rect 19812 5137 19840 5578
rect 19798 5128 19854 5137
rect 19798 5063 19854 5072
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20364 3738 20392 5782
rect 20548 4554 20576 11096
rect 20732 9654 20760 11096
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20916 9194 20944 11096
rect 20640 9166 20944 9194
rect 21100 9178 21128 11096
rect 21088 9172 21140 9178
rect 20640 7426 20668 9166
rect 21088 9114 21140 9120
rect 21284 9058 21312 11096
rect 20824 9030 21312 9058
rect 20718 8392 20774 8401
rect 20718 8327 20774 8336
rect 20732 7546 20760 8327
rect 20824 7585 20852 9030
rect 20904 8900 20956 8906
rect 20904 8842 20956 8848
rect 21364 8900 21416 8906
rect 21364 8842 21416 8848
rect 20810 7576 20866 7585
rect 20720 7540 20772 7546
rect 20810 7511 20866 7520
rect 20720 7482 20772 7488
rect 20640 7398 20760 7426
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20640 3738 20668 5646
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 20456 2378 20484 3470
rect 20732 3369 20760 7398
rect 20916 6118 20944 8842
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21272 7540 21324 7546
rect 21376 7528 21404 8842
rect 21324 7500 21404 7528
rect 21272 7482 21324 7488
rect 21178 7440 21234 7449
rect 21178 7375 21180 7384
rect 21232 7375 21234 7384
rect 21180 7346 21232 7352
rect 21192 7206 21220 7346
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21100 3738 21128 3878
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 21468 3505 21496 11096
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21454 3496 21510 3505
rect 21454 3431 21510 3440
rect 21364 3392 21416 3398
rect 20718 3360 20774 3369
rect 21364 3334 21416 3340
rect 20718 3295 20774 3304
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 20444 2372 20496 2378
rect 20444 2314 20496 2320
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 20272 56 20300 2246
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 21376 2106 21404 3334
rect 21560 2990 21588 7482
rect 21652 3097 21680 11096
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 21638 3088 21694 3097
rect 21638 3023 21694 3032
rect 21548 2984 21600 2990
rect 21744 2961 21772 9114
rect 21836 8945 21864 11096
rect 22020 9194 22048 11096
rect 21928 9166 22048 9194
rect 21822 8936 21878 8945
rect 21822 8871 21878 8880
rect 21928 7313 21956 9166
rect 22006 8936 22062 8945
rect 22006 8871 22062 8880
rect 21914 7304 21970 7313
rect 21914 7239 21970 7248
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21928 6322 21956 6734
rect 22020 6322 22048 8871
rect 22204 7750 22232 11096
rect 22282 9752 22338 9761
rect 22282 9687 22338 9696
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22296 6322 22324 9687
rect 22388 6905 22416 11096
rect 22572 8809 22600 11096
rect 22756 8974 22784 11096
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22558 8800 22614 8809
rect 22558 8735 22614 8744
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 22374 6896 22430 6905
rect 22374 6831 22430 6840
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 21822 5672 21878 5681
rect 21822 5607 21878 5616
rect 21548 2926 21600 2932
rect 21730 2952 21786 2961
rect 21730 2887 21786 2896
rect 21364 2100 21416 2106
rect 21364 2042 21416 2048
rect 21836 56 21864 5607
rect 22664 4078 22692 8366
rect 22940 8362 22968 11096
rect 22928 8356 22980 8362
rect 22928 8298 22980 8304
rect 22928 8084 22980 8090
rect 22928 8026 22980 8032
rect 22940 6186 22968 8026
rect 23124 6934 23152 11096
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 23308 6866 23336 11096
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23492 6798 23520 11096
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23676 6322 23704 11096
rect 23860 6390 23888 11096
rect 23848 6384 23900 6390
rect 23848 6326 23900 6332
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 24044 6254 24072 11096
rect 24228 6458 24256 11096
rect 24412 9602 24440 11096
rect 24320 9574 24440 9602
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24032 6248 24084 6254
rect 24032 6190 24084 6196
rect 24320 6186 24348 9574
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24412 6662 24440 9454
rect 24596 8945 24624 11096
rect 24780 9761 24808 11096
rect 24766 9752 24822 9761
rect 24766 9687 24822 9696
rect 24676 9240 24728 9246
rect 24676 9182 24728 9188
rect 24582 8936 24638 8945
rect 24582 8871 24638 8880
rect 24582 8800 24638 8809
rect 24582 8735 24638 8744
rect 24492 8492 24544 8498
rect 24492 8434 24544 8440
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24504 6458 24532 8434
rect 24596 7002 24624 8735
rect 24584 6996 24636 7002
rect 24584 6938 24636 6944
rect 24688 6662 24716 9182
rect 24964 8634 24992 11096
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24780 7410 24808 8230
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 22928 6180 22980 6186
rect 22928 6122 22980 6128
rect 24308 6180 24360 6186
rect 24308 6122 24360 6128
rect 23204 6112 23256 6118
rect 23204 6054 23256 6060
rect 23216 5914 23244 6054
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 23386 5128 23442 5137
rect 23386 5063 23442 5072
rect 22652 4072 22704 4078
rect 22652 4014 22704 4020
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 3194 22876 3334
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 23400 56 23428 5063
rect 24872 3738 24900 7754
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24872 66 24900 3470
rect 24860 60 24912 66
rect 14096 2 14148 8
rect 15566 0 15622 56
rect 17130 0 17186 56
rect 18694 0 18750 56
rect 20258 0 20314 56
rect 21822 0 21878 56
rect 23386 0 23442 56
rect 24964 56 24992 7346
rect 25056 6662 25084 8774
rect 25148 8634 25176 11096
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25134 8528 25190 8537
rect 25134 8463 25136 8472
rect 25188 8463 25190 8472
rect 25228 8492 25280 8498
rect 25136 8434 25188 8440
rect 25228 8434 25280 8440
rect 25136 8356 25188 8362
rect 25136 8298 25188 8304
rect 25148 6798 25176 8298
rect 25240 7546 25268 8434
rect 25332 8362 25360 11096
rect 25516 8634 25544 11096
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25504 8492 25556 8498
rect 25504 8434 25556 8440
rect 25320 8356 25372 8362
rect 25320 8298 25372 8304
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25332 3942 25360 7822
rect 25516 6662 25544 8434
rect 25608 6798 25636 8910
rect 25700 8566 25728 11096
rect 25688 8560 25740 8566
rect 25688 8502 25740 8508
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 25412 6656 25464 6662
rect 25412 6598 25464 6604
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 25424 5778 25452 6598
rect 25412 5772 25464 5778
rect 25412 5714 25464 5720
rect 25792 4049 25820 8434
rect 25884 8090 25912 11096
rect 26068 8362 26096 11096
rect 26252 8514 26280 11096
rect 26436 9602 26464 11096
rect 26436 9574 26556 9602
rect 26422 9208 26478 9217
rect 26422 9143 26478 9152
rect 26252 8486 26372 8514
rect 26436 8498 26464 9143
rect 26056 8356 26108 8362
rect 26056 8298 26108 8304
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 26344 8090 26372 8486
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 26528 8430 26556 9574
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 26620 8090 26648 11096
rect 26700 9580 26752 9586
rect 26700 9522 26752 9528
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 26332 8084 26384 8090
rect 26332 8026 26384 8032
rect 26608 8084 26660 8090
rect 26608 8026 26660 8032
rect 26712 7834 26740 9522
rect 26804 8634 26832 11096
rect 26988 9160 27016 11096
rect 26896 9132 27016 9160
rect 26792 8628 26844 8634
rect 26792 8570 26844 8576
rect 26896 8090 26924 9132
rect 27172 8838 27200 11096
rect 27160 8832 27212 8838
rect 27160 8774 27212 8780
rect 27356 8786 27384 11096
rect 27540 8974 27568 11096
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27528 8832 27580 8838
rect 27356 8758 27476 8786
rect 27528 8774 27580 8780
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 26884 8084 26936 8090
rect 26884 8026 26936 8032
rect 26620 7806 26740 7834
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 26514 7032 26570 7041
rect 26514 6967 26570 6976
rect 26330 6896 26386 6905
rect 26330 6831 26386 6840
rect 26344 6798 26372 6831
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 26436 6458 26464 6598
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25778 4040 25834 4049
rect 25778 3975 25834 3984
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26528 56 26556 6967
rect 26620 6662 26648 7806
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 26712 6798 26740 7686
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26974 7304 27030 7313
rect 26804 6934 26832 7278
rect 26884 7268 26936 7274
rect 26974 7239 27030 7248
rect 26884 7210 26936 7216
rect 26896 7002 26924 7210
rect 26884 6996 26936 7002
rect 26884 6938 26936 6944
rect 26792 6928 26844 6934
rect 26792 6870 26844 6876
rect 26988 6798 27016 7239
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 26792 5024 26844 5030
rect 26792 4966 26844 4972
rect 26804 4282 26832 4966
rect 26884 4820 26936 4826
rect 26884 4762 26936 4768
rect 26896 4282 26924 4762
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 26792 4276 26844 4282
rect 26792 4218 26844 4224
rect 26884 4276 26936 4282
rect 26884 4218 26936 4224
rect 27356 3738 27384 8434
rect 27448 8090 27476 8758
rect 27540 8566 27568 8774
rect 27528 8560 27580 8566
rect 27528 8502 27580 8508
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 27632 8378 27660 8434
rect 27540 8350 27660 8378
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 27448 3670 27476 5646
rect 27436 3664 27488 3670
rect 27436 3606 27488 3612
rect 27540 3466 27568 8350
rect 27724 8090 27752 11096
rect 27908 8362 27936 11096
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 27896 8356 27948 8362
rect 27896 8298 27948 8304
rect 27712 8084 27764 8090
rect 27712 8026 27764 8032
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27632 4826 27660 7822
rect 27724 7274 27752 7822
rect 27816 7546 27844 7822
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 27712 7268 27764 7274
rect 27712 7210 27764 7216
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 28000 3670 28028 8434
rect 28092 8090 28120 11096
rect 28080 8084 28132 8090
rect 28276 8072 28304 11096
rect 28356 8084 28408 8090
rect 28276 8044 28356 8072
rect 28080 8026 28132 8032
rect 28356 8026 28408 8032
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 28080 7404 28132 7410
rect 28080 7346 28132 7352
rect 28092 5137 28120 7346
rect 28078 5128 28134 5137
rect 28078 5063 28134 5072
rect 28368 3738 28396 7754
rect 28460 7750 28488 11096
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 28552 8634 28580 8910
rect 28644 8634 28672 11096
rect 31758 9616 31814 9625
rect 31758 9551 31814 9560
rect 31668 9444 31720 9450
rect 31668 9386 31720 9392
rect 31298 9344 31354 9353
rect 31298 9279 31354 9288
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 31312 8498 31340 9279
rect 31482 8936 31538 8945
rect 31482 8871 31538 8880
rect 31496 8634 31524 8871
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31680 8498 31708 9386
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28448 7404 28500 7410
rect 28448 7346 28500 7352
rect 28460 5681 28488 7346
rect 28644 6662 28672 8434
rect 28736 7546 28764 8434
rect 28816 7880 28868 7886
rect 28816 7822 28868 7828
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 28828 7274 28856 7822
rect 28920 7546 28948 8434
rect 29092 7812 29144 7818
rect 29092 7754 29144 7760
rect 29104 7546 29132 7754
rect 29840 7546 29868 8434
rect 31668 8288 31720 8294
rect 31668 8230 31720 8236
rect 31680 7886 31708 8230
rect 31772 8090 31800 9551
rect 32586 9344 32642 9353
rect 32312 9308 32364 9314
rect 32586 9279 32642 9288
rect 32312 9250 32364 9256
rect 31852 8628 31904 8634
rect 31852 8570 31904 8576
rect 31864 8537 31892 8570
rect 31850 8528 31906 8537
rect 32324 8498 32352 9250
rect 31850 8463 31906 8472
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32496 8356 32548 8362
rect 32496 8298 32548 8304
rect 32508 8265 32536 8298
rect 32494 8256 32550 8265
rect 31950 8188 32258 8197
rect 32494 8191 32550 8200
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 32404 7948 32456 7954
rect 32404 7890 32456 7896
rect 30656 7880 30708 7886
rect 30656 7822 30708 7828
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 32312 7880 32364 7886
rect 32312 7822 32364 7828
rect 30668 7546 30696 7822
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 29092 7540 29144 7546
rect 29092 7482 29144 7488
rect 29828 7540 29880 7546
rect 29828 7482 29880 7488
rect 30656 7540 30708 7546
rect 30656 7482 30708 7488
rect 29092 7404 29144 7410
rect 29092 7346 29144 7352
rect 29368 7404 29420 7410
rect 29368 7346 29420 7352
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 28816 7268 28868 7274
rect 28816 7210 28868 7216
rect 29104 7041 29132 7346
rect 29090 7032 29146 7041
rect 29090 6967 29146 6976
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 28632 6656 28684 6662
rect 28632 6598 28684 6604
rect 28446 5672 28502 5681
rect 28446 5607 28502 5616
rect 28908 5092 28960 5098
rect 28908 5034 28960 5040
rect 28920 4486 28948 5034
rect 28908 4480 28960 4486
rect 28908 4422 28960 4428
rect 28356 3732 28408 3738
rect 28356 3674 28408 3680
rect 27988 3664 28040 3670
rect 27988 3606 28040 3612
rect 27528 3460 27580 3466
rect 27528 3402 27580 3408
rect 27620 3460 27672 3466
rect 27620 3402 27672 3408
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27632 2009 27660 3402
rect 28078 2680 28134 2689
rect 28078 2615 28134 2624
rect 27618 2000 27674 2009
rect 27618 1935 27674 1944
rect 28092 56 28120 2615
rect 29288 2310 29316 6734
rect 29380 2689 29408 7346
rect 29644 7336 29696 7342
rect 29644 7278 29696 7284
rect 29366 2680 29422 2689
rect 29366 2615 29422 2624
rect 29276 2304 29328 2310
rect 29276 2246 29328 2252
rect 29656 56 29684 7278
rect 30196 7200 30248 7206
rect 30196 7142 30248 7148
rect 30208 6934 30236 7142
rect 30196 6928 30248 6934
rect 30196 6870 30248 6876
rect 30656 6792 30708 6798
rect 30656 6734 30708 6740
rect 30472 6248 30524 6254
rect 30472 6190 30524 6196
rect 30378 5264 30434 5273
rect 30378 5199 30434 5208
rect 30392 2922 30420 5199
rect 30484 3641 30512 6190
rect 30564 5636 30616 5642
rect 30564 5578 30616 5584
rect 30470 3632 30526 3641
rect 30470 3567 30526 3576
rect 30380 2916 30432 2922
rect 30380 2858 30432 2864
rect 30576 2854 30604 5578
rect 30668 5166 30696 6734
rect 30656 5160 30708 5166
rect 30656 5102 30708 5108
rect 30656 3528 30708 3534
rect 30656 3470 30708 3476
rect 30668 2990 30696 3470
rect 30656 2984 30708 2990
rect 30656 2926 30708 2932
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31128 2009 31156 2246
rect 31114 2000 31170 2009
rect 31114 1935 31170 1944
rect 31220 56 31248 7346
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 32324 7002 32352 7822
rect 32416 7410 32444 7890
rect 32496 7744 32548 7750
rect 32496 7686 32548 7692
rect 32508 7449 32536 7686
rect 32600 7546 32628 9279
rect 33414 9072 33470 9081
rect 33414 9007 33470 9016
rect 32680 8900 32732 8906
rect 32680 8842 32732 8848
rect 32692 8498 32720 8842
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32864 8356 32916 8362
rect 32864 8298 32916 8304
rect 32876 7993 32904 8298
rect 33428 8090 33456 9007
rect 33416 8084 33468 8090
rect 33416 8026 33468 8032
rect 32862 7984 32918 7993
rect 32862 7919 32918 7928
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 32588 7540 32640 7546
rect 32588 7482 32640 7488
rect 32494 7440 32550 7449
rect 32404 7404 32456 7410
rect 32494 7375 32550 7384
rect 32404 7346 32456 7352
rect 32692 7274 32720 7822
rect 33600 7744 33652 7750
rect 33598 7712 33600 7721
rect 33652 7712 33654 7721
rect 33010 7644 33318 7653
rect 33598 7647 33654 7656
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 32772 7472 32824 7478
rect 32772 7414 32824 7420
rect 32680 7268 32732 7274
rect 32680 7210 32732 7216
rect 32312 6996 32364 7002
rect 32312 6938 32364 6944
rect 32404 6792 32456 6798
rect 32404 6734 32456 6740
rect 32312 6316 32364 6322
rect 32312 6258 32364 6264
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32324 5914 32352 6258
rect 32312 5908 32364 5914
rect 32312 5850 32364 5856
rect 32416 5778 32444 6734
rect 32496 6112 32548 6118
rect 32494 6080 32496 6089
rect 32548 6080 32550 6089
rect 32494 6015 32550 6024
rect 32404 5772 32456 5778
rect 32404 5714 32456 5720
rect 32312 5228 32364 5234
rect 32312 5170 32364 5176
rect 31760 5024 31812 5030
rect 31760 4966 31812 4972
rect 31668 4752 31720 4758
rect 31668 4694 31720 4700
rect 31680 4146 31708 4694
rect 31668 4140 31720 4146
rect 31668 4082 31720 4088
rect 31300 2644 31352 2650
rect 31300 2586 31352 2592
rect 31312 2446 31340 2586
rect 31772 2446 31800 4966
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 32324 4593 32352 5170
rect 32496 5024 32548 5030
rect 32494 4992 32496 5001
rect 32548 4992 32550 5001
rect 32494 4927 32550 4936
rect 32310 4584 32366 4593
rect 32310 4519 32366 4528
rect 32404 4480 32456 4486
rect 32404 4422 32456 4428
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 32416 3534 32444 4422
rect 32496 3936 32548 3942
rect 32494 3904 32496 3913
rect 32548 3904 32550 3913
rect 32494 3839 32550 3848
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 31852 3120 31904 3126
rect 32036 3120 32088 3126
rect 31904 3068 32036 3074
rect 31852 3062 32088 3068
rect 31864 3046 32076 3062
rect 31852 2848 31904 2854
rect 32496 2848 32548 2854
rect 31852 2790 31904 2796
rect 32494 2816 32496 2825
rect 32548 2816 32550 2825
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 31760 2440 31812 2446
rect 31760 2382 31812 2388
rect 31864 2394 31892 2790
rect 31950 2748 32258 2757
rect 32494 2751 32550 2760
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 31864 2366 31984 2394
rect 31484 2304 31536 2310
rect 31484 2246 31536 2252
rect 31852 2304 31904 2310
rect 31852 2246 31904 2252
rect 31496 1465 31524 2246
rect 31482 1456 31538 1465
rect 31482 1391 31538 1400
rect 31864 1193 31892 2246
rect 31956 1737 31984 2366
rect 31942 1728 31998 1737
rect 31942 1663 31998 1672
rect 31850 1184 31906 1193
rect 31850 1119 31906 1128
rect 32784 56 32812 7414
rect 32864 7200 32916 7206
rect 32862 7168 32864 7177
rect 32916 7168 32918 7177
rect 32862 7103 32918 7112
rect 32862 6896 32918 6905
rect 32862 6831 32918 6840
rect 32876 6662 32904 6831
rect 33416 6724 33468 6730
rect 33416 6666 33468 6672
rect 32864 6656 32916 6662
rect 33428 6633 33456 6666
rect 32864 6598 32916 6604
rect 33414 6624 33470 6633
rect 33010 6556 33318 6565
rect 33414 6559 33470 6568
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 32864 6452 32916 6458
rect 32864 6394 32916 6400
rect 32876 6361 32904 6394
rect 32862 6352 32918 6361
rect 32862 6287 32918 6296
rect 32864 5840 32916 5846
rect 32862 5808 32864 5817
rect 32916 5808 32918 5817
rect 32862 5743 32918 5752
rect 33416 5568 33468 5574
rect 33414 5536 33416 5545
rect 33468 5536 33470 5545
rect 33010 5468 33318 5477
rect 33414 5471 33470 5480
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 32876 5273 32904 5306
rect 32862 5264 32918 5273
rect 32862 5199 32918 5208
rect 32864 4752 32916 4758
rect 32862 4720 32864 4729
rect 32916 4720 32918 4729
rect 32862 4655 32918 4664
rect 33416 4480 33468 4486
rect 33414 4448 33416 4457
rect 33468 4448 33470 4457
rect 33010 4380 33318 4389
rect 33414 4383 33470 4392
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 32862 4176 32918 4185
rect 32862 4111 32918 4120
rect 32876 4010 32904 4111
rect 32864 4004 32916 4010
rect 32864 3946 32916 3952
rect 32864 3664 32916 3670
rect 32862 3632 32864 3641
rect 32916 3632 32918 3641
rect 32862 3567 32918 3576
rect 33416 3392 33468 3398
rect 33414 3360 33416 3369
rect 33468 3360 33470 3369
rect 33010 3292 33318 3301
rect 33414 3295 33470 3304
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32864 3188 32916 3194
rect 32864 3130 32916 3136
rect 32876 3097 32904 3130
rect 32862 3088 32918 3097
rect 32862 3023 32918 3032
rect 32864 2576 32916 2582
rect 32862 2544 32864 2553
rect 32916 2544 32918 2553
rect 32862 2479 32918 2488
rect 33416 2304 33468 2310
rect 33414 2272 33416 2281
rect 33468 2272 33470 2281
rect 33010 2204 33318 2213
rect 33414 2207 33470 2216
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 24860 2 24912 8
rect 24950 0 25006 56
rect 26514 0 26570 56
rect 28078 0 28134 56
rect 29642 0 29698 56
rect 31206 0 31262 56
rect 32770 0 32826 56
<< via2 >>
rect 5078 9560 5134 9616
rect 1030 8200 1086 8256
rect 2870 9152 2926 9208
rect 2870 8744 2926 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1306 7656 1362 7712
rect 294 7384 350 7440
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 3514 6840 3570 6896
rect 2778 6568 2834 6624
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 2870 5480 2926 5536
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2962 5208 3018 5264
rect 2870 4664 2926 4720
rect 3422 4392 3478 4448
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 5354 9288 5410 9344
rect 5078 7248 5134 7304
rect 4894 6704 4950 6760
rect 5354 7384 5410 7440
rect 4710 6296 4766 6352
rect 4066 6160 4122 6216
rect 6826 6860 6882 6896
rect 6826 6840 6828 6860
rect 6828 6840 6880 6860
rect 6880 6840 6882 6860
rect 7378 9424 7434 9480
rect 7378 8472 7434 8528
rect 7470 8200 7526 8256
rect 7562 7928 7618 7984
rect 8298 11056 8354 11112
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 7746 6316 7802 6352
rect 7746 6296 7748 6316
rect 7748 6296 7800 6316
rect 7800 6296 7802 6316
rect 8482 9696 8538 9752
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 7378 5752 7434 5808
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 8482 5072 8538 5128
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 8482 4664 8538 4720
rect 8666 4664 8722 4720
rect 7286 3440 7342 3496
rect 8666 4392 8722 4448
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 9954 9832 10010 9888
rect 10506 8472 10562 8528
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 8390 3732 8446 3768
rect 10598 7928 10654 7984
rect 10782 7520 10838 7576
rect 8390 3712 8392 3732
rect 8392 3712 8444 3732
rect 8444 3712 8446 3732
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 9402 2896 9458 2952
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 11426 9968 11482 10024
rect 12162 10104 12218 10160
rect 12162 8608 12218 8664
rect 12990 8744 13046 8800
rect 12714 7540 12770 7576
rect 12714 7520 12716 7540
rect 12716 7520 12768 7540
rect 12768 7520 12770 7540
rect 12806 3712 12862 3768
rect 11978 3440 12034 3496
rect 10966 1128 11022 1184
rect 14002 10240 14058 10296
rect 14002 8608 14058 8664
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 14738 9016 14794 9072
rect 14370 7928 14426 7984
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 15382 10104 15438 10160
rect 15566 9968 15622 10024
rect 16302 9832 16358 9888
rect 15934 9696 15990 9752
rect 15566 9560 15622 9616
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 14738 7928 14794 7984
rect 13174 4664 13230 4720
rect 12990 1944 13046 2000
rect 14002 6160 14058 6216
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13818 4800 13874 4856
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 14002 3440 14058 3496
rect 14186 3476 14188 3496
rect 14188 3476 14240 3496
rect 14240 3476 14242 3496
rect 14186 3440 14242 3476
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 16394 9152 16450 9208
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 16394 6160 16450 6216
rect 14554 3304 14610 3360
rect 14370 2760 14426 2816
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 14830 5616 14886 5672
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 15014 4664 15070 4720
rect 15474 4528 15530 4584
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 14922 3984 14978 4040
rect 15106 3984 15162 4040
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 13634 1672 13690 1728
rect 15842 3032 15898 3088
rect 16578 7792 16634 7848
rect 16762 6840 16818 6896
rect 17130 9152 17186 9208
rect 16946 6704 17002 6760
rect 16670 5652 16672 5672
rect 16672 5652 16724 5672
rect 16724 5652 16726 5672
rect 16670 5616 16726 5652
rect 16486 5072 16542 5128
rect 16486 3440 16542 3496
rect 16394 3032 16450 3088
rect 16670 2896 16726 2952
rect 18326 11056 18382 11112
rect 18510 10240 18566 10296
rect 17774 9424 17830 9480
rect 17958 9288 18014 9344
rect 18142 7268 18198 7304
rect 18142 7248 18144 7268
rect 18144 7248 18196 7268
rect 18196 7248 18198 7268
rect 17406 5752 17462 5808
rect 17590 3576 17646 3632
rect 17774 3612 17776 3632
rect 17776 3612 17828 3632
rect 17828 3612 17830 3632
rect 17774 3576 17830 3612
rect 18142 4120 18198 4176
rect 18602 7928 18658 7984
rect 19338 7520 19394 7576
rect 18878 6296 18934 6352
rect 16946 2352 17002 2408
rect 17130 1944 17186 2000
rect 15658 1400 15714 1456
rect 19614 9560 19670 9616
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19614 5208 19670 5264
rect 19798 5072 19854 5128
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 20718 8336 20774 8392
rect 20810 7520 20866 7576
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21178 7404 21234 7440
rect 21178 7384 21180 7404
rect 21180 7384 21232 7404
rect 21232 7384 21234 7404
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21454 3440 21510 3496
rect 20718 3304 20774 3360
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 21638 3032 21694 3088
rect 21822 8880 21878 8936
rect 22006 8880 22062 8936
rect 21914 7248 21970 7304
rect 22282 9696 22338 9752
rect 22558 8744 22614 8800
rect 22374 6840 22430 6896
rect 21822 5616 21878 5672
rect 21730 2896 21786 2952
rect 24766 9696 24822 9752
rect 24582 8880 24638 8936
rect 24582 8744 24638 8800
rect 23386 5072 23442 5128
rect 25134 8492 25190 8528
rect 25134 8472 25136 8492
rect 25136 8472 25188 8492
rect 25188 8472 25190 8492
rect 26422 9152 26478 9208
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 26514 6976 26570 7032
rect 26330 6840 26386 6896
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25778 3984 25834 4040
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 26974 7248 27030 7304
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 28078 5072 28134 5128
rect 31758 9560 31814 9616
rect 31298 9288 31354 9344
rect 31482 8880 31538 8936
rect 32586 9288 32642 9344
rect 31850 8472 31906 8528
rect 32494 8200 32550 8256
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 29090 6976 29146 7032
rect 28446 5616 28502 5672
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 28078 2624 28134 2680
rect 27618 1944 27674 2000
rect 29366 2624 29422 2680
rect 30378 5208 30434 5264
rect 30470 3576 30526 3632
rect 31114 1944 31170 2000
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 33414 9016 33470 9072
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 32862 7928 32918 7984
rect 32494 7384 32550 7440
rect 33598 7692 33600 7712
rect 33600 7692 33652 7712
rect 33652 7692 33654 7712
rect 33598 7656 33654 7692
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 32494 6060 32496 6080
rect 32496 6060 32548 6080
rect 32548 6060 32550 6080
rect 32494 6024 32550 6060
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 32494 4972 32496 4992
rect 32496 4972 32548 4992
rect 32548 4972 32550 4992
rect 32494 4936 32550 4972
rect 32310 4528 32366 4584
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 32494 3884 32496 3904
rect 32496 3884 32548 3904
rect 32548 3884 32550 3904
rect 32494 3848 32550 3884
rect 32494 2796 32496 2816
rect 32496 2796 32548 2816
rect 32548 2796 32550 2816
rect 32494 2760 32550 2796
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 31482 1400 31538 1456
rect 31942 1672 31998 1728
rect 31850 1128 31906 1184
rect 32862 7148 32864 7168
rect 32864 7148 32916 7168
rect 32916 7148 32918 7168
rect 32862 7112 32918 7148
rect 32862 6840 32918 6896
rect 33414 6568 33470 6624
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 32862 6296 32918 6352
rect 32862 5788 32864 5808
rect 32864 5788 32916 5808
rect 32916 5788 32918 5808
rect 32862 5752 32918 5788
rect 33414 5516 33416 5536
rect 33416 5516 33468 5536
rect 33468 5516 33470 5536
rect 33414 5480 33470 5516
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 32862 5208 32918 5264
rect 32862 4700 32864 4720
rect 32864 4700 32916 4720
rect 32916 4700 32918 4720
rect 32862 4664 32918 4700
rect 33414 4428 33416 4448
rect 33416 4428 33468 4448
rect 33468 4428 33470 4448
rect 33414 4392 33470 4428
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 32862 4120 32918 4176
rect 32862 3612 32864 3632
rect 32864 3612 32916 3632
rect 32916 3612 32918 3632
rect 32862 3576 32918 3612
rect 33414 3340 33416 3360
rect 33416 3340 33468 3360
rect 33468 3340 33470 3360
rect 33414 3304 33470 3340
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 32862 3032 32918 3088
rect 32862 2524 32864 2544
rect 32864 2524 32916 2544
rect 32916 2524 32918 2544
rect 32862 2488 32918 2524
rect 33414 2252 33416 2272
rect 33416 2252 33468 2272
rect 33468 2252 33470 2272
rect 33414 2216 33470 2252
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
<< metal3 >>
rect 8293 11114 8359 11117
rect 18321 11114 18387 11117
rect 8293 11112 18387 11114
rect 8293 11056 8298 11112
rect 8354 11056 18326 11112
rect 18382 11056 18387 11112
rect 8293 11054 18387 11056
rect 8293 11051 8359 11054
rect 18321 11051 18387 11054
rect 13997 10298 14063 10301
rect 18505 10298 18571 10301
rect 13997 10296 18571 10298
rect 13997 10240 14002 10296
rect 14058 10240 18510 10296
rect 18566 10240 18571 10296
rect 13997 10238 18571 10240
rect 13997 10235 14063 10238
rect 18505 10235 18571 10238
rect 12157 10162 12223 10165
rect 15377 10162 15443 10165
rect 12157 10160 15443 10162
rect 12157 10104 12162 10160
rect 12218 10104 15382 10160
rect 15438 10104 15443 10160
rect 12157 10102 15443 10104
rect 12157 10099 12223 10102
rect 15377 10099 15443 10102
rect 11421 10026 11487 10029
rect 15561 10026 15627 10029
rect 11421 10024 15627 10026
rect 11421 9968 11426 10024
rect 11482 9968 15566 10024
rect 15622 9968 15627 10024
rect 11421 9966 15627 9968
rect 11421 9963 11487 9966
rect 15561 9963 15627 9966
rect 9949 9890 10015 9893
rect 16297 9890 16363 9893
rect 9949 9888 16363 9890
rect 9949 9832 9954 9888
rect 10010 9832 16302 9888
rect 16358 9832 16363 9888
rect 9949 9830 16363 9832
rect 9949 9827 10015 9830
rect 16297 9827 16363 9830
rect 8477 9754 8543 9757
rect 15929 9754 15995 9757
rect 8477 9752 15995 9754
rect 8477 9696 8482 9752
rect 8538 9696 15934 9752
rect 15990 9696 15995 9752
rect 8477 9694 15995 9696
rect 8477 9691 8543 9694
rect 15929 9691 15995 9694
rect 22277 9754 22343 9757
rect 24761 9754 24827 9757
rect 22277 9752 24827 9754
rect 22277 9696 22282 9752
rect 22338 9696 24766 9752
rect 24822 9696 24827 9752
rect 22277 9694 24827 9696
rect 22277 9691 22343 9694
rect 24761 9691 24827 9694
rect 0 9618 120 9648
rect 5073 9618 5139 9621
rect 0 9616 5139 9618
rect 0 9560 5078 9616
rect 5134 9560 5139 9616
rect 0 9558 5139 9560
rect 0 9528 120 9558
rect 5073 9555 5139 9558
rect 15561 9618 15627 9621
rect 19609 9618 19675 9621
rect 15561 9616 19675 9618
rect 15561 9560 15566 9616
rect 15622 9560 19614 9616
rect 19670 9560 19675 9616
rect 15561 9558 19675 9560
rect 15561 9555 15627 9558
rect 19609 9555 19675 9558
rect 31753 9618 31819 9621
rect 34288 9618 34408 9648
rect 31753 9616 34408 9618
rect 31753 9560 31758 9616
rect 31814 9560 34408 9616
rect 31753 9558 34408 9560
rect 31753 9555 31819 9558
rect 34288 9528 34408 9558
rect 7373 9482 7439 9485
rect 17769 9482 17835 9485
rect 7373 9480 17835 9482
rect 7373 9424 7378 9480
rect 7434 9424 17774 9480
rect 17830 9424 17835 9480
rect 7373 9422 17835 9424
rect 7373 9419 7439 9422
rect 17769 9419 17835 9422
rect 0 9346 120 9376
rect 5349 9346 5415 9349
rect 0 9344 5415 9346
rect 0 9288 5354 9344
rect 5410 9288 5415 9344
rect 0 9286 5415 9288
rect 0 9256 120 9286
rect 5349 9283 5415 9286
rect 17953 9346 18019 9349
rect 31293 9346 31359 9349
rect 17953 9344 31359 9346
rect 17953 9288 17958 9344
rect 18014 9288 31298 9344
rect 31354 9288 31359 9344
rect 17953 9286 31359 9288
rect 17953 9283 18019 9286
rect 31293 9283 31359 9286
rect 32581 9346 32647 9349
rect 34288 9346 34408 9376
rect 32581 9344 34408 9346
rect 32581 9288 32586 9344
rect 32642 9288 34408 9344
rect 32581 9286 34408 9288
rect 32581 9283 32647 9286
rect 34288 9256 34408 9286
rect 2865 9210 2931 9213
rect 16389 9210 16455 9213
rect 2865 9208 16455 9210
rect 2865 9152 2870 9208
rect 2926 9152 16394 9208
rect 16450 9152 16455 9208
rect 2865 9150 16455 9152
rect 2865 9147 2931 9150
rect 16389 9147 16455 9150
rect 17125 9210 17191 9213
rect 26417 9210 26483 9213
rect 17125 9208 26483 9210
rect 17125 9152 17130 9208
rect 17186 9152 26422 9208
rect 26478 9152 26483 9208
rect 17125 9150 26483 9152
rect 17125 9147 17191 9150
rect 26417 9147 26483 9150
rect 0 9074 120 9104
rect 14733 9074 14799 9077
rect 0 9072 14799 9074
rect 0 9016 14738 9072
rect 14794 9016 14799 9072
rect 0 9014 14799 9016
rect 0 8984 120 9014
rect 14733 9011 14799 9014
rect 33409 9074 33475 9077
rect 34288 9074 34408 9104
rect 33409 9072 34408 9074
rect 33409 9016 33414 9072
rect 33470 9016 34408 9072
rect 33409 9014 34408 9016
rect 33409 9011 33475 9014
rect 34288 8984 34408 9014
rect 21817 8938 21883 8941
rect 14782 8936 21883 8938
rect 14782 8880 21822 8936
rect 21878 8880 21883 8936
rect 14782 8878 21883 8880
rect 0 8802 120 8832
rect 2865 8802 2931 8805
rect 0 8800 2931 8802
rect 0 8744 2870 8800
rect 2926 8744 2931 8800
rect 0 8742 2931 8744
rect 0 8712 120 8742
rect 2865 8739 2931 8742
rect 12985 8802 13051 8805
rect 14782 8802 14842 8878
rect 21817 8875 21883 8878
rect 22001 8938 22067 8941
rect 24577 8938 24643 8941
rect 22001 8936 24643 8938
rect 22001 8880 22006 8936
rect 22062 8880 24582 8936
rect 24638 8880 24643 8936
rect 22001 8878 24643 8880
rect 22001 8875 22067 8878
rect 24577 8875 24643 8878
rect 31477 8938 31543 8941
rect 31477 8936 33610 8938
rect 31477 8880 31482 8936
rect 31538 8880 33610 8936
rect 31477 8878 33610 8880
rect 31477 8875 31543 8878
rect 12985 8800 14842 8802
rect 12985 8744 12990 8800
rect 13046 8744 14842 8800
rect 12985 8742 14842 8744
rect 22553 8802 22619 8805
rect 24577 8802 24643 8805
rect 22553 8800 24643 8802
rect 22553 8744 22558 8800
rect 22614 8744 24582 8800
rect 24638 8744 24643 8800
rect 22553 8742 24643 8744
rect 33550 8802 33610 8878
rect 34288 8802 34408 8832
rect 33550 8742 34408 8802
rect 12985 8739 13051 8742
rect 22553 8739 22619 8742
rect 24577 8739 24643 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 34288 8712 34408 8742
rect 33006 8671 33322 8672
rect 12157 8666 12223 8669
rect 13997 8666 14063 8669
rect 12157 8664 14063 8666
rect 12157 8608 12162 8664
rect 12218 8608 14002 8664
rect 14058 8608 14063 8664
rect 12157 8606 14063 8608
rect 12157 8603 12223 8606
rect 13997 8603 14063 8606
rect 0 8530 120 8560
rect 7373 8530 7439 8533
rect 0 8528 7439 8530
rect 0 8472 7378 8528
rect 7434 8472 7439 8528
rect 0 8470 7439 8472
rect 0 8440 120 8470
rect 7373 8467 7439 8470
rect 10501 8530 10567 8533
rect 25129 8530 25195 8533
rect 10501 8528 25195 8530
rect 10501 8472 10506 8528
rect 10562 8472 25134 8528
rect 25190 8472 25195 8528
rect 10501 8470 25195 8472
rect 10501 8467 10567 8470
rect 25129 8467 25195 8470
rect 31845 8530 31911 8533
rect 34288 8530 34408 8560
rect 31845 8528 34408 8530
rect 31845 8472 31850 8528
rect 31906 8472 34408 8528
rect 31845 8470 34408 8472
rect 31845 8467 31911 8470
rect 34288 8440 34408 8470
rect 20713 8394 20779 8397
rect 1350 8392 20779 8394
rect 1350 8336 20718 8392
rect 20774 8336 20779 8392
rect 1350 8334 20779 8336
rect 0 8258 120 8288
rect 1025 8258 1091 8261
rect 0 8256 1091 8258
rect 0 8200 1030 8256
rect 1086 8200 1091 8256
rect 0 8198 1091 8200
rect 0 8168 120 8198
rect 1025 8195 1091 8198
rect 0 7986 120 8016
rect 1350 7986 1410 8334
rect 20713 8331 20779 8334
rect 7465 8258 7531 8261
rect 7422 8256 7531 8258
rect 7422 8200 7470 8256
rect 7526 8200 7531 8256
rect 7422 8195 7531 8200
rect 32489 8258 32555 8261
rect 34288 8258 34408 8288
rect 32489 8256 34408 8258
rect 32489 8200 32494 8256
rect 32550 8200 34408 8256
rect 32489 8198 34408 8200
rect 32489 8195 32555 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 0 7926 1410 7986
rect 7422 7986 7482 8195
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 34288 8168 34408 8198
rect 31946 8127 32262 8128
rect 7557 7986 7623 7989
rect 7422 7984 7623 7986
rect 7422 7928 7562 7984
rect 7618 7928 7623 7984
rect 7422 7926 7623 7928
rect 0 7896 120 7926
rect 7557 7923 7623 7926
rect 10593 7986 10659 7989
rect 14365 7986 14431 7989
rect 10593 7984 14431 7986
rect 10593 7928 10598 7984
rect 10654 7928 14370 7984
rect 14426 7928 14431 7984
rect 10593 7926 14431 7928
rect 10593 7923 10659 7926
rect 14365 7923 14431 7926
rect 14733 7986 14799 7989
rect 18597 7986 18663 7989
rect 14733 7984 18663 7986
rect 14733 7928 14738 7984
rect 14794 7928 18602 7984
rect 18658 7928 18663 7984
rect 14733 7926 18663 7928
rect 14733 7923 14799 7926
rect 18597 7923 18663 7926
rect 32857 7986 32923 7989
rect 34288 7986 34408 8016
rect 32857 7984 34408 7986
rect 32857 7928 32862 7984
rect 32918 7928 34408 7984
rect 32857 7926 34408 7928
rect 32857 7923 32923 7926
rect 34288 7896 34408 7926
rect 16573 7850 16639 7853
rect 1718 7848 16639 7850
rect 1718 7792 16578 7848
rect 16634 7792 16639 7848
rect 1718 7790 16639 7792
rect 0 7714 120 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 120 7654
rect 1301 7651 1367 7654
rect 0 7442 120 7472
rect 289 7442 355 7445
rect 0 7440 355 7442
rect 0 7384 294 7440
rect 350 7384 355 7440
rect 0 7382 355 7384
rect 0 7352 120 7382
rect 289 7379 355 7382
rect 0 7170 120 7200
rect 1718 7170 1778 7790
rect 16573 7787 16639 7790
rect 33593 7714 33659 7717
rect 34288 7714 34408 7744
rect 33593 7712 34408 7714
rect 33593 7656 33598 7712
rect 33654 7656 34408 7712
rect 33593 7654 34408 7656
rect 33593 7651 33659 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 34288 7624 34408 7654
rect 33006 7583 33322 7584
rect 10777 7578 10843 7581
rect 12709 7578 12775 7581
rect 10777 7576 12775 7578
rect 10777 7520 10782 7576
rect 10838 7520 12714 7576
rect 12770 7520 12775 7576
rect 10777 7518 12775 7520
rect 10777 7515 10843 7518
rect 12709 7515 12775 7518
rect 19333 7578 19399 7581
rect 20805 7578 20871 7581
rect 19333 7576 20871 7578
rect 19333 7520 19338 7576
rect 19394 7520 20810 7576
rect 20866 7520 20871 7576
rect 19333 7518 20871 7520
rect 19333 7515 19399 7518
rect 20805 7515 20871 7518
rect 5349 7442 5415 7445
rect 21173 7442 21239 7445
rect 5349 7440 21239 7442
rect 5349 7384 5354 7440
rect 5410 7384 21178 7440
rect 21234 7384 21239 7440
rect 5349 7382 21239 7384
rect 5349 7379 5415 7382
rect 21173 7379 21239 7382
rect 32489 7442 32555 7445
rect 34288 7442 34408 7472
rect 32489 7440 34408 7442
rect 32489 7384 32494 7440
rect 32550 7384 34408 7440
rect 32489 7382 34408 7384
rect 32489 7379 32555 7382
rect 34288 7352 34408 7382
rect 5073 7306 5139 7309
rect 18137 7306 18203 7309
rect 5073 7304 18203 7306
rect 5073 7248 5078 7304
rect 5134 7248 18142 7304
rect 18198 7248 18203 7304
rect 5073 7246 18203 7248
rect 5073 7243 5139 7246
rect 18137 7243 18203 7246
rect 21909 7306 21975 7309
rect 26969 7306 27035 7309
rect 21909 7304 27035 7306
rect 21909 7248 21914 7304
rect 21970 7248 26974 7304
rect 27030 7248 27035 7304
rect 21909 7246 27035 7248
rect 21909 7243 21975 7246
rect 26969 7243 27035 7246
rect 0 7110 1778 7170
rect 32857 7170 32923 7173
rect 34288 7170 34408 7200
rect 32857 7168 34408 7170
rect 32857 7112 32862 7168
rect 32918 7112 34408 7168
rect 32857 7110 34408 7112
rect 0 7080 120 7110
rect 32857 7107 32923 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 34288 7080 34408 7110
rect 31946 7039 32262 7040
rect 26509 7034 26575 7037
rect 29085 7034 29151 7037
rect 26509 7032 29151 7034
rect 26509 6976 26514 7032
rect 26570 6976 29090 7032
rect 29146 6976 29151 7032
rect 26509 6974 29151 6976
rect 26509 6971 26575 6974
rect 29085 6971 29151 6974
rect 0 6898 120 6928
rect 3509 6898 3575 6901
rect 0 6896 3575 6898
rect 0 6840 3514 6896
rect 3570 6840 3575 6896
rect 0 6838 3575 6840
rect 0 6808 120 6838
rect 3509 6835 3575 6838
rect 6821 6898 6887 6901
rect 16757 6898 16823 6901
rect 6821 6896 16823 6898
rect 6821 6840 6826 6896
rect 6882 6840 16762 6896
rect 16818 6840 16823 6896
rect 6821 6838 16823 6840
rect 6821 6835 6887 6838
rect 16757 6835 16823 6838
rect 22369 6898 22435 6901
rect 26325 6898 26391 6901
rect 22369 6896 26391 6898
rect 22369 6840 22374 6896
rect 22430 6840 26330 6896
rect 26386 6840 26391 6896
rect 22369 6838 26391 6840
rect 22369 6835 22435 6838
rect 26325 6835 26391 6838
rect 32857 6898 32923 6901
rect 34288 6898 34408 6928
rect 32857 6896 34408 6898
rect 32857 6840 32862 6896
rect 32918 6840 34408 6896
rect 32857 6838 34408 6840
rect 32857 6835 32923 6838
rect 34288 6808 34408 6838
rect 4889 6762 4955 6765
rect 16941 6762 17007 6765
rect 4889 6760 17007 6762
rect 4889 6704 4894 6760
rect 4950 6704 16946 6760
rect 17002 6704 17007 6760
rect 4889 6702 17007 6704
rect 4889 6699 4955 6702
rect 16941 6699 17007 6702
rect 0 6626 120 6656
rect 2773 6626 2839 6629
rect 0 6624 2839 6626
rect 0 6568 2778 6624
rect 2834 6568 2839 6624
rect 0 6566 2839 6568
rect 0 6536 120 6566
rect 2773 6563 2839 6566
rect 33409 6626 33475 6629
rect 34288 6626 34408 6656
rect 33409 6624 34408 6626
rect 33409 6568 33414 6624
rect 33470 6568 34408 6624
rect 33409 6566 34408 6568
rect 33409 6563 33475 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 34288 6536 34408 6566
rect 33006 6495 33322 6496
rect 0 6354 120 6384
rect 4705 6354 4771 6357
rect 0 6352 4771 6354
rect 0 6296 4710 6352
rect 4766 6296 4771 6352
rect 0 6294 4771 6296
rect 0 6264 120 6294
rect 4705 6291 4771 6294
rect 7741 6354 7807 6357
rect 18873 6354 18939 6357
rect 7741 6352 18939 6354
rect 7741 6296 7746 6352
rect 7802 6296 18878 6352
rect 18934 6296 18939 6352
rect 7741 6294 18939 6296
rect 7741 6291 7807 6294
rect 18873 6291 18939 6294
rect 32857 6354 32923 6357
rect 34288 6354 34408 6384
rect 32857 6352 34408 6354
rect 32857 6296 32862 6352
rect 32918 6296 34408 6352
rect 32857 6294 34408 6296
rect 32857 6291 32923 6294
rect 34288 6264 34408 6294
rect 4061 6218 4127 6221
rect 1718 6216 4127 6218
rect 1718 6160 4066 6216
rect 4122 6160 4127 6216
rect 1718 6158 4127 6160
rect 0 6082 120 6112
rect 1718 6082 1778 6158
rect 4061 6155 4127 6158
rect 13997 6218 14063 6221
rect 16389 6218 16455 6221
rect 13997 6216 16455 6218
rect 13997 6160 14002 6216
rect 14058 6160 16394 6216
rect 16450 6160 16455 6216
rect 13997 6158 16455 6160
rect 13997 6155 14063 6158
rect 16389 6155 16455 6158
rect 0 6022 1778 6082
rect 32489 6082 32555 6085
rect 34288 6082 34408 6112
rect 32489 6080 34408 6082
rect 32489 6024 32494 6080
rect 32550 6024 34408 6080
rect 32489 6022 34408 6024
rect 0 5992 120 6022
rect 32489 6019 32555 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 34288 5992 34408 6022
rect 31946 5951 32262 5952
rect 0 5810 120 5840
rect 7373 5810 7439 5813
rect 17401 5810 17467 5813
rect 0 5750 2790 5810
rect 0 5720 120 5750
rect 2730 5674 2790 5750
rect 7373 5808 17467 5810
rect 7373 5752 7378 5808
rect 7434 5752 17406 5808
rect 17462 5752 17467 5808
rect 7373 5750 17467 5752
rect 7373 5747 7439 5750
rect 17401 5747 17467 5750
rect 32857 5810 32923 5813
rect 34288 5810 34408 5840
rect 32857 5808 34408 5810
rect 32857 5752 32862 5808
rect 32918 5752 34408 5808
rect 32857 5750 34408 5752
rect 32857 5747 32923 5750
rect 34288 5720 34408 5750
rect 14825 5674 14891 5677
rect 16665 5676 16731 5677
rect 16614 5674 16620 5676
rect 2730 5672 14891 5674
rect 2730 5616 14830 5672
rect 14886 5616 14891 5672
rect 2730 5614 14891 5616
rect 16574 5614 16620 5674
rect 16684 5672 16731 5676
rect 16726 5616 16731 5672
rect 14825 5611 14891 5614
rect 16614 5612 16620 5614
rect 16684 5612 16731 5616
rect 16665 5611 16731 5612
rect 21817 5674 21883 5677
rect 28441 5674 28507 5677
rect 21817 5672 28507 5674
rect 21817 5616 21822 5672
rect 21878 5616 28446 5672
rect 28502 5616 28507 5672
rect 21817 5614 28507 5616
rect 21817 5611 21883 5614
rect 28441 5611 28507 5614
rect 0 5538 120 5568
rect 2865 5538 2931 5541
rect 0 5536 2931 5538
rect 0 5480 2870 5536
rect 2926 5480 2931 5536
rect 0 5478 2931 5480
rect 0 5448 120 5478
rect 2865 5475 2931 5478
rect 33409 5538 33475 5541
rect 34288 5538 34408 5568
rect 33409 5536 34408 5538
rect 33409 5480 33414 5536
rect 33470 5480 34408 5536
rect 33409 5478 34408 5480
rect 33409 5475 33475 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 34288 5448 34408 5478
rect 33006 5407 33322 5408
rect 0 5266 120 5296
rect 2814 5266 2820 5268
rect 0 5206 2820 5266
rect 0 5176 120 5206
rect 2814 5204 2820 5206
rect 2884 5204 2890 5268
rect 2957 5266 3023 5269
rect 19609 5266 19675 5269
rect 30373 5266 30439 5269
rect 2957 5264 19675 5266
rect 2957 5208 2962 5264
rect 3018 5208 19614 5264
rect 19670 5208 19675 5264
rect 2957 5206 19675 5208
rect 2957 5203 3023 5206
rect 19609 5203 19675 5206
rect 22050 5264 30439 5266
rect 22050 5208 30378 5264
rect 30434 5208 30439 5264
rect 22050 5206 30439 5208
rect 8477 5130 8543 5133
rect 16481 5130 16547 5133
rect 1718 5070 8402 5130
rect 0 4994 120 5024
rect 1718 4994 1778 5070
rect 0 4934 1778 4994
rect 0 4904 120 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 2814 4796 2820 4860
rect 2884 4858 2890 4860
rect 8342 4858 8402 5070
rect 8477 5128 16547 5130
rect 8477 5072 8482 5128
rect 8538 5072 16486 5128
rect 16542 5072 16547 5128
rect 8477 5070 16547 5072
rect 8477 5067 8543 5070
rect 16481 5067 16547 5070
rect 19793 5130 19859 5133
rect 22050 5130 22110 5206
rect 30373 5203 30439 5206
rect 32857 5266 32923 5269
rect 34288 5266 34408 5296
rect 32857 5264 34408 5266
rect 32857 5208 32862 5264
rect 32918 5208 34408 5264
rect 32857 5206 34408 5208
rect 32857 5203 32923 5206
rect 34288 5176 34408 5206
rect 19793 5128 22110 5130
rect 19793 5072 19798 5128
rect 19854 5072 22110 5128
rect 19793 5070 22110 5072
rect 23381 5130 23447 5133
rect 28073 5130 28139 5133
rect 23381 5128 28139 5130
rect 23381 5072 23386 5128
rect 23442 5072 28078 5128
rect 28134 5072 28139 5128
rect 23381 5070 28139 5072
rect 19793 5067 19859 5070
rect 23381 5067 23447 5070
rect 28073 5067 28139 5070
rect 32489 4994 32555 4997
rect 34288 4994 34408 5024
rect 32489 4992 34408 4994
rect 32489 4936 32494 4992
rect 32550 4936 34408 4992
rect 32489 4934 34408 4936
rect 32489 4931 32555 4934
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 34288 4904 34408 4934
rect 31946 4863 32262 4864
rect 13813 4858 13879 4861
rect 2884 4798 3066 4858
rect 8342 4856 13879 4858
rect 8342 4800 13818 4856
rect 13874 4800 13879 4856
rect 8342 4798 13879 4800
rect 2884 4796 2890 4798
rect 0 4722 120 4752
rect 2865 4722 2931 4725
rect 0 4720 2931 4722
rect 0 4664 2870 4720
rect 2926 4664 2931 4720
rect 0 4662 2931 4664
rect 3006 4722 3066 4798
rect 13813 4795 13879 4798
rect 8477 4722 8543 4725
rect 3006 4720 8543 4722
rect 3006 4664 8482 4720
rect 8538 4664 8543 4720
rect 3006 4662 8543 4664
rect 0 4632 120 4662
rect 2865 4659 2931 4662
rect 8477 4659 8543 4662
rect 8661 4722 8727 4725
rect 13169 4722 13235 4725
rect 8661 4720 13235 4722
rect 8661 4664 8666 4720
rect 8722 4664 13174 4720
rect 13230 4664 13235 4720
rect 8661 4662 13235 4664
rect 8661 4659 8727 4662
rect 13169 4659 13235 4662
rect 15009 4722 15075 4725
rect 32857 4722 32923 4725
rect 34288 4722 34408 4752
rect 15009 4720 22110 4722
rect 15009 4664 15014 4720
rect 15070 4664 22110 4720
rect 15009 4662 22110 4664
rect 15009 4659 15075 4662
rect 15469 4586 15535 4589
rect 2730 4584 15535 4586
rect 2730 4528 15474 4584
rect 15530 4528 15535 4584
rect 2730 4526 15535 4528
rect 22050 4586 22110 4662
rect 32857 4720 34408 4722
rect 32857 4664 32862 4720
rect 32918 4664 34408 4720
rect 32857 4662 34408 4664
rect 32857 4659 32923 4662
rect 34288 4632 34408 4662
rect 32305 4586 32371 4589
rect 22050 4584 32371 4586
rect 22050 4528 32310 4584
rect 32366 4528 32371 4584
rect 22050 4526 32371 4528
rect 0 4450 120 4480
rect 2730 4450 2790 4526
rect 15469 4523 15535 4526
rect 32305 4523 32371 4526
rect 0 4390 2790 4450
rect 3417 4450 3483 4453
rect 8661 4450 8727 4453
rect 3417 4448 8727 4450
rect 3417 4392 3422 4448
rect 3478 4392 8666 4448
rect 8722 4392 8727 4448
rect 3417 4390 8727 4392
rect 0 4360 120 4390
rect 3417 4387 3483 4390
rect 8661 4387 8727 4390
rect 33409 4450 33475 4453
rect 34288 4450 34408 4480
rect 33409 4448 34408 4450
rect 33409 4392 33414 4448
rect 33470 4392 34408 4448
rect 33409 4390 34408 4392
rect 33409 4387 33475 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 34288 4360 34408 4390
rect 33006 4319 33322 4320
rect 0 4178 120 4208
rect 18137 4178 18203 4181
rect 0 4176 18203 4178
rect 0 4120 18142 4176
rect 18198 4120 18203 4176
rect 0 4118 18203 4120
rect 0 4088 120 4118
rect 18137 4115 18203 4118
rect 32857 4178 32923 4181
rect 34288 4178 34408 4208
rect 32857 4176 34408 4178
rect 32857 4120 32862 4176
rect 32918 4120 34408 4176
rect 32857 4118 34408 4120
rect 32857 4115 32923 4118
rect 34288 4088 34408 4118
rect 14917 4042 14983 4045
rect 1718 4040 14983 4042
rect 1718 3984 14922 4040
rect 14978 3984 14983 4040
rect 1718 3982 14983 3984
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 14917 3979 14983 3982
rect 15101 4042 15167 4045
rect 25773 4042 25839 4045
rect 15101 4040 25839 4042
rect 15101 3984 15106 4040
rect 15162 3984 25778 4040
rect 25834 3984 25839 4040
rect 15101 3982 25839 3984
rect 15101 3979 15167 3982
rect 25773 3979 25839 3982
rect 0 3846 1778 3906
rect 32489 3906 32555 3909
rect 34288 3906 34408 3936
rect 32489 3904 34408 3906
rect 32489 3848 32494 3904
rect 32550 3848 34408 3904
rect 32489 3846 34408 3848
rect 0 3816 120 3846
rect 32489 3843 32555 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 34288 3816 34408 3846
rect 31946 3775 32262 3776
rect 8385 3770 8451 3773
rect 12801 3770 12867 3773
rect 8385 3768 12867 3770
rect 8385 3712 8390 3768
rect 8446 3712 12806 3768
rect 12862 3712 12867 3768
rect 8385 3710 12867 3712
rect 8385 3707 8451 3710
rect 12801 3707 12867 3710
rect 0 3634 120 3664
rect 17585 3634 17651 3637
rect 0 3632 17651 3634
rect 0 3576 17590 3632
rect 17646 3576 17651 3632
rect 0 3574 17651 3576
rect 0 3544 120 3574
rect 17585 3571 17651 3574
rect 17769 3634 17835 3637
rect 30465 3634 30531 3637
rect 17769 3632 30531 3634
rect 17769 3576 17774 3632
rect 17830 3576 30470 3632
rect 30526 3576 30531 3632
rect 17769 3574 30531 3576
rect 17769 3571 17835 3574
rect 30465 3571 30531 3574
rect 32857 3634 32923 3637
rect 34288 3634 34408 3664
rect 32857 3632 34408 3634
rect 32857 3576 32862 3632
rect 32918 3576 34408 3632
rect 32857 3574 34408 3576
rect 32857 3571 32923 3574
rect 34288 3544 34408 3574
rect 7281 3498 7347 3501
rect 11973 3498 12039 3501
rect 13997 3498 14063 3501
rect 2730 3496 7347 3498
rect 2730 3440 7286 3496
rect 7342 3440 7347 3496
rect 2730 3438 7347 3440
rect 0 3362 120 3392
rect 2730 3362 2790 3438
rect 7281 3435 7347 3438
rect 7422 3438 9506 3498
rect 0 3302 2790 3362
rect 0 3272 120 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 0 3090 120 3120
rect 7422 3090 7482 3438
rect 9446 3362 9506 3438
rect 11973 3496 14063 3498
rect 11973 3440 11978 3496
rect 12034 3440 14002 3496
rect 14058 3440 14063 3496
rect 11973 3438 14063 3440
rect 11973 3435 12039 3438
rect 13997 3435 14063 3438
rect 14181 3498 14247 3501
rect 16481 3498 16547 3501
rect 21449 3498 21515 3501
rect 14181 3496 16314 3498
rect 14181 3440 14186 3496
rect 14242 3440 16314 3496
rect 14181 3438 16314 3440
rect 14181 3435 14247 3438
rect 14549 3362 14615 3365
rect 9446 3360 14615 3362
rect 9446 3304 14554 3360
rect 14610 3304 14615 3360
rect 9446 3302 14615 3304
rect 16254 3362 16314 3438
rect 16481 3496 21515 3498
rect 16481 3440 16486 3496
rect 16542 3440 21454 3496
rect 21510 3440 21515 3496
rect 16481 3438 21515 3440
rect 16481 3435 16547 3438
rect 21449 3435 21515 3438
rect 20713 3362 20779 3365
rect 16254 3360 20779 3362
rect 16254 3304 20718 3360
rect 20774 3304 20779 3360
rect 16254 3302 20779 3304
rect 14549 3299 14615 3302
rect 20713 3299 20779 3302
rect 33409 3362 33475 3365
rect 34288 3362 34408 3392
rect 33409 3360 34408 3362
rect 33409 3304 33414 3360
rect 33470 3304 34408 3360
rect 33409 3302 34408 3304
rect 33409 3299 33475 3302
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 34288 3272 34408 3302
rect 33006 3231 33322 3232
rect 15837 3090 15903 3093
rect 0 3030 7482 3090
rect 7606 3088 15903 3090
rect 7606 3032 15842 3088
rect 15898 3032 15903 3088
rect 7606 3030 15903 3032
rect 0 3000 120 3030
rect 7606 2954 7666 3030
rect 15837 3027 15903 3030
rect 16389 3090 16455 3093
rect 21633 3090 21699 3093
rect 16389 3088 21699 3090
rect 16389 3032 16394 3088
rect 16450 3032 21638 3088
rect 21694 3032 21699 3088
rect 16389 3030 21699 3032
rect 16389 3027 16455 3030
rect 21633 3027 21699 3030
rect 32857 3090 32923 3093
rect 34288 3090 34408 3120
rect 32857 3088 34408 3090
rect 32857 3032 32862 3088
rect 32918 3032 34408 3088
rect 32857 3030 34408 3032
rect 32857 3027 32923 3030
rect 34288 3000 34408 3030
rect 1718 2894 7666 2954
rect 9397 2954 9463 2957
rect 16665 2954 16731 2957
rect 21725 2954 21791 2957
rect 9397 2952 16731 2954
rect 9397 2896 9402 2952
rect 9458 2896 16670 2952
rect 16726 2896 16731 2952
rect 9397 2894 16731 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 9397 2891 9463 2894
rect 16665 2891 16731 2894
rect 19750 2952 21791 2954
rect 19750 2896 21730 2952
rect 21786 2896 21791 2952
rect 19750 2894 21791 2896
rect 0 2758 1778 2818
rect 14365 2818 14431 2821
rect 19750 2818 19810 2894
rect 21725 2891 21791 2894
rect 14365 2816 19810 2818
rect 14365 2760 14370 2816
rect 14426 2760 19810 2816
rect 14365 2758 19810 2760
rect 32489 2818 32555 2821
rect 34288 2818 34408 2848
rect 32489 2816 34408 2818
rect 32489 2760 32494 2816
rect 32550 2760 34408 2816
rect 32489 2758 34408 2760
rect 0 2728 120 2758
rect 14365 2755 14431 2758
rect 32489 2755 32555 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 34288 2728 34408 2758
rect 31946 2687 32262 2688
rect 28073 2682 28139 2685
rect 29361 2682 29427 2685
rect 28073 2680 29427 2682
rect 28073 2624 28078 2680
rect 28134 2624 29366 2680
rect 29422 2624 29427 2680
rect 28073 2622 29427 2624
rect 28073 2619 28139 2622
rect 29361 2619 29427 2622
rect 0 2546 120 2576
rect 16614 2546 16620 2548
rect 0 2486 16620 2546
rect 0 2456 120 2486
rect 16614 2484 16620 2486
rect 16684 2484 16690 2548
rect 32857 2546 32923 2549
rect 34288 2546 34408 2576
rect 32857 2544 34408 2546
rect 32857 2488 32862 2544
rect 32918 2488 34408 2544
rect 32857 2486 34408 2488
rect 32857 2483 32923 2486
rect 34288 2456 34408 2486
rect 16941 2410 17007 2413
rect 2822 2408 17007 2410
rect 2822 2352 16946 2408
rect 17002 2352 17007 2408
rect 2822 2350 17007 2352
rect 0 2274 120 2304
rect 2822 2274 2882 2350
rect 16941 2347 17007 2350
rect 0 2214 2882 2274
rect 33409 2274 33475 2277
rect 34288 2274 34408 2304
rect 33409 2272 34408 2274
rect 33409 2216 33414 2272
rect 33470 2216 34408 2272
rect 33409 2214 34408 2216
rect 0 2184 120 2214
rect 33409 2211 33475 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 34288 2184 34408 2214
rect 33006 2143 33322 2144
rect 0 2002 120 2032
rect 12985 2002 13051 2005
rect 0 2000 13051 2002
rect 0 1944 12990 2000
rect 13046 1944 13051 2000
rect 0 1942 13051 1944
rect 0 1912 120 1942
rect 12985 1939 13051 1942
rect 17125 2002 17191 2005
rect 27613 2002 27679 2005
rect 17125 2000 27679 2002
rect 17125 1944 17130 2000
rect 17186 1944 27618 2000
rect 27674 1944 27679 2000
rect 17125 1942 27679 1944
rect 17125 1939 17191 1942
rect 27613 1939 27679 1942
rect 31109 2002 31175 2005
rect 34288 2002 34408 2032
rect 31109 2000 34408 2002
rect 31109 1944 31114 2000
rect 31170 1944 34408 2000
rect 31109 1942 34408 1944
rect 31109 1939 31175 1942
rect 34288 1912 34408 1942
rect 0 1730 120 1760
rect 13629 1730 13695 1733
rect 0 1728 13695 1730
rect 0 1672 13634 1728
rect 13690 1672 13695 1728
rect 0 1670 13695 1672
rect 0 1640 120 1670
rect 13629 1667 13695 1670
rect 31937 1730 32003 1733
rect 34288 1730 34408 1760
rect 31937 1728 34408 1730
rect 31937 1672 31942 1728
rect 31998 1672 34408 1728
rect 31937 1670 34408 1672
rect 31937 1667 32003 1670
rect 34288 1640 34408 1670
rect 0 1458 120 1488
rect 15653 1458 15719 1461
rect 0 1456 15719 1458
rect 0 1400 15658 1456
rect 15714 1400 15719 1456
rect 0 1398 15719 1400
rect 0 1368 120 1398
rect 15653 1395 15719 1398
rect 31477 1458 31543 1461
rect 34288 1458 34408 1488
rect 31477 1456 34408 1458
rect 31477 1400 31482 1456
rect 31538 1400 34408 1456
rect 31477 1398 34408 1400
rect 31477 1395 31543 1398
rect 34288 1368 34408 1398
rect 0 1186 120 1216
rect 10961 1186 11027 1189
rect 0 1184 11027 1186
rect 0 1128 10966 1184
rect 11022 1128 11027 1184
rect 0 1126 11027 1128
rect 0 1096 120 1126
rect 10961 1123 11027 1126
rect 31845 1186 31911 1189
rect 34288 1186 34408 1216
rect 31845 1184 34408 1186
rect 31845 1128 31850 1184
rect 31906 1128 34408 1184
rect 31845 1126 34408 1128
rect 31845 1123 31911 1126
rect 34288 1096 34408 1126
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 16620 5672 16684 5676
rect 16620 5616 16670 5672
rect 16670 5616 16684 5672
rect 16620 5612 16684 5616
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 2820 5204 2884 5268
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 2820 4796 2884 4860
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 16620 2484 16684 2548
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
<< metal4 >>
rect 1944 8192 2264 11152
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 3004 8736 3324 11152
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 2819 5268 2885 5269
rect 2819 5204 2820 5268
rect 2884 5204 2885 5268
rect 2819 5203 2885 5204
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 2822 4861 2882 5203
rect 2819 4860 2885 4861
rect 2819 4796 2820 4860
rect 2884 4796 2885 4860
rect 2819 4795 2885 4796
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11152
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11152
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11152
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11152
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 19944 8192 20264 11152
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 16619 5676 16685 5677
rect 16619 5612 16620 5676
rect 16684 5612 16685 5676
rect 16619 5611 16685 5612
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 16622 2549 16682 5611
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 16619 2548 16685 2549
rect 16619 2484 16620 2548
rect 16684 2484 16685 2548
rect 16619 2483 16685 2484
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 0 20264 2688
rect 21004 8736 21324 11152
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11152
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11152
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11152
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11152
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 14352 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _002_
timestamp -3599
transform 1 0 15180 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _003_
timestamp -3599
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _004_
timestamp -3599
transform 1 0 13524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _005_
timestamp -3599
transform 1 0 17296 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform 1 0 16652 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 17572 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _009_
timestamp -3599
transform 1 0 14076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 17848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 15640 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _014_
timestamp -3599
transform 1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _015_
timestamp -3599
transform 1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _016_
timestamp -3599
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _018_
timestamp -3599
transform 1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _021_
timestamp -3599
transform 1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 20424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _023_
timestamp -3599
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 20424 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _025_
timestamp -3599
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _026_
timestamp -3599
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 19320 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _029_
timestamp -3599
transform 1 0 16744 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_
timestamp -3599
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _032_
timestamp -3599
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _033_
timestamp -3599
transform 1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _034_
timestamp -3599
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _035_
timestamp -3599
transform 1 0 14260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _036_
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp -3599
transform -1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp -3599
transform -1 0 21804 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp -3599
transform -1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform -1 0 27324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp -3599
transform 1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp -3599
transform 1 0 29624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp -3599
transform 1 0 28796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp -3599
transform 1 0 29072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform 1 0 28612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform -1 0 28612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform 1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform 1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform 1 0 29992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform 1 0 30636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp -3599
transform 1 0 29716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp -3599
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp -3599
transform -1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp -3599
transform -1 0 3128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp -3599
transform -1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp -3599
transform -1 0 5060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp -3599
transform -1 0 4784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp -3599
transform -1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp -3599
transform -1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp -3599
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp -3599
transform -1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp -3599
transform -1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp -3599
transform -1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp -3599
transform 1 0 7544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp -3599
transform 1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp -3599
transform 1 0 8096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp -3599
transform -1 0 7544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp -3599
transform -1 0 7268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp -3599
transform -1 0 7544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp -3599
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp -3599
transform -1 0 7452 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp -3599
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp -3599
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp -3599
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform 1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp -3599
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp -3599
transform 1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp -3599
transform 1 0 12236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp -3599
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp -3599
transform 1 0 12788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform 1 0 11960 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform 1 0 11684 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp -3599
transform 1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform -1 0 11408 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp -3599
transform 1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp -3599
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _092_
timestamp -3599
transform -1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp -3599
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp -3599
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp -3599
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp -3599
transform -1 0 24196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp -3599
transform -1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _098_
timestamp -3599
transform -1 0 24932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _099_
timestamp -3599
transform -1 0 25208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _100_
timestamp -3599
transform -1 0 25668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _101_
timestamp -3599
transform -1 0 26036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp -3599
transform -1 0 26404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _103_
timestamp -3599
transform -1 0 26772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _104_
timestamp -3599
transform -1 0 27048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp -3599
transform 1 0 10304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 17112 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 18860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 15640 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform 1 0 13156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 15640 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 17112 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform 1 0 19780 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 15364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 15824 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform 1 0 17020 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 20884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 19320 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 16560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 19044 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 16008 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 21620 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform -1 0 18308 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform 1 0 12972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform 1 0 16928 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform -1 0 17848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform 1 0 16744 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform 1 0 12788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 19044 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform -1 0 28796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 21528 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 23000 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform -1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform -1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 2576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform -1 0 4048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6
timestamp -3599
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp -3599
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12
timestamp -3599
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18
timestamp -3599
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21
timestamp -3599
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp -3599
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35
timestamp -3599
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp -3599
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp -3599
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp -3599
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47
timestamp -3599
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50
timestamp -3599
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60
timestamp -3599
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp -3599
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp -3599
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75
timestamp -3599
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_78
timestamp -3599
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_88
timestamp -3599
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91
timestamp -3599
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp -3599
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp -3599
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100
timestamp -3599
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103
timestamp -3599
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106
timestamp -3599
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_116
timestamp -3599
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp -3599
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_122
timestamp -3599
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp -3599
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_128
timestamp -3599
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_131
timestamp -3599
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_134
timestamp -3599
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_144
timestamp -3599
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_147
timestamp -3599
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_150
timestamp -3599
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_153
timestamp -3599
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp -3599
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_159
timestamp -3599
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_162
timestamp -3599
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_172
timestamp -3599
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_175
timestamp -3599
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_178
timestamp -3599
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp -3599
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_184
timestamp -3599
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp -3599
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_190
timestamp -3599
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_200
timestamp -3599
transform 1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_203
timestamp -3599
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_206
timestamp -3599
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_209
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_212
timestamp -3599
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_215
timestamp -3599
transform 1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp -3599
transform 1 0 21160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_228
timestamp -3599
transform 1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_231
timestamp -3599
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_234
timestamp -3599
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_237
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_240
timestamp -3599
transform 1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_243
timestamp -3599
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_246
timestamp -3599
transform 1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_256
timestamp -3599
transform 1 0 24656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_259
timestamp -3599
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_262
timestamp -3599
transform 1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_265
timestamp -3599
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_268
timestamp -3599
transform 1 0 25760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_271
timestamp -3599
transform 1 0 26036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_274
timestamp -3599
transform 1 0 26312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_281
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_284
timestamp -3599
transform 1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_287
timestamp -3599
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_290
timestamp -3599
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_293
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp -3599
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_299
timestamp -3599
transform 1 0 28612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_302
timestamp -3599
transform 1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_309
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_312
timestamp -3599
transform 1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_315
timestamp -3599
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_318
timestamp -3599
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_321
timestamp -3599
transform 1 0 30636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6
timestamp -3599
transform 1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_9
timestamp -3599
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_12
timestamp -3599
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_15
timestamp -3599
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_18
timestamp -3599
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_21
timestamp -3599
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_24
timestamp -3599
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp -3599
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_30
timestamp -3599
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_33
timestamp -3599
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_36
timestamp -3599
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_39
timestamp -3599
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_42
timestamp -3599
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_45
timestamp -3599
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_48
timestamp -3599
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -3599
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_60
timestamp -3599
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_63
timestamp -3599
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_66
timestamp -3599
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp -3599
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_72
timestamp -3599
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_75
timestamp -3599
transform 1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp -3599
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp -3599
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_84
timestamp -3599
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_87
timestamp -3599
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_90
timestamp -3599
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_93
timestamp -3599
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_96
timestamp -3599
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_99
timestamp -3599
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp -3599
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_108
timestamp -3599
transform 1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_116
timestamp -3599
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp -3599
transform 1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_122
timestamp -3599
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp -3599
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_128
timestamp -3599
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_131
timestamp -3599
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_134
timestamp -3599
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_137
timestamp -3599
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_140
timestamp -3599
transform 1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp -3599
transform 1 0 14260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_146
timestamp -3599
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_149
timestamp -3599
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp -3599
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_155
timestamp -3599
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_158
timestamp -3599
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_164
timestamp -3599
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_172
timestamp -3599
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_175
timestamp -3599
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_178
timestamp -3599
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_181
timestamp -3599
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp -3599
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_187
timestamp -3599
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_190
timestamp -3599
transform 1 0 18584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_193
timestamp -3599
transform 1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_196
timestamp -3599
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_199
timestamp -3599
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_202
timestamp -3599
transform 1 0 19688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_205
timestamp -3599
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp -3599
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_211
timestamp -3599
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_214
timestamp -3599
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_217
timestamp -3599
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp -3599
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -3599
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_228
timestamp -3599
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_231
timestamp -3599
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_234
timestamp -3599
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_237
timestamp -3599
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_240
timestamp -3599
transform 1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_243
timestamp -3599
transform 1 0 23460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_246
timestamp -3599
transform 1 0 23736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_249
timestamp -3599
transform 1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_252
timestamp -3599
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_255
timestamp -3599
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_258
timestamp -3599
transform 1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_261
timestamp -3599
transform 1 0 25116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_264
timestamp -3599
transform 1 0 25392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_267
timestamp -3599
transform 1 0 25668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_270
timestamp -3599
transform 1 0 25944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_273
timestamp -3599
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_276
timestamp -3599
transform 1 0 26496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -3599
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_284
timestamp -3599
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_287
timestamp -3599
transform 1 0 27508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_290
timestamp -3599
transform 1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_293
timestamp -3599
transform 1 0 28060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_296
timestamp -3599
transform 1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_299
timestamp -3599
transform 1 0 28612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_302
timestamp -3599
transform 1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_305
timestamp -3599
transform 1 0 29164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_308
timestamp -3599
transform 1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_311
timestamp -3599
transform 1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_314
timestamp -3599
transform 1 0 29992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_317
timestamp -3599
transform 1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_320
timestamp -3599
transform 1 0 30544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_323
timestamp -3599
transform 1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_326
timestamp -3599
transform 1 0 31096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_329
timestamp -3599
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_6
timestamp -3599
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_9
timestamp -3599
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_12
timestamp -3599
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_18
timestamp -3599
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_21
timestamp -3599
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_24
timestamp -3599
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp -3599
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_35
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_38
timestamp -3599
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp -3599
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_44
timestamp -3599
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_47
timestamp -3599
transform 1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp -3599
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp -3599
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp -3599
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_59
timestamp -3599
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_62
timestamp -3599
transform 1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_65
timestamp -3599
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp -3599
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_71
timestamp -3599
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_74
timestamp -3599
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_80
timestamp -3599
transform 1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_88
timestamp -3599
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_91
timestamp -3599
transform 1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_94
timestamp -3599
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_97
timestamp -3599
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_104
timestamp -3599
transform 1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp -3599
transform 1 0 10948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_112
timestamp -3599
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_115
timestamp -3599
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_118
timestamp -3599
transform 1 0 11960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_122
timestamp -3599
transform 1 0 12328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_125
timestamp -3599
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_128
timestamp -3599
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_131
timestamp -3599
transform 1 0 13156 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_134
timestamp -3599
transform 1 0 13432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp -3599
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_146
timestamp -3599
transform 1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_149
timestamp -3599
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_152
timestamp -3599
transform 1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_160
timestamp -3599
transform 1 0 15824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_163
timestamp -3599
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_166
timestamp -3599
transform 1 0 16376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_169
timestamp -3599
transform 1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_172
timestamp -3599
transform 1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_175
timestamp -3599
transform 1 0 17204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_178
timestamp -3599
transform 1 0 17480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_185
timestamp -3599
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_188
timestamp -3599
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_191
timestamp -3599
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp -3599
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_200
timestamp -3599
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp -3599
transform 1 0 20240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_213
timestamp -3599
transform 1 0 20700 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp -3599
transform 1 0 21160 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_225
timestamp -3599
transform 1 0 21804 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_228
timestamp -3599
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_231
timestamp -3599
transform 1 0 22356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_234
timestamp -3599
transform 1 0 22632 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_241
timestamp -3599
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_244
timestamp -3599
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_247
timestamp -3599
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp -3599
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_256
timestamp -3599
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_259
timestamp -3599
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_262
timestamp -3599
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_265
timestamp -3599
transform 1 0 25484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_268
timestamp -3599
transform 1 0 25760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_271
timestamp -3599
transform 1 0 26036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_274
timestamp -3599
transform 1 0 26312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_277
timestamp -3599
transform 1 0 26588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_280
timestamp -3599
transform 1 0 26864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_285
timestamp -3599
transform 1 0 27324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_288
timestamp -3599
transform 1 0 27600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_291
timestamp -3599
transform 1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_294
timestamp -3599
transform 1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_297
timestamp -3599
transform 1 0 28428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_300
timestamp -3599
transform 1 0 28704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp -3599
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_309
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_313
timestamp -3599
transform 1 0 29900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_316
timestamp -3599
transform 1 0 30176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_319
timestamp -3599
transform 1 0 30452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_322
timestamp -3599
transform 1 0 30728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_325
timestamp -3599
transform 1 0 31004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_328
timestamp -3599
transform 1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_331
timestamp -3599
transform 1 0 31556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_334
timestamp -3599
transform 1 0 31832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_337
timestamp -3599
transform 1 0 32108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_6
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_9
timestamp -3599
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_12
timestamp -3599
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_18
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_21
timestamp -3599
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_24
timestamp -3599
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp -3599
transform 1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_30
timestamp -3599
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_33
timestamp -3599
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_36
timestamp -3599
transform 1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_39
timestamp -3599
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_42
timestamp -3599
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_45
timestamp -3599
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_48
timestamp -3599
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp -3599
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_60
timestamp -3599
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_63
timestamp -3599
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_66
timestamp -3599
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp -3599
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_73
timestamp -3599
transform 1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_76
timestamp -3599
transform 1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_79
timestamp -3599
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_82
timestamp -3599
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_85
timestamp -3599
transform 1 0 8924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_88
timestamp -3599
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_91
timestamp -3599
transform 1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_94
timestamp -3599
transform 1 0 9752 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_97
timestamp -3599
transform 1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_100
timestamp -3599
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_103
timestamp -3599
transform 1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_106
timestamp -3599
transform 1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp -3599
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_131
timestamp -3599
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_134
timestamp -3599
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_137
timestamp -3599
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_140
timestamp -3599
transform 1 0 13984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_143
timestamp -3599
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_146
timestamp -3599
transform 1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_149
timestamp -3599
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_152
timestamp -3599
transform 1 0 15088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_155
timestamp -3599
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_158
timestamp -3599
transform 1 0 15640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_164
timestamp -3599
transform 1 0 16192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_172
timestamp -3599
transform 1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_175
timestamp -3599
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_178
timestamp -3599
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp -3599
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp -3599
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_187
timestamp -3599
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_190
timestamp -3599
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_193
timestamp -3599
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_196
timestamp -3599
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_199
timestamp -3599
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_202
timestamp -3599
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_205
timestamp -3599
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_208
timestamp -3599
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_211
timestamp -3599
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_214
timestamp -3599
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp -3599
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp -3599
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_228
timestamp -3599
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_231
timestamp -3599
transform 1 0 22356 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_234
timestamp -3599
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_237
timestamp -3599
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_240
timestamp -3599
transform 1 0 23184 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_243
timestamp -3599
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_246
timestamp -3599
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_249
timestamp -3599
transform 1 0 24012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_252
timestamp -3599
transform 1 0 24288 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_255
timestamp -3599
transform 1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_258
timestamp -3599
transform 1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_261
timestamp -3599
transform 1 0 25116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_264
timestamp -3599
transform 1 0 25392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_267
timestamp -3599
transform 1 0 25668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_270
timestamp -3599
transform 1 0 25944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_273
timestamp -3599
transform 1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_276
timestamp -3599
transform 1 0 26496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_281
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_284
timestamp -3599
transform 1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_287
timestamp -3599
transform 1 0 27508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_290
timestamp -3599
transform 1 0 27784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_293
timestamp -3599
transform 1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_296
timestamp -3599
transform 1 0 28336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_299
timestamp -3599
transform 1 0 28612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_302
timestamp -3599
transform 1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_305
timestamp -3599
transform 1 0 29164 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_308
timestamp -3599
transform 1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_311
timestamp -3599
transform 1 0 29716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_314
timestamp -3599
transform 1 0 29992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_317
timestamp -3599
transform 1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_320
timestamp -3599
transform 1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_323
timestamp -3599
transform 1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_326
timestamp -3599
transform 1 0 31096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_329
timestamp -3599
transform 1 0 31372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_332
timestamp -3599
transform 1 0 31648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp -3599
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_6
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp -3599
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_12
timestamp -3599
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_18
timestamp -3599
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_21
timestamp -3599
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_24
timestamp -3599
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp -3599
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_35
timestamp -3599
transform 1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp -3599
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_44
timestamp -3599
transform 1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_47
timestamp -3599
transform 1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_50
timestamp -3599
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp -3599
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_56
timestamp -3599
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_59
timestamp -3599
transform 1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_62
timestamp -3599
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp -3599
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_68
timestamp -3599
transform 1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_71
timestamp -3599
transform 1 0 7636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_74
timestamp -3599
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_80
timestamp -3599
transform 1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_88
timestamp -3599
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_91
timestamp -3599
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_94
timestamp -3599
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_100
timestamp -3599
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_103
timestamp -3599
transform 1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_106
timestamp -3599
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp -3599
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_112
timestamp -3599
transform 1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_115
timestamp -3599
transform 1 0 11684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_120
timestamp -3599
transform 1 0 12144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_123
timestamp -3599
transform 1 0 12420 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_126
timestamp -3599
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_129
timestamp -3599
transform 1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_132
timestamp -3599
transform 1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_135
timestamp -3599
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp -3599
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_144
timestamp -3599
transform 1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_147
timestamp -3599
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp -3599
transform 1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_153
timestamp -3599
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp -3599
transform 1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_159
timestamp -3599
transform 1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_162
timestamp -3599
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp -3599
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_168
timestamp -3599
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_171
timestamp -3599
transform 1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_174
timestamp -3599
transform 1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_177
timestamp -3599
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_180
timestamp -3599
transform 1 0 17664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_183
timestamp -3599
transform 1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_186
timestamp -3599
transform 1 0 18216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_189
timestamp -3599
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_192
timestamp -3599
transform 1 0 18768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_200
timestamp -3599
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_203
timestamp -3599
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_206
timestamp -3599
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp -3599
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_212
timestamp -3599
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_215
timestamp -3599
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_218
timestamp -3599
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp -3599
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_224
timestamp -3599
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_227
timestamp -3599
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_230
timestamp -3599
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_233
timestamp -3599
transform 1 0 22540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_236
timestamp -3599
transform 1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_239
timestamp -3599
transform 1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_242
timestamp -3599
transform 1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_245
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_248
timestamp -3599
transform 1 0 23920 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_256
timestamp -3599
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_259
timestamp -3599
transform 1 0 24932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_262
timestamp -3599
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_265
timestamp -3599
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_268
timestamp -3599
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_271
timestamp -3599
transform 1 0 26036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_274
timestamp -3599
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_277
timestamp -3599
transform 1 0 26588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_280
timestamp -3599
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_283
timestamp -3599
transform 1 0 27140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_286
timestamp -3599
transform 1 0 27416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_289
timestamp -3599
transform 1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_292
timestamp -3599
transform 1 0 27968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_295
timestamp -3599
transform 1 0 28244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp -3599
transform 1 0 28520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_304
timestamp -3599
transform 1 0 29072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_312
timestamp -3599
transform 1 0 29808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_315
timestamp -3599
transform 1 0 30084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_318
timestamp -3599
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_324
timestamp -3599
transform 1 0 30912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_327
timestamp -3599
transform 1 0 31188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_330
timestamp -3599
transform 1 0 31464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp -3599
transform 1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_336
timestamp -3599
transform 1 0 32016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_6
timestamp -3599
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_9
timestamp -3599
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp -3599
transform 1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_18
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_21
timestamp -3599
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp -3599
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp -3599
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_33
timestamp -3599
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_36
timestamp -3599
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_42
timestamp -3599
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_45
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_48
timestamp -3599
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -3599
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_60
timestamp -3599
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_63
timestamp -3599
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_66
timestamp -3599
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_72
timestamp -3599
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp -3599
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_84
timestamp -3599
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_87
timestamp -3599
transform 1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_90
timestamp -3599
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp -3599
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_96
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_99
timestamp -3599
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_102
timestamp -3599
transform 1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_108
timestamp -3599
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_116
timestamp -3599
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp -3599
transform 1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_122
timestamp -3599
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp -3599
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_128
timestamp -3599
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_131
timestamp -3599
transform 1 0 13156 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_134
timestamp -3599
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_137
timestamp -3599
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_140
timestamp -3599
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp -3599
transform 1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_146
timestamp -3599
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp -3599
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_152
timestamp -3599
transform 1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_155
timestamp -3599
transform 1 0 15364 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_158
timestamp -3599
transform 1 0 15640 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_164
timestamp -3599
transform 1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_195
timestamp -3599
transform 1 0 19044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_198
timestamp -3599
transform 1 0 19320 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_201
timestamp -3599
transform 1 0 19596 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_204
timestamp -3599
transform 1 0 19872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_207
timestamp -3599
transform 1 0 20148 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_210
timestamp -3599
transform 1 0 20424 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_213
timestamp -3599
transform 1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_216
timestamp -3599
transform 1 0 20976 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_219
timestamp -3599
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp -3599
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_228
timestamp -3599
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_231
timestamp -3599
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_234
timestamp -3599
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_237
timestamp -3599
transform 1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_240
timestamp -3599
transform 1 0 23184 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_243
timestamp -3599
transform 1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_246
timestamp -3599
transform 1 0 23736 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_249
timestamp -3599
transform 1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_252
timestamp -3599
transform 1 0 24288 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_255
timestamp -3599
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_258
timestamp -3599
transform 1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_261
timestamp -3599
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_264
timestamp -3599
transform 1 0 25392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_267
timestamp -3599
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_270
timestamp -3599
transform 1 0 25944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_276
timestamp -3599
transform 1 0 26496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_284
timestamp -3599
transform 1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_287
timestamp -3599
transform 1 0 27508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_290
timestamp -3599
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_293
timestamp -3599
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_296
timestamp -3599
transform 1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_299
timestamp -3599
transform 1 0 28612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_302
timestamp -3599
transform 1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_305
timestamp -3599
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_308
timestamp -3599
transform 1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_311
timestamp -3599
transform 1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_314
timestamp -3599
transform 1 0 29992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_317
timestamp -3599
transform 1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_320
timestamp -3599
transform 1 0 30544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_323
timestamp -3599
transform 1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_326
timestamp -3599
transform 1 0 31096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_329
timestamp -3599
transform 1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_332
timestamp -3599
transform 1 0 31648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp -3599
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_6
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_9
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_12
timestamp -3599
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_15
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_18
timestamp -3599
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_21
timestamp -3599
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_24
timestamp -3599
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp -3599
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_38
timestamp -3599
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_44
timestamp -3599
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_47
timestamp -3599
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_50
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp -3599
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp -3599
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_59
timestamp -3599
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_62
timestamp -3599
transform 1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_70
timestamp -3599
transform 1 0 7544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_73
timestamp -3599
transform 1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_76
timestamp -3599
transform 1 0 8096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_79
timestamp -3599
transform 1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp -3599
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_88
timestamp -3599
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_91
timestamp -3599
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_94
timestamp -3599
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_97
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_100
timestamp -3599
transform 1 0 10304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_103
timestamp -3599
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_106
timestamp -3599
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_109
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_112
timestamp -3599
transform 1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_115
timestamp -3599
transform 1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_118
timestamp -3599
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp -3599
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_124
timestamp -3599
transform 1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_127
timestamp -3599
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_130
timestamp -3599
transform 1 0 13064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_136
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_144
timestamp -3599
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_147
timestamp -3599
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp -3599
transform 1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_153
timestamp -3599
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_161
timestamp -3599
transform 1 0 15916 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_164
timestamp -3599
transform 1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_167
timestamp -3599
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_182
timestamp -3599
transform 1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_185
timestamp -3599
transform 1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_188
timestamp -3599
transform 1 0 18400 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_191
timestamp -3599
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp -3599
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_200
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_203
timestamp -3599
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_206
timestamp -3599
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_212
timestamp -3599
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp -3599
transform 1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_218
timestamp -3599
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_221
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_224
timestamp -3599
transform 1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_227
timestamp -3599
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_230
timestamp -3599
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_233
timestamp -3599
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_236
timestamp -3599
transform 1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_239
timestamp -3599
transform 1 0 23092 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_242
timestamp -3599
transform 1 0 23368 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_245
timestamp -3599
transform 1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_248
timestamp -3599
transform 1 0 23920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -3599
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_256
timestamp -3599
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_259
timestamp -3599
transform 1 0 24932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_262
timestamp -3599
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_268
timestamp -3599
transform 1 0 25760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_271
timestamp -3599
transform 1 0 26036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_274
timestamp -3599
transform 1 0 26312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_277
timestamp -3599
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_280
timestamp -3599
transform 1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_283
timestamp -3599
transform 1 0 27140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_286
timestamp -3599
transform 1 0 27416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_289
timestamp -3599
transform 1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_292
timestamp -3599
transform 1 0 27968 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_295
timestamp -3599
transform 1 0 28244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_298
timestamp -3599
transform 1 0 28520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_301
timestamp -3599
transform 1 0 28796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_304
timestamp -3599
transform 1 0 29072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_312
timestamp -3599
transform 1 0 29808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_315
timestamp -3599
transform 1 0 30084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_318
timestamp -3599
transform 1 0 30360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_321
timestamp -3599
transform 1 0 30636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_324
timestamp -3599
transform 1 0 30912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_327
timestamp -3599
transform 1 0 31188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_330
timestamp -3599
transform 1 0 31464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_333
timestamp -3599
transform 1 0 31740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_336
timestamp -3599
transform 1 0 32016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_6
timestamp -3599
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_9
timestamp -3599
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_12
timestamp -3599
transform 1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_18
timestamp -3599
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_21
timestamp -3599
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp -3599
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp -3599
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp -3599
transform 1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_46
timestamp -3599
transform 1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_49
timestamp -3599
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_52
timestamp -3599
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_73
timestamp -3599
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_82
timestamp -3599
transform 1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_85
timestamp -3599
transform 1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_88
timestamp -3599
transform 1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_91
timestamp -3599
transform 1 0 9476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_94
timestamp -3599
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_97
timestamp -3599
transform 1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_100
timestamp -3599
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_103
timestamp -3599
transform 1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_106
timestamp -3599
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp -3599
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_116
timestamp -3599
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp -3599
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp -3599
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_125
timestamp -3599
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_162
timestamp -3599
transform 1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp -3599
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_172
timestamp -3599
transform 1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_175
timestamp -3599
transform 1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_178
timestamp -3599
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp -3599
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_184
timestamp -3599
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_187
timestamp -3599
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_190
timestamp -3599
transform 1 0 18584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_193
timestamp -3599
transform 1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_196
timestamp -3599
transform 1 0 19136 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_199
timestamp -3599
transform 1 0 19412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_202
timestamp -3599
transform 1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_205
timestamp -3599
transform 1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_208
timestamp -3599
transform 1 0 20240 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_211
timestamp -3599
transform 1 0 20516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_214
timestamp -3599
transform 1 0 20792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp -3599
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_220
timestamp -3599
transform 1 0 21344 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_243
timestamp -3599
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_246
timestamp -3599
transform 1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_249
timestamp -3599
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_252
timestamp -3599
transform 1 0 24288 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_255
timestamp -3599
transform 1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_258
timestamp -3599
transform 1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_261
timestamp -3599
transform 1 0 25116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_264
timestamp -3599
transform 1 0 25392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_267
timestamp -3599
transform 1 0 25668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_270
timestamp -3599
transform 1 0 25944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_273
timestamp -3599
transform 1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_276
timestamp -3599
transform 1 0 26496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -3599
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_284
timestamp -3599
transform 1 0 27232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_287
timestamp -3599
transform 1 0 27508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_290
timestamp -3599
transform 1 0 27784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_296
timestamp -3599
transform 1 0 28336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_299
timestamp -3599
transform 1 0 28612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_302
timestamp -3599
transform 1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_305
timestamp -3599
transform 1 0 29164 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_308
timestamp -3599
transform 1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_311
timestamp -3599
transform 1 0 29716 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_314
timestamp -3599
transform 1 0 29992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_317
timestamp -3599
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_320
timestamp -3599
transform 1 0 30544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_323
timestamp -3599
transform 1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_326
timestamp -3599
transform 1 0 31096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_332
timestamp -3599
transform 1 0 31648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_6
timestamp -3599
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_9
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_12
timestamp -3599
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp -3599
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_18
timestamp -3599
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_21
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_35
timestamp -3599
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp -3599
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp -3599
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_47
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_50
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp -3599
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_56
timestamp -3599
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_59
timestamp -3599
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_69
timestamp -3599
transform 1 0 7452 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_72
timestamp -3599
transform 1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_75
timestamp -3599
transform 1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_78
timestamp -3599
transform 1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp -3599
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_88
timestamp -3599
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_91
timestamp -3599
transform 1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_94
timestamp -3599
transform 1 0 9752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp -3599
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_100
timestamp -3599
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_103
timestamp -3599
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_106
timestamp -3599
transform 1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_109
timestamp -3599
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_112
timestamp -3599
transform 1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_115
timestamp -3599
transform 1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_118
timestamp -3599
transform 1 0 11960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_125
timestamp -3599
transform 1 0 12604 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_128
timestamp -3599
transform 1 0 12880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_131
timestamp -3599
transform 1 0 13156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_134
timestamp -3599
transform 1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp -3599
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_144
timestamp -3599
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_147
timestamp -3599
transform 1 0 14628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp -3599
transform 1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_156
timestamp -3599
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_159
timestamp -3599
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_162
timestamp -3599
transform 1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp -3599
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp -3599
transform 1 0 16560 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_171
timestamp -3599
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_174
timestamp -3599
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_180
timestamp -3599
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_183
timestamp -3599
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_186
timestamp -3599
transform 1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_192
timestamp -3599
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_200
timestamp -3599
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_203
timestamp -3599
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_206
timestamp -3599
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp -3599
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_212
timestamp -3599
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_215
timestamp -3599
transform 1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_218
timestamp -3599
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_221
timestamp -3599
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_224
timestamp -3599
transform 1 0 21712 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_227
timestamp -3599
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_230
timestamp -3599
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_233
timestamp -3599
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_236
timestamp -3599
transform 1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_239
timestamp -3599
transform 1 0 23092 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_242
timestamp -3599
transform 1 0 23368 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_245
timestamp -3599
transform 1 0 23644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_262
timestamp -3599
transform 1 0 25208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_267
timestamp -3599
transform 1 0 25668 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_271
timestamp -3599
transform 1 0 26036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_275
timestamp -3599
transform 1 0 26404 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_282
timestamp -3599
transform 1 0 27048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_285
timestamp -3599
transform 1 0 27324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_288
timestamp -3599
transform 1 0 27600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_291
timestamp -3599
transform 1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_294
timestamp -3599
transform 1 0 28152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_297
timestamp -3599
transform 1 0 28428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_300
timestamp -3599
transform 1 0 28704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_303
timestamp -3599
transform 1 0 28980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_312
timestamp -3599
transform 1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_315
timestamp -3599
transform 1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_318
timestamp -3599
transform 1 0 30360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_321
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_324
timestamp -3599
transform 1 0 30912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_327
timestamp -3599
transform 1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_330
timestamp -3599
transform 1 0 31464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_333
timestamp -3599
transform 1 0 31740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_336
timestamp -3599
transform 1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6
timestamp -3599
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_9
timestamp -3599
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_25
timestamp -3599
transform 1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_28
timestamp -3599
transform 1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_31
timestamp -3599
transform 1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_34
timestamp -3599
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_37
timestamp -3599
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_40
timestamp -3599
transform 1 0 4784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_43
timestamp -3599
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_46
timestamp -3599
transform 1 0 5336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_49
timestamp -3599
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_52
timestamp -3599
transform 1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_60
timestamp -3599
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_63
timestamp -3599
transform 1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_70
timestamp -3599
transform 1 0 7544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_73
timestamp -3599
transform 1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_76
timestamp -3599
transform 1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_79
timestamp -3599
transform 1 0 8372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_82
timestamp -3599
transform 1 0 8648 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_85
timestamp -3599
transform 1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_92
timestamp -3599
transform 1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_98
timestamp -3599
transform 1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_101
timestamp -3599
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_104
timestamp -3599
transform 1 0 10672 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_107
timestamp -3599
transform 1 0 10948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_130
timestamp -3599
transform 1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_133
timestamp -3599
transform 1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_136
timestamp -3599
transform 1 0 13616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_139
timestamp -3599
transform 1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_142
timestamp -3599
transform 1 0 14168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_145
timestamp -3599
transform 1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_148
timestamp -3599
transform 1 0 14720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_151
timestamp -3599
transform 1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_154
timestamp -3599
transform 1 0 15272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_157
timestamp -3599
transform 1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_160
timestamp -3599
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_163
timestamp -3599
transform 1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_178
timestamp -3599
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_181
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp -3599
transform 1 0 18032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_195
timestamp -3599
transform 1 0 19044 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_204
timestamp -3599
transform 1 0 19872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp -3599
transform 1 0 20240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_228
timestamp -3599
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_231
timestamp -3599
transform 1 0 22356 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_234
timestamp -3599
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_237
timestamp -3599
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_240
timestamp -3599
transform 1 0 23184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_243
timestamp -3599
transform 1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_246
timestamp -3599
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_249
timestamp -3599
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_252
timestamp -3599
transform 1 0 24288 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_255
timestamp -3599
transform 1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_258
timestamp -3599
transform 1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_261
timestamp -3599
transform 1 0 25116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_264
timestamp -3599
transform 1 0 25392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_267
timestamp -3599
transform 1 0 25668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_270
timestamp -3599
transform 1 0 25944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_273
timestamp -3599
transform 1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_276
timestamp -3599
transform 1 0 26496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -3599
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_284
timestamp -3599
transform 1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_287
timestamp -3599
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_293
timestamp -3599
transform 1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_308
timestamp -3599
transform 1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_320
timestamp -3599
transform 1 0 30544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_324
timestamp -3599
transform 1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_327
timestamp -3599
transform 1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_330
timestamp -3599
transform 1 0 31464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp -3599
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_6
timestamp -3599
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_9
timestamp -3599
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_12
timestamp -3599
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_18
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_24
timestamp -3599
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp -3599
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_35
timestamp -3599
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_38
timestamp -3599
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_44
timestamp -3599
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_47
timestamp -3599
transform 1 0 5428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_148
timestamp -3599
transform 1 0 14720 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_151
timestamp -3599
transform 1 0 14996 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp -3599
transform 1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_157
timestamp -3599
transform 1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_160
timestamp -3599
transform 1 0 15824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_163
timestamp -3599
transform 1 0 16100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_166
timestamp -3599
transform 1 0 16376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_169
timestamp -3599
transform 1 0 16652 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_172
timestamp -3599
transform 1 0 16928 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_175
timestamp -3599
transform 1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_178
timestamp -3599
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_181
timestamp -3599
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_184
timestamp -3599
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_187
timestamp -3599
transform 1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_190
timestamp -3599
transform 1 0 18584 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp -3599
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_200
timestamp -3599
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_203
timestamp -3599
transform 1 0 19780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_206
timestamp -3599
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp -3599
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_212
timestamp -3599
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp -3599
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_218
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_221
timestamp -3599
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_224
timestamp -3599
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_227
timestamp -3599
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp -3599
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_233
timestamp -3599
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_236
timestamp -3599
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_239
timestamp -3599
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_242
timestamp -3599
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_245
timestamp -3599
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_248
timestamp -3599
transform 1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_256
timestamp -3599
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_259
timestamp -3599
transform 1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_262
timestamp -3599
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_265
timestamp -3599
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_268
timestamp -3599
transform 1 0 25760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp -3599
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_312
timestamp -3599
transform 1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_315
timestamp -3599
transform 1 0 30084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_318
timestamp -3599
transform 1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_321
timestamp -3599
transform 1 0 30636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_324
timestamp -3599
transform 1 0 30912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_327
timestamp -3599
transform 1 0 31188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_330
timestamp -3599
transform 1 0 31464 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_6
timestamp -3599
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_9
timestamp -3599
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_12
timestamp -3599
transform 1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_15
timestamp -3599
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_18
timestamp -3599
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_21
timestamp -3599
transform 1 0 3036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_24
timestamp -3599
transform 1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp -3599
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_32
timestamp -3599
transform 1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_35
timestamp -3599
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_38
timestamp -3599
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_163
timestamp -3599
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp -3599
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_172
timestamp -3599
transform 1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_175
timestamp -3599
transform 1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_178
timestamp -3599
transform 1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_181
timestamp -3599
transform 1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_184
timestamp -3599
transform 1 0 18032 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_187
timestamp -3599
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_190
timestamp -3599
transform 1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_193
timestamp -3599
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_200
timestamp -3599
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_203
timestamp -3599
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_206
timestamp -3599
transform 1 0 20056 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_209
timestamp -3599
transform 1 0 20332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_212
timestamp -3599
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_215
timestamp -3599
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_218
timestamp -3599
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp -3599
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_228
timestamp -3599
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_231
timestamp -3599
transform 1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_234
timestamp -3599
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_237
timestamp -3599
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_240
timestamp -3599
transform 1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_243
timestamp -3599
transform 1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_246
timestamp -3599
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_249
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_253
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_256
timestamp -3599
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp -3599
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp -3599
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_313
timestamp -3599
transform 1 0 29900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_316
timestamp -3599
transform 1 0 30176 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_319
timestamp -3599
transform 1 0 30452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_322
timestamp -3599
transform 1 0 30728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_325
timestamp -3599
transform 1 0 31004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 32292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 32660 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 32292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 32660 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 32292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 32660 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 32292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 32660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 32292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 32660 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 31280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 32292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 32660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 32660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 32292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 32660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 32660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 32292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 31280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 31924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 32292 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 30912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 32292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 32660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 32292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 32660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform 1 0 25208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform -1 0 27416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform -1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform -1 0 27784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform -1 0 28796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 27784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform -1 0 29164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform -1 0 28520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform -1 0 28888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform -1 0 29256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform -1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform 1 0 25576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 25944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 26312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform 1 0 26312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform 1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 27048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform -1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 5888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 6624 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 6624 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform -1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 9200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform -1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform -1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform -1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform -1 0 10120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform -1 0 9936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform -1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform -1 0 10672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform -1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform -1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 13248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 13984 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform -1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 33304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 33304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 33304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 33304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 33304 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 33304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 33304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 33304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 33304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 33304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_term_single_106
timestamp -3599
transform -1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_36
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_42
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_43
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_44
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_48
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_49
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_50
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_51
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_54
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_55
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_57
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_58
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_60
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_61
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_62
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_63
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_64
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_65
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_66
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_67
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_68
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_69
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_70
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_71
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_72
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_73
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_74
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_75
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_76
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_77
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_79
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_80
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_81
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_82
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_84
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_85
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_89
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_92
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_94
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_97
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_101
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_102
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_103
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_104
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_105
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_106
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_107
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 15198 11096 15254 11152 0 FreeSans 224 0 0 0 Co
port 0 nsew signal output
flabel metal3 s 0 1096 120 1216 0 FreeSans 480 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 34288 1096 34408 1216 0 FreeSans 480 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 34288 3816 34408 3936 0 FreeSans 480 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 34288 4088 34408 4208 0 FreeSans 480 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 34288 4360 34408 4480 0 FreeSans 480 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 34288 4632 34408 4752 0 FreeSans 480 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 34288 4904 34408 5024 0 FreeSans 480 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 34288 5176 34408 5296 0 FreeSans 480 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 34288 5448 34408 5568 0 FreeSans 480 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 34288 5720 34408 5840 0 FreeSans 480 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 34288 5992 34408 6112 0 FreeSans 480 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 34288 6264 34408 6384 0 FreeSans 480 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 34288 1368 34408 1488 0 FreeSans 480 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 34288 6536 34408 6656 0 FreeSans 480 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 34288 6808 34408 6928 0 FreeSans 480 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 34288 7080 34408 7200 0 FreeSans 480 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 34288 7352 34408 7472 0 FreeSans 480 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 34288 7624 34408 7744 0 FreeSans 480 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 34288 7896 34408 8016 0 FreeSans 480 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 34288 8168 34408 8288 0 FreeSans 480 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 34288 8440 34408 8560 0 FreeSans 480 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 34288 8712 34408 8832 0 FreeSans 480 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 34288 8984 34408 9104 0 FreeSans 480 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 34288 1640 34408 1760 0 FreeSans 480 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 34288 9256 34408 9376 0 FreeSans 480 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 34288 9528 34408 9648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 34288 1912 34408 2032 0 FreeSans 480 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 34288 2184 34408 2304 0 FreeSans 480 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 34288 2456 34408 2576 0 FreeSans 480 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 34288 2728 34408 2848 0 FreeSans 480 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 34288 3000 34408 3120 0 FreeSans 480 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 34288 3272 34408 3392 0 FreeSans 480 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 34288 3544 34408 3664 0 FreeSans 480 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 3054 0 3110 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 18694 0 18750 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 20258 0 20314 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 21822 0 21878 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 23386 0 23442 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 24950 0 25006 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 26514 0 26570 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 28078 0 28134 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 29642 0 29698 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 31206 0 31262 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 32770 0 32826 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 4618 0 4674 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 6182 0 6238 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 7746 0 7802 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 9310 0 9366 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 10874 0 10930 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 12438 0 12494 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 14002 0 14058 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 15566 0 15622 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 17130 0 17186 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 25134 11096 25190 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 26974 11096 27030 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 27158 11096 27214 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 27342 11096 27398 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 27526 11096 27582 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 27710 11096 27766 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 27894 11096 27950 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 28078 11096 28134 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 28262 11096 28318 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 28446 11096 28502 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 28630 11096 28686 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 25318 11096 25374 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 25502 11096 25558 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 25686 11096 25742 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 25870 11096 25926 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 26054 11096 26110 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 26238 11096 26294 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 26422 11096 26478 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 26606 11096 26662 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 26790 11096 26846 11152 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 5630 11096 5686 11152 0 FreeSans 224 0 0 0 N1BEG[0]
port 105 nsew signal output
flabel metal2 s 5814 11096 5870 11152 0 FreeSans 224 0 0 0 N1BEG[1]
port 106 nsew signal output
flabel metal2 s 5998 11096 6054 11152 0 FreeSans 224 0 0 0 N1BEG[2]
port 107 nsew signal output
flabel metal2 s 6182 11096 6238 11152 0 FreeSans 224 0 0 0 N1BEG[3]
port 108 nsew signal output
flabel metal2 s 6366 11096 6422 11152 0 FreeSans 224 0 0 0 N2BEG[0]
port 109 nsew signal output
flabel metal2 s 6550 11096 6606 11152 0 FreeSans 224 0 0 0 N2BEG[1]
port 110 nsew signal output
flabel metal2 s 6734 11096 6790 11152 0 FreeSans 224 0 0 0 N2BEG[2]
port 111 nsew signal output
flabel metal2 s 6918 11096 6974 11152 0 FreeSans 224 0 0 0 N2BEG[3]
port 112 nsew signal output
flabel metal2 s 7102 11096 7158 11152 0 FreeSans 224 0 0 0 N2BEG[4]
port 113 nsew signal output
flabel metal2 s 7286 11096 7342 11152 0 FreeSans 224 0 0 0 N2BEG[5]
port 114 nsew signal output
flabel metal2 s 7470 11096 7526 11152 0 FreeSans 224 0 0 0 N2BEG[6]
port 115 nsew signal output
flabel metal2 s 7654 11096 7710 11152 0 FreeSans 224 0 0 0 N2BEG[7]
port 116 nsew signal output
flabel metal2 s 7838 11096 7894 11152 0 FreeSans 224 0 0 0 N2BEGb[0]
port 117 nsew signal output
flabel metal2 s 8022 11096 8078 11152 0 FreeSans 224 0 0 0 N2BEGb[1]
port 118 nsew signal output
flabel metal2 s 8206 11096 8262 11152 0 FreeSans 224 0 0 0 N2BEGb[2]
port 119 nsew signal output
flabel metal2 s 8390 11096 8446 11152 0 FreeSans 224 0 0 0 N2BEGb[3]
port 120 nsew signal output
flabel metal2 s 8574 11096 8630 11152 0 FreeSans 224 0 0 0 N2BEGb[4]
port 121 nsew signal output
flabel metal2 s 8758 11096 8814 11152 0 FreeSans 224 0 0 0 N2BEGb[5]
port 122 nsew signal output
flabel metal2 s 8942 11096 8998 11152 0 FreeSans 224 0 0 0 N2BEGb[6]
port 123 nsew signal output
flabel metal2 s 9126 11096 9182 11152 0 FreeSans 224 0 0 0 N2BEGb[7]
port 124 nsew signal output
flabel metal2 s 9310 11096 9366 11152 0 FreeSans 224 0 0 0 N4BEG[0]
port 125 nsew signal output
flabel metal2 s 11150 11096 11206 11152 0 FreeSans 224 0 0 0 N4BEG[10]
port 126 nsew signal output
flabel metal2 s 11334 11096 11390 11152 0 FreeSans 224 0 0 0 N4BEG[11]
port 127 nsew signal output
flabel metal2 s 11518 11096 11574 11152 0 FreeSans 224 0 0 0 N4BEG[12]
port 128 nsew signal output
flabel metal2 s 11702 11096 11758 11152 0 FreeSans 224 0 0 0 N4BEG[13]
port 129 nsew signal output
flabel metal2 s 11886 11096 11942 11152 0 FreeSans 224 0 0 0 N4BEG[14]
port 130 nsew signal output
flabel metal2 s 12070 11096 12126 11152 0 FreeSans 224 0 0 0 N4BEG[15]
port 131 nsew signal output
flabel metal2 s 9494 11096 9550 11152 0 FreeSans 224 0 0 0 N4BEG[1]
port 132 nsew signal output
flabel metal2 s 9678 11096 9734 11152 0 FreeSans 224 0 0 0 N4BEG[2]
port 133 nsew signal output
flabel metal2 s 9862 11096 9918 11152 0 FreeSans 224 0 0 0 N4BEG[3]
port 134 nsew signal output
flabel metal2 s 10046 11096 10102 11152 0 FreeSans 224 0 0 0 N4BEG[4]
port 135 nsew signal output
flabel metal2 s 10230 11096 10286 11152 0 FreeSans 224 0 0 0 N4BEG[5]
port 136 nsew signal output
flabel metal2 s 10414 11096 10470 11152 0 FreeSans 224 0 0 0 N4BEG[6]
port 137 nsew signal output
flabel metal2 s 10598 11096 10654 11152 0 FreeSans 224 0 0 0 N4BEG[7]
port 138 nsew signal output
flabel metal2 s 10782 11096 10838 11152 0 FreeSans 224 0 0 0 N4BEG[8]
port 139 nsew signal output
flabel metal2 s 10966 11096 11022 11152 0 FreeSans 224 0 0 0 N4BEG[9]
port 140 nsew signal output
flabel metal2 s 12254 11096 12310 11152 0 FreeSans 224 0 0 0 NN4BEG[0]
port 141 nsew signal output
flabel metal2 s 14094 11096 14150 11152 0 FreeSans 224 0 0 0 NN4BEG[10]
port 142 nsew signal output
flabel metal2 s 14278 11096 14334 11152 0 FreeSans 224 0 0 0 NN4BEG[11]
port 143 nsew signal output
flabel metal2 s 14462 11096 14518 11152 0 FreeSans 224 0 0 0 NN4BEG[12]
port 144 nsew signal output
flabel metal2 s 14646 11096 14702 11152 0 FreeSans 224 0 0 0 NN4BEG[13]
port 145 nsew signal output
flabel metal2 s 14830 11096 14886 11152 0 FreeSans 224 0 0 0 NN4BEG[14]
port 146 nsew signal output
flabel metal2 s 15014 11096 15070 11152 0 FreeSans 224 0 0 0 NN4BEG[15]
port 147 nsew signal output
flabel metal2 s 12438 11096 12494 11152 0 FreeSans 224 0 0 0 NN4BEG[1]
port 148 nsew signal output
flabel metal2 s 12622 11096 12678 11152 0 FreeSans 224 0 0 0 NN4BEG[2]
port 149 nsew signal output
flabel metal2 s 12806 11096 12862 11152 0 FreeSans 224 0 0 0 NN4BEG[3]
port 150 nsew signal output
flabel metal2 s 12990 11096 13046 11152 0 FreeSans 224 0 0 0 NN4BEG[4]
port 151 nsew signal output
flabel metal2 s 13174 11096 13230 11152 0 FreeSans 224 0 0 0 NN4BEG[5]
port 152 nsew signal output
flabel metal2 s 13358 11096 13414 11152 0 FreeSans 224 0 0 0 NN4BEG[6]
port 153 nsew signal output
flabel metal2 s 13542 11096 13598 11152 0 FreeSans 224 0 0 0 NN4BEG[7]
port 154 nsew signal output
flabel metal2 s 13726 11096 13782 11152 0 FreeSans 224 0 0 0 NN4BEG[8]
port 155 nsew signal output
flabel metal2 s 13910 11096 13966 11152 0 FreeSans 224 0 0 0 NN4BEG[9]
port 156 nsew signal output
flabel metal2 s 15382 11096 15438 11152 0 FreeSans 224 0 0 0 S1END[0]
port 157 nsew signal input
flabel metal2 s 15566 11096 15622 11152 0 FreeSans 224 0 0 0 S1END[1]
port 158 nsew signal input
flabel metal2 s 15750 11096 15806 11152 0 FreeSans 224 0 0 0 S1END[2]
port 159 nsew signal input
flabel metal2 s 15934 11096 15990 11152 0 FreeSans 224 0 0 0 S1END[3]
port 160 nsew signal input
flabel metal2 s 17590 11096 17646 11152 0 FreeSans 224 0 0 0 S2END[0]
port 161 nsew signal input
flabel metal2 s 17774 11096 17830 11152 0 FreeSans 224 0 0 0 S2END[1]
port 162 nsew signal input
flabel metal2 s 17958 11096 18014 11152 0 FreeSans 224 0 0 0 S2END[2]
port 163 nsew signal input
flabel metal2 s 18142 11096 18198 11152 0 FreeSans 224 0 0 0 S2END[3]
port 164 nsew signal input
flabel metal2 s 18326 11096 18382 11152 0 FreeSans 224 0 0 0 S2END[4]
port 165 nsew signal input
flabel metal2 s 18510 11096 18566 11152 0 FreeSans 224 0 0 0 S2END[5]
port 166 nsew signal input
flabel metal2 s 18694 11096 18750 11152 0 FreeSans 224 0 0 0 S2END[6]
port 167 nsew signal input
flabel metal2 s 18878 11096 18934 11152 0 FreeSans 224 0 0 0 S2END[7]
port 168 nsew signal input
flabel metal2 s 16118 11096 16174 11152 0 FreeSans 224 0 0 0 S2MID[0]
port 169 nsew signal input
flabel metal2 s 16302 11096 16358 11152 0 FreeSans 224 0 0 0 S2MID[1]
port 170 nsew signal input
flabel metal2 s 16486 11096 16542 11152 0 FreeSans 224 0 0 0 S2MID[2]
port 171 nsew signal input
flabel metal2 s 16670 11096 16726 11152 0 FreeSans 224 0 0 0 S2MID[3]
port 172 nsew signal input
flabel metal2 s 16854 11096 16910 11152 0 FreeSans 224 0 0 0 S2MID[4]
port 173 nsew signal input
flabel metal2 s 17038 11096 17094 11152 0 FreeSans 224 0 0 0 S2MID[5]
port 174 nsew signal input
flabel metal2 s 17222 11096 17278 11152 0 FreeSans 224 0 0 0 S2MID[6]
port 175 nsew signal input
flabel metal2 s 17406 11096 17462 11152 0 FreeSans 224 0 0 0 S2MID[7]
port 176 nsew signal input
flabel metal2 s 19062 11096 19118 11152 0 FreeSans 224 0 0 0 S4END[0]
port 177 nsew signal input
flabel metal2 s 20902 11096 20958 11152 0 FreeSans 224 0 0 0 S4END[10]
port 178 nsew signal input
flabel metal2 s 21086 11096 21142 11152 0 FreeSans 224 0 0 0 S4END[11]
port 179 nsew signal input
flabel metal2 s 21270 11096 21326 11152 0 FreeSans 224 0 0 0 S4END[12]
port 180 nsew signal input
flabel metal2 s 21454 11096 21510 11152 0 FreeSans 224 0 0 0 S4END[13]
port 181 nsew signal input
flabel metal2 s 21638 11096 21694 11152 0 FreeSans 224 0 0 0 S4END[14]
port 182 nsew signal input
flabel metal2 s 21822 11096 21878 11152 0 FreeSans 224 0 0 0 S4END[15]
port 183 nsew signal input
flabel metal2 s 19246 11096 19302 11152 0 FreeSans 224 0 0 0 S4END[1]
port 184 nsew signal input
flabel metal2 s 19430 11096 19486 11152 0 FreeSans 224 0 0 0 S4END[2]
port 185 nsew signal input
flabel metal2 s 19614 11096 19670 11152 0 FreeSans 224 0 0 0 S4END[3]
port 186 nsew signal input
flabel metal2 s 19798 11096 19854 11152 0 FreeSans 224 0 0 0 S4END[4]
port 187 nsew signal input
flabel metal2 s 19982 11096 20038 11152 0 FreeSans 224 0 0 0 S4END[5]
port 188 nsew signal input
flabel metal2 s 20166 11096 20222 11152 0 FreeSans 224 0 0 0 S4END[6]
port 189 nsew signal input
flabel metal2 s 20350 11096 20406 11152 0 FreeSans 224 0 0 0 S4END[7]
port 190 nsew signal input
flabel metal2 s 20534 11096 20590 11152 0 FreeSans 224 0 0 0 S4END[8]
port 191 nsew signal input
flabel metal2 s 20718 11096 20774 11152 0 FreeSans 224 0 0 0 S4END[9]
port 192 nsew signal input
flabel metal2 s 22006 11096 22062 11152 0 FreeSans 224 0 0 0 SS4END[0]
port 193 nsew signal input
flabel metal2 s 23846 11096 23902 11152 0 FreeSans 224 0 0 0 SS4END[10]
port 194 nsew signal input
flabel metal2 s 24030 11096 24086 11152 0 FreeSans 224 0 0 0 SS4END[11]
port 195 nsew signal input
flabel metal2 s 24214 11096 24270 11152 0 FreeSans 224 0 0 0 SS4END[12]
port 196 nsew signal input
flabel metal2 s 24398 11096 24454 11152 0 FreeSans 224 0 0 0 SS4END[13]
port 197 nsew signal input
flabel metal2 s 24582 11096 24638 11152 0 FreeSans 224 0 0 0 SS4END[14]
port 198 nsew signal input
flabel metal2 s 24766 11096 24822 11152 0 FreeSans 224 0 0 0 SS4END[15]
port 199 nsew signal input
flabel metal2 s 22190 11096 22246 11152 0 FreeSans 224 0 0 0 SS4END[1]
port 200 nsew signal input
flabel metal2 s 22374 11096 22430 11152 0 FreeSans 224 0 0 0 SS4END[2]
port 201 nsew signal input
flabel metal2 s 22558 11096 22614 11152 0 FreeSans 224 0 0 0 SS4END[3]
port 202 nsew signal input
flabel metal2 s 22742 11096 22798 11152 0 FreeSans 224 0 0 0 SS4END[4]
port 203 nsew signal input
flabel metal2 s 22926 11096 22982 11152 0 FreeSans 224 0 0 0 SS4END[5]
port 204 nsew signal input
flabel metal2 s 23110 11096 23166 11152 0 FreeSans 224 0 0 0 SS4END[6]
port 205 nsew signal input
flabel metal2 s 23294 11096 23350 11152 0 FreeSans 224 0 0 0 SS4END[7]
port 206 nsew signal input
flabel metal2 s 23478 11096 23534 11152 0 FreeSans 224 0 0 0 SS4END[8]
port 207 nsew signal input
flabel metal2 s 23662 11096 23718 11152 0 FreeSans 224 0 0 0 SS4END[9]
port 208 nsew signal input
flabel metal2 s 1490 0 1546 56 0 FreeSans 224 0 0 0 UserCLK
port 209 nsew signal input
flabel metal2 s 24950 11096 25006 11152 0 FreeSans 224 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal4 s 3004 0 3324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 3004 11092 3324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 9004 11092 9324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 15004 11092 15324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 21004 11092 21324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 27004 11092 27324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11152 0 FreeSans 1920 90 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 33004 11092 33324 11152 0 FreeSans 480 0 0 0 VGND
port 211 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 1944 11092 2264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 0 8264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 7944 11092 8264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 0 14264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 13944 11092 14264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 0 20264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 19944 11092 20264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 0 26264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 25944 11092 26264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 0 32264 11152 0 FreeSans 1920 90 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
flabel metal4 s 31944 11092 32264 11152 0 FreeSans 480 0 0 0 VPWR
port 212 nsew power bidirectional
rlabel metal1 17214 8704 17214 8704 0 VGND
rlabel metal1 17204 8160 17204 8160 0 VPWR
rlabel metal3 5542 1156 5542 1156 0 FrameData[0]
rlabel metal3 919 3876 919 3876 0 FrameData[10]
rlabel metal2 18170 4675 18170 4675 0 FrameData[11]
rlabel metal2 15502 5049 15502 5049 0 FrameData[12]
rlabel metal2 2898 4624 2898 4624 0 FrameData[13]
rlabel metal3 919 4964 919 4964 0 FrameData[14]
rlabel metal1 16744 5610 16744 5610 0 FrameData[15]
rlabel metal1 19734 3706 19734 3706 0 FrameData[16]
rlabel metal2 15410 3944 15410 3944 0 FrameData[17]
rlabel metal3 919 6052 919 6052 0 FrameData[18]
rlabel metal2 16790 4318 16790 4318 0 FrameData[19]
rlabel metal3 7888 1428 7888 1428 0 FrameData[1]
rlabel metal2 17894 4114 17894 4114 0 FrameData[20]
rlabel metal1 12006 2346 12006 2346 0 FrameData[21]
rlabel metal3 919 7140 919 7140 0 FrameData[22]
rlabel metal3 206 7412 206 7412 0 FrameData[23]
rlabel metal3 712 7684 712 7684 0 FrameData[24]
rlabel metal3 735 7956 735 7956 0 FrameData[25]
rlabel metal3 574 8228 574 8228 0 FrameData[26]
rlabel metal1 18492 7174 18492 7174 0 FrameData[27]
rlabel metal2 16422 8347 16422 8347 0 FrameData[28]
rlabel metal2 18630 7667 18630 7667 0 FrameData[29]
rlabel metal3 6876 1700 6876 1700 0 FrameData[2]
rlabel via2 21206 7395 21206 7395 0 FrameData[30]
rlabel via2 18170 7259 18170 7259 0 FrameData[31]
rlabel metal3 6554 1972 6554 1972 0 FrameData[3]
rlabel metal3 1471 2244 1471 2244 0 FrameData[4]
rlabel metal3 8371 2516 8371 2516 0 FrameData[5]
rlabel metal3 919 2788 919 2788 0 FrameData[6]
rlabel metal1 15686 4998 15686 4998 0 FrameData[7]
rlabel metal3 1425 3332 1425 3332 0 FrameData[8]
rlabel metal1 18354 5202 18354 5202 0 FrameData[9]
rlabel metal3 33098 1156 33098 1156 0 FrameData_O[0]
rlabel metal3 33420 3876 33420 3876 0 FrameData_O[10]
rlabel metal3 33604 4148 33604 4148 0 FrameData_O[11]
rlabel metal3 33880 4420 33880 4420 0 FrameData_O[12]
rlabel metal3 33604 4692 33604 4692 0 FrameData_O[13]
rlabel metal3 33420 4964 33420 4964 0 FrameData_O[14]
rlabel metal3 33604 5236 33604 5236 0 FrameData_O[15]
rlabel metal3 33880 5508 33880 5508 0 FrameData_O[16]
rlabel metal3 33604 5780 33604 5780 0 FrameData_O[17]
rlabel metal3 33420 6052 33420 6052 0 FrameData_O[18]
rlabel metal3 33604 6324 33604 6324 0 FrameData_O[19]
rlabel metal3 32914 1428 32914 1428 0 FrameData_O[1]
rlabel metal3 33880 6596 33880 6596 0 FrameData_O[20]
rlabel metal3 33604 6868 33604 6868 0 FrameData_O[21]
rlabel metal3 33604 7140 33604 7140 0 FrameData_O[22]
rlabel metal3 33420 7412 33420 7412 0 FrameData_O[23]
rlabel metal3 33972 7684 33972 7684 0 FrameData_O[24]
rlabel metal3 33604 7956 33604 7956 0 FrameData_O[25]
rlabel metal3 33420 8228 33420 8228 0 FrameData_O[26]
rlabel metal3 33098 8500 33098 8500 0 FrameData_O[27]
rlabel metal3 33949 8772 33949 8772 0 FrameData_O[28]
rlabel metal1 32798 8058 32798 8058 0 FrameData_O[29]
rlabel metal3 33144 1700 33144 1700 0 FrameData_O[2]
rlabel metal1 32568 7514 32568 7514 0 FrameData_O[30]
rlabel metal2 31786 8823 31786 8823 0 FrameData_O[31]
rlabel metal3 32730 1972 32730 1972 0 FrameData_O[3]
rlabel metal3 33880 2244 33880 2244 0 FrameData_O[4]
rlabel metal3 33604 2516 33604 2516 0 FrameData_O[5]
rlabel metal3 33420 2788 33420 2788 0 FrameData_O[6]
rlabel metal3 33604 3060 33604 3060 0 FrameData_O[7]
rlabel metal3 33880 3332 33880 3332 0 FrameData_O[8]
rlabel metal3 33604 3604 33604 3604 0 FrameData_O[9]
rlabel metal2 3082 55 3082 55 0 FrameStrobe[0]
rlabel metal2 18722 2248 18722 2248 0 FrameStrobe[10]
rlabel metal2 20286 1160 20286 1160 0 FrameStrobe[11]
rlabel metal2 21850 2843 21850 2843 0 FrameStrobe[12]
rlabel metal3 25760 5100 25760 5100 0 FrameStrobe[13]
rlabel metal1 26496 7378 26496 7378 0 FrameStrobe[14]
rlabel metal3 27830 7004 27830 7004 0 FrameStrobe[15]
rlabel metal2 28106 1347 28106 1347 0 FrameStrobe[16]
rlabel metal1 29946 7310 29946 7310 0 FrameStrobe[17]
rlabel metal1 31050 7378 31050 7378 0 FrameStrobe[18]
rlabel metal2 32798 3744 32798 3744 0 FrameStrobe[19]
rlabel metal1 7912 3434 7912 3434 0 FrameStrobe[1]
rlabel metal2 14306 3298 14306 3298 0 FrameStrobe[2]
rlabel metal1 13271 4590 13271 4590 0 FrameStrobe[3]
rlabel metal2 9338 735 9338 735 0 FrameStrobe[4]
rlabel metal2 10902 1058 10902 1058 0 FrameStrobe[5]
rlabel metal2 12466 1602 12466 1602 0 FrameStrobe[6]
rlabel metal2 14030 55 14030 55 0 FrameStrobe[7]
rlabel metal1 16468 3638 16468 3638 0 FrameStrobe[8]
rlabel metal2 17158 1007 17158 1007 0 FrameStrobe[9]
rlabel metal1 25300 8602 25300 8602 0 FrameStrobe_O[0]
rlabel metal1 27048 8058 27048 8058 0 FrameStrobe_O[10]
rlabel metal1 28198 8568 28198 8568 0 FrameStrobe_O[11]
rlabel metal1 27508 8058 27508 8058 0 FrameStrobe_O[12]
rlabel metal2 28566 8772 28566 8772 0 FrameStrobe_O[13]
rlabel metal1 27876 8058 27876 8058 0 FrameStrobe_O[14]
rlabel metal1 28428 8330 28428 8330 0 FrameStrobe_O[15]
rlabel metal1 28198 8058 28198 8058 0 FrameStrobe_O[16]
rlabel metal1 28520 8058 28520 8058 0 FrameStrobe_O[17]
rlabel metal1 28750 7718 28750 7718 0 FrameStrobe_O[18]
rlabel metal1 29164 8602 29164 8602 0 FrameStrobe_O[19]
rlabel metal1 25576 8330 25576 8330 0 FrameStrobe_O[1]
rlabel metal1 25852 8602 25852 8602 0 FrameStrobe_O[2]
rlabel metal1 26542 8568 26542 8568 0 FrameStrobe_O[3]
rlabel metal1 26036 8058 26036 8058 0 FrameStrobe_O[4]
rlabel metal1 26634 8330 26634 8330 0 FrameStrobe_O[5]
rlabel metal1 26450 8058 26450 8058 0 FrameStrobe_O[6]
rlabel metal1 27554 8364 27554 8364 0 FrameStrobe_O[7]
rlabel metal1 26726 8058 26726 8058 0 FrameStrobe_O[8]
rlabel metal1 27324 8602 27324 8602 0 FrameStrobe_O[9]
rlabel metal1 5336 8602 5336 8602 0 N1BEG[0]
rlabel metal1 5796 8058 5796 8058 0 N1BEG[1]
rlabel metal1 5704 8330 5704 8330 0 N1BEG[2]
rlabel metal1 6164 8058 6164 8058 0 N1BEG[3]
rlabel metal1 5750 8568 5750 8568 0 N2BEG[0]
rlabel metal1 6532 8058 6532 8058 0 N2BEG[1]
rlabel metal1 6440 8602 6440 8602 0 N2BEG[2]
rlabel metal1 6900 8058 6900 8058 0 N2BEG[3]
rlabel metal1 7268 7514 7268 7514 0 N2BEG[4]
rlabel metal1 7268 8058 7268 8058 0 N2BEG[5]
rlabel metal1 7176 8602 7176 8602 0 N2BEG[6]
rlabel metal1 7636 8058 7636 8058 0 N2BEG[7]
rlabel metal1 7130 8432 7130 8432 0 N2BEGb[0]
rlabel metal2 7866 8755 7866 8755 0 N2BEGb[1]
rlabel metal1 7544 8330 7544 8330 0 N2BEGb[2]
rlabel metal1 8372 8058 8372 8058 0 N2BEGb[3]
rlabel metal1 7958 8568 7958 8568 0 N2BEGb[4]
rlabel metal1 8740 8058 8740 8058 0 N2BEGb[5]
rlabel metal1 8602 8602 8602 8602 0 N2BEGb[6]
rlabel metal2 9430 8347 9430 8347 0 N2BEGb[7]
rlabel metal1 8648 8330 8648 8330 0 N4BEG[0]
rlabel metal1 10488 8602 10488 8602 0 N4BEG[10]
rlabel metal1 11270 8058 11270 8058 0 N4BEG[11]
rlabel metal1 11178 8330 11178 8330 0 N4BEG[12]
rlabel metal1 11638 8058 11638 8058 0 N4BEG[13]
rlabel metal1 11546 8602 11546 8602 0 N4BEG[14]
rlabel metal1 12052 8058 12052 8058 0 N4BEG[15]
rlabel metal1 9430 8058 9430 8058 0 N4BEG[1]
rlabel metal1 9798 7514 9798 7514 0 N4BEG[2]
rlabel metal1 9798 8058 9798 8058 0 N4BEG[3]
rlabel metal1 9706 8602 9706 8602 0 N4BEG[4]
rlabel metal1 10166 8058 10166 8058 0 N4BEG[5]
rlabel metal1 10074 8330 10074 8330 0 N4BEG[6]
rlabel metal1 10534 8058 10534 8058 0 N4BEG[7]
rlabel metal2 10074 8381 10074 8381 0 N4BEG[8]
rlabel metal1 10902 8058 10902 8058 0 N4BEG[9]
rlabel metal2 12282 9584 12282 9584 0 NN4BEG[0]
rlabel metal1 13938 8602 13938 8602 0 NN4BEG[10]
rlabel metal1 14398 8058 14398 8058 0 NN4BEG[11]
rlabel metal2 14490 9856 14490 9856 0 NN4BEG[12]
rlabel metal1 14766 8602 14766 8602 0 NN4BEG[13]
rlabel metal1 15456 8262 15456 8262 0 NN4BEG[14]
rlabel metal1 15088 8602 15088 8602 0 NN4BEG[15]
rlabel metal1 12558 8058 12558 8058 0 NN4BEG[1]
rlabel metal1 12282 8262 12282 8262 0 NN4BEG[2]
rlabel metal1 12926 8058 12926 8058 0 NN4BEG[3]
rlabel metal2 13018 9992 13018 9992 0 NN4BEG[4]
rlabel metal1 13294 8058 13294 8058 0 NN4BEG[5]
rlabel metal1 13018 8602 13018 8602 0 NN4BEG[6]
rlabel metal1 13662 8058 13662 8058 0 NN4BEG[7]
rlabel metal1 13156 8330 13156 8330 0 NN4BEG[8]
rlabel metal1 13616 8330 13616 8330 0 NN4BEG[9]
rlabel metal2 15410 10621 15410 10621 0 S1END[0]
rlabel metal2 15594 10553 15594 10553 0 S1END[1]
rlabel metal2 2530 7616 2530 7616 0 S1END[2]
rlabel metal2 2162 7684 2162 7684 0 S1END[3]
rlabel metal2 17618 10009 17618 10009 0 S2END[0]
rlabel metal2 17802 10808 17802 10808 0 S2END[1]
rlabel metal2 17986 11046 17986 11046 0 S2END[2]
rlabel metal2 18170 11097 18170 11097 0 S2END[3]
rlabel via2 18354 11097 18354 11097 0 S2END[4]
rlabel metal2 18538 10689 18538 10689 0 S2END[5]
rlabel metal2 18722 10978 18722 10978 0 S2END[6]
rlabel metal2 18906 8717 18906 8717 0 S2END[7]
rlabel metal2 16146 10876 16146 10876 0 S2MID[0]
rlabel metal2 16330 10485 16330 10485 0 S2MID[1]
rlabel metal2 16514 8462 16514 8462 0 S2MID[2]
rlabel metal2 16698 10621 16698 10621 0 S2MID[3]
rlabel metal2 16882 10009 16882 10009 0 S2MID[4]
rlabel metal2 17066 8972 17066 8972 0 S2MID[5]
rlabel metal2 17250 8734 17250 8734 0 S2MID[6]
rlabel metal2 17434 8445 17434 8445 0 S2MID[7]
rlabel metal2 19090 9006 19090 9006 0 S4END[0]
rlabel metal2 20930 10145 20930 10145 0 S4END[10]
rlabel metal2 21114 10128 21114 10128 0 S4END[11]
rlabel metal2 21298 10077 21298 10077 0 S4END[12]
rlabel metal2 21482 7289 21482 7289 0 S4END[13]
rlabel metal2 21666 7085 21666 7085 0 S4END[14]
rlabel metal2 21850 10009 21850 10009 0 S4END[15]
rlabel metal2 19274 10434 19274 10434 0 S4END[1]
rlabel metal2 19458 8598 19458 8598 0 S4END[2]
rlabel metal2 19642 10349 19642 10349 0 S4END[3]
rlabel metal2 19826 10638 19826 10638 0 S4END[4]
rlabel metal2 20010 9686 20010 9686 0 S4END[5]
rlabel metal2 20194 10536 20194 10536 0 S4END[6]
rlabel metal2 20378 9584 20378 9584 0 S4END[7]
rlabel metal2 20562 7816 20562 7816 0 S4END[8]
rlabel metal2 20746 10366 20746 10366 0 S4END[9]
rlabel metal2 22034 10145 22034 10145 0 SS4END[0]
rlabel metal2 23874 8734 23874 8734 0 SS4END[10]
rlabel metal2 24058 8666 24058 8666 0 SS4END[11]
rlabel metal2 24242 8768 24242 8768 0 SS4END[12]
rlabel metal1 21666 6324 21666 6324 0 SS4END[13]
rlabel metal2 22034 7599 22034 7599 0 SS4END[14]
rlabel metal2 24794 10417 24794 10417 0 SS4END[15]
rlabel metal2 22218 9414 22218 9414 0 SS4END[1]
rlabel metal2 22402 8989 22402 8989 0 SS4END[2]
rlabel metal2 22586 9941 22586 9941 0 SS4END[3]
rlabel metal2 22770 10026 22770 10026 0 SS4END[4]
rlabel metal2 22954 9720 22954 9720 0 SS4END[5]
rlabel metal2 23138 9006 23138 9006 0 SS4END[6]
rlabel metal2 23322 8972 23322 8972 0 SS4END[7]
rlabel metal2 23506 8938 23506 8938 0 SS4END[8]
rlabel metal2 23690 8700 23690 8700 0 SS4END[9]
rlabel metal2 1518 1772 1518 1772 0 UserCLK
rlabel metal2 24978 9856 24978 9856 0 UserCLKo
rlabel metal1 31050 2414 31050 2414 0 net1
rlabel metal2 32338 6086 32338 6086 0 net10
rlabel metal1 17802 8024 17802 8024 0 net100
rlabel metal2 18078 7412 18078 7412 0 net101
rlabel metal2 20378 7208 20378 7208 0 net102
rlabel metal2 13478 8976 13478 8976 0 net103
rlabel metal2 13846 8840 13846 8840 0 net104
rlabel metal2 10534 6103 10534 6103 0 net105
rlabel metal1 15640 8330 15640 8330 0 net106
rlabel via2 17802 3621 17802 3621 0 net11
rlabel metal2 31326 2516 31326 2516 0 net12
rlabel metal1 18446 3706 18446 3706 0 net13
rlabel metal2 32430 6256 32430 6256 0 net14
rlabel metal1 17664 7514 17664 7514 0 net15
rlabel metal2 32338 7412 32338 7412 0 net16
rlabel metal1 20194 7276 20194 7276 0 net17
rlabel metal1 21206 7514 21206 7514 0 net18
rlabel metal2 19826 8398 19826 8398 0 net19
rlabel metal2 18078 4862 18078 4862 0 net2
rlabel metal2 19550 8466 19550 8466 0 net20
rlabel metal1 17480 7242 17480 7242 0 net21
rlabel metal1 21298 7412 21298 7412 0 net22
rlabel metal2 14490 4726 14490 4726 0 net23
rlabel metal1 21390 7480 21390 7480 0 net24
rlabel metal2 18538 7718 18538 7718 0 net25
rlabel metal2 13754 4420 13754 4420 0 net26
rlabel metal1 32062 2414 32062 2414 0 net27
rlabel metal1 31142 2516 31142 2516 0 net28
rlabel metal2 19826 5355 19826 5355 0 net29
rlabel metal2 18354 4896 18354 4896 0 net3
rlabel metal2 18538 4080 18538 4080 0 net30
rlabel metal2 14398 4488 14398 4488 0 net31
rlabel metal2 32430 3978 32430 3978 0 net32
rlabel metal2 21574 5236 21574 5236 0 net33
rlabel metal1 28244 4794 28244 4794 0 net34
rlabel metal1 28888 6630 28888 6630 0 net35
rlabel metal1 28198 7242 28198 7242 0 net36
rlabel metal1 28658 7514 28658 7514 0 net37
rlabel metal2 27830 7684 27830 7684 0 net38
rlabel metal2 28934 7990 28934 7990 0 net39
rlabel metal2 16606 5100 16606 5100 0 net4
rlabel metal1 29164 7514 29164 7514 0 net40
rlabel metal1 29440 7242 29440 7242 0 net41
rlabel metal2 30682 7684 30682 7684 0 net42
rlabel metal1 29808 7514 29808 7514 0 net43
rlabel metal2 17250 3808 17250 3808 0 net44
rlabel metal1 14812 3706 14812 3706 0 net45
rlabel metal1 15732 4454 15732 4454 0 net46
rlabel metal2 21114 3808 21114 3808 0 net47
rlabel metal1 21919 3366 21919 3366 0 net48
rlabel metal1 24058 3706 24058 3706 0 net49
rlabel metal2 16422 5389 16422 5389 0 net5
rlabel metal1 27324 3706 27324 3706 0 net50
rlabel metal1 28658 3706 28658 3706 0 net51
rlabel metal1 28842 3638 28842 3638 0 net52
rlabel metal1 2553 7242 2553 7242 0 net53
rlabel metal2 2806 7684 2806 7684 0 net54
rlabel metal1 4140 7242 4140 7242 0 net55
rlabel metal1 4646 7514 4646 7514 0 net56
rlabel metal1 5152 6426 5152 6426 0 net57
rlabel metal1 5520 6086 5520 6086 0 net58
rlabel metal1 5382 6154 5382 6154 0 net59
rlabel metal2 15042 4964 15042 4964 0 net6
rlabel metal1 4278 6188 4278 6188 0 net60
rlabel metal2 4002 7174 4002 7174 0 net61
rlabel metal1 5520 6630 5520 6630 0 net62
rlabel metal1 3910 6630 3910 6630 0 net63
rlabel metal1 3358 6664 3358 6664 0 net64
rlabel metal2 7590 7191 7590 7191 0 net65
rlabel metal2 8418 7106 8418 7106 0 net66
rlabel metal1 7958 6426 7958 6426 0 net67
rlabel metal2 7498 7174 7498 7174 0 net68
rlabel metal2 7222 7650 7222 7650 0 net69
rlabel metal2 19734 5508 19734 5508 0 net7
rlabel metal1 8004 5882 8004 5882 0 net70
rlabel metal1 6624 6426 6624 6426 0 net71
rlabel metal1 8326 6630 8326 6630 0 net72
rlabel metal2 12650 5899 12650 5899 0 net73
rlabel metal1 12788 7514 12788 7514 0 net74
rlabel metal1 11960 7514 11960 7514 0 net75
rlabel metal1 11500 7242 11500 7242 0 net76
rlabel metal1 11914 6970 11914 6970 0 net77
rlabel metal1 12006 6630 12006 6630 0 net78
rlabel metal1 11592 7514 11592 7514 0 net79
rlabel metal2 27462 4658 27462 4658 0 net8
rlabel metal1 12144 3910 12144 3910 0 net80
rlabel metal2 12374 5712 12374 5712 0 net81
rlabel metal1 12098 4012 12098 4012 0 net82
rlabel metal1 10810 3910 10810 3910 0 net83
rlabel metal1 11592 3706 11592 3706 0 net84
rlabel metal1 10948 3978 10948 3978 0 net85
rlabel metal1 11730 4794 11730 4794 0 net86
rlabel metal1 12190 7514 12190 7514 0 net87
rlabel metal2 12558 7616 12558 7616 0 net88
rlabel metal1 21850 6188 21850 6188 0 net89
rlabel metal2 15778 3094 15778 3094 0 net9
rlabel metal2 14582 8636 14582 8636 0 net90
rlabel metal2 14674 6800 14674 6800 0 net91
rlabel metal1 18354 8568 18354 8568 0 net92
rlabel metal2 14950 7582 14950 7582 0 net93
rlabel metal1 26496 6630 26496 6630 0 net94
rlabel metal2 15686 9010 15686 9010 0 net95
rlabel metal1 21712 6086 21712 6086 0 net96
rlabel metal1 21206 6086 21206 6086 0 net97
rlabel metal2 17618 6528 17618 6528 0 net98
rlabel metal1 21942 6256 21942 6256 0 net99
<< properties >>
string FIXED_BBOX 0 0 34408 11152
<< end >>
