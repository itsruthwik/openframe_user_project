VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DSP
  CLASS BLOCK ;
  FOREIGN DSP ;
  ORIGIN 0.000 0.000 ;
  SIZE 199.640 BY 519.520 ;
  PIN Tile_X0Y0_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 367.240 199.640 367.840 ;
    END
  END Tile_X0Y0_E1BEG[0]
  PIN Tile_X0Y0_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 368.600 199.640 369.200 ;
    END
  END Tile_X0Y0_E1BEG[1]
  PIN Tile_X0Y0_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 369.960 199.640 370.560 ;
    END
  END Tile_X0Y0_E1BEG[2]
  PIN Tile_X0Y0_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 371.320 199.640 371.920 ;
    END
  END Tile_X0Y0_E1BEG[3]
  PIN Tile_X0Y0_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 0.600 367.840 ;
    END
  END Tile_X0Y0_E1END[0]
  PIN Tile_X0Y0_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 0.600 369.200 ;
    END
  END Tile_X0Y0_E1END[1]
  PIN Tile_X0Y0_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 0.600 370.560 ;
    END
  END Tile_X0Y0_E1END[2]
  PIN Tile_X0Y0_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 0.600 371.920 ;
    END
  END Tile_X0Y0_E1END[3]
  PIN Tile_X0Y0_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 372.680 199.640 373.280 ;
    END
  END Tile_X0Y0_E2BEG[0]
  PIN Tile_X0Y0_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 374.040 199.640 374.640 ;
    END
  END Tile_X0Y0_E2BEG[1]
  PIN Tile_X0Y0_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 375.400 199.640 376.000 ;
    END
  END Tile_X0Y0_E2BEG[2]
  PIN Tile_X0Y0_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 376.760 199.640 377.360 ;
    END
  END Tile_X0Y0_E2BEG[3]
  PIN Tile_X0Y0_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 378.120 199.640 378.720 ;
    END
  END Tile_X0Y0_E2BEG[4]
  PIN Tile_X0Y0_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 379.480 199.640 380.080 ;
    END
  END Tile_X0Y0_E2BEG[5]
  PIN Tile_X0Y0_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 380.840 199.640 381.440 ;
    END
  END Tile_X0Y0_E2BEG[6]
  PIN Tile_X0Y0_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 382.200 199.640 382.800 ;
    END
  END Tile_X0Y0_E2BEG[7]
  PIN Tile_X0Y0_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 383.560 199.640 384.160 ;
    END
  END Tile_X0Y0_E2BEGb[0]
  PIN Tile_X0Y0_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 384.920 199.640 385.520 ;
    END
  END Tile_X0Y0_E2BEGb[1]
  PIN Tile_X0Y0_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 386.280 199.640 386.880 ;
    END
  END Tile_X0Y0_E2BEGb[2]
  PIN Tile_X0Y0_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 387.640 199.640 388.240 ;
    END
  END Tile_X0Y0_E2BEGb[3]
  PIN Tile_X0Y0_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 389.000 199.640 389.600 ;
    END
  END Tile_X0Y0_E2BEGb[4]
  PIN Tile_X0Y0_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 390.360 199.640 390.960 ;
    END
  END Tile_X0Y0_E2BEGb[5]
  PIN Tile_X0Y0_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 391.720 199.640 392.320 ;
    END
  END Tile_X0Y0_E2BEGb[6]
  PIN Tile_X0Y0_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 393.080 199.640 393.680 ;
    END
  END Tile_X0Y0_E2BEGb[7]
  PIN Tile_X0Y0_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 0.600 384.160 ;
    END
  END Tile_X0Y0_E2END[0]
  PIN Tile_X0Y0_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 0.600 385.520 ;
    END
  END Tile_X0Y0_E2END[1]
  PIN Tile_X0Y0_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 0.600 386.880 ;
    END
  END Tile_X0Y0_E2END[2]
  PIN Tile_X0Y0_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 0.600 388.240 ;
    END
  END Tile_X0Y0_E2END[3]
  PIN Tile_X0Y0_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 0.600 389.600 ;
    END
  END Tile_X0Y0_E2END[4]
  PIN Tile_X0Y0_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 0.600 390.960 ;
    END
  END Tile_X0Y0_E2END[5]
  PIN Tile_X0Y0_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 0.600 392.320 ;
    END
  END Tile_X0Y0_E2END[6]
  PIN Tile_X0Y0_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 0.600 393.680 ;
    END
  END Tile_X0Y0_E2END[7]
  PIN Tile_X0Y0_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 0.600 373.280 ;
    END
  END Tile_X0Y0_E2MID[0]
  PIN Tile_X0Y0_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 0.600 374.640 ;
    END
  END Tile_X0Y0_E2MID[1]
  PIN Tile_X0Y0_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 0.600 376.000 ;
    END
  END Tile_X0Y0_E2MID[2]
  PIN Tile_X0Y0_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 0.600 377.360 ;
    END
  END Tile_X0Y0_E2MID[3]
  PIN Tile_X0Y0_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 0.600 378.720 ;
    END
  END Tile_X0Y0_E2MID[4]
  PIN Tile_X0Y0_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 0.600 380.080 ;
    END
  END Tile_X0Y0_E2MID[5]
  PIN Tile_X0Y0_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 0.600 381.440 ;
    END
  END Tile_X0Y0_E2MID[6]
  PIN Tile_X0Y0_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 0.600 382.800 ;
    END
  END Tile_X0Y0_E2MID[7]
  PIN Tile_X0Y0_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 416.200 199.640 416.800 ;
    END
  END Tile_X0Y0_E6BEG[0]
  PIN Tile_X0Y0_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 429.800 199.640 430.400 ;
    END
  END Tile_X0Y0_E6BEG[10]
  PIN Tile_X0Y0_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 431.160 199.640 431.760 ;
    END
  END Tile_X0Y0_E6BEG[11]
  PIN Tile_X0Y0_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 417.560 199.640 418.160 ;
    END
  END Tile_X0Y0_E6BEG[1]
  PIN Tile_X0Y0_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 418.920 199.640 419.520 ;
    END
  END Tile_X0Y0_E6BEG[2]
  PIN Tile_X0Y0_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 420.280 199.640 420.880 ;
    END
  END Tile_X0Y0_E6BEG[3]
  PIN Tile_X0Y0_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 421.640 199.640 422.240 ;
    END
  END Tile_X0Y0_E6BEG[4]
  PIN Tile_X0Y0_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 423.000 199.640 423.600 ;
    END
  END Tile_X0Y0_E6BEG[5]
  PIN Tile_X0Y0_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 424.360 199.640 424.960 ;
    END
  END Tile_X0Y0_E6BEG[6]
  PIN Tile_X0Y0_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 425.720 199.640 426.320 ;
    END
  END Tile_X0Y0_E6BEG[7]
  PIN Tile_X0Y0_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 427.080 199.640 427.680 ;
    END
  END Tile_X0Y0_E6BEG[8]
  PIN Tile_X0Y0_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 428.440 199.640 429.040 ;
    END
  END Tile_X0Y0_E6BEG[9]
  PIN Tile_X0Y0_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 0.600 416.800 ;
    END
  END Tile_X0Y0_E6END[0]
  PIN Tile_X0Y0_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 0.600 430.400 ;
    END
  END Tile_X0Y0_E6END[10]
  PIN Tile_X0Y0_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 0.600 431.760 ;
    END
  END Tile_X0Y0_E6END[11]
  PIN Tile_X0Y0_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 0.600 418.160 ;
    END
  END Tile_X0Y0_E6END[1]
  PIN Tile_X0Y0_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 0.600 419.520 ;
    END
  END Tile_X0Y0_E6END[2]
  PIN Tile_X0Y0_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 0.600 420.880 ;
    END
  END Tile_X0Y0_E6END[3]
  PIN Tile_X0Y0_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 0.600 422.240 ;
    END
  END Tile_X0Y0_E6END[4]
  PIN Tile_X0Y0_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 0.600 423.600 ;
    END
  END Tile_X0Y0_E6END[5]
  PIN Tile_X0Y0_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 0.600 424.960 ;
    END
  END Tile_X0Y0_E6END[6]
  PIN Tile_X0Y0_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 0.600 426.320 ;
    END
  END Tile_X0Y0_E6END[7]
  PIN Tile_X0Y0_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 0.600 427.680 ;
    END
  END Tile_X0Y0_E6END[8]
  PIN Tile_X0Y0_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 0.600 429.040 ;
    END
  END Tile_X0Y0_E6END[9]
  PIN Tile_X0Y0_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 394.440 199.640 395.040 ;
    END
  END Tile_X0Y0_EE4BEG[0]
  PIN Tile_X0Y0_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 408.040 199.640 408.640 ;
    END
  END Tile_X0Y0_EE4BEG[10]
  PIN Tile_X0Y0_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 409.400 199.640 410.000 ;
    END
  END Tile_X0Y0_EE4BEG[11]
  PIN Tile_X0Y0_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 410.760 199.640 411.360 ;
    END
  END Tile_X0Y0_EE4BEG[12]
  PIN Tile_X0Y0_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 412.120 199.640 412.720 ;
    END
  END Tile_X0Y0_EE4BEG[13]
  PIN Tile_X0Y0_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 413.480 199.640 414.080 ;
    END
  END Tile_X0Y0_EE4BEG[14]
  PIN Tile_X0Y0_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 414.840 199.640 415.440 ;
    END
  END Tile_X0Y0_EE4BEG[15]
  PIN Tile_X0Y0_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 395.800 199.640 396.400 ;
    END
  END Tile_X0Y0_EE4BEG[1]
  PIN Tile_X0Y0_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 397.160 199.640 397.760 ;
    END
  END Tile_X0Y0_EE4BEG[2]
  PIN Tile_X0Y0_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 398.520 199.640 399.120 ;
    END
  END Tile_X0Y0_EE4BEG[3]
  PIN Tile_X0Y0_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 399.880 199.640 400.480 ;
    END
  END Tile_X0Y0_EE4BEG[4]
  PIN Tile_X0Y0_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 401.240 199.640 401.840 ;
    END
  END Tile_X0Y0_EE4BEG[5]
  PIN Tile_X0Y0_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 402.600 199.640 403.200 ;
    END
  END Tile_X0Y0_EE4BEG[6]
  PIN Tile_X0Y0_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 403.960 199.640 404.560 ;
    END
  END Tile_X0Y0_EE4BEG[7]
  PIN Tile_X0Y0_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 405.320 199.640 405.920 ;
    END
  END Tile_X0Y0_EE4BEG[8]
  PIN Tile_X0Y0_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 406.680 199.640 407.280 ;
    END
  END Tile_X0Y0_EE4BEG[9]
  PIN Tile_X0Y0_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 0.600 395.040 ;
    END
  END Tile_X0Y0_EE4END[0]
  PIN Tile_X0Y0_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 0.600 408.640 ;
    END
  END Tile_X0Y0_EE4END[10]
  PIN Tile_X0Y0_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 0.600 410.000 ;
    END
  END Tile_X0Y0_EE4END[11]
  PIN Tile_X0Y0_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 0.600 411.360 ;
    END
  END Tile_X0Y0_EE4END[12]
  PIN Tile_X0Y0_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 0.600 412.720 ;
    END
  END Tile_X0Y0_EE4END[13]
  PIN Tile_X0Y0_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 0.600 414.080 ;
    END
  END Tile_X0Y0_EE4END[14]
  PIN Tile_X0Y0_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 0.600 415.440 ;
    END
  END Tile_X0Y0_EE4END[15]
  PIN Tile_X0Y0_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 0.600 396.400 ;
    END
  END Tile_X0Y0_EE4END[1]
  PIN Tile_X0Y0_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 0.600 397.760 ;
    END
  END Tile_X0Y0_EE4END[2]
  PIN Tile_X0Y0_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 0.600 399.120 ;
    END
  END Tile_X0Y0_EE4END[3]
  PIN Tile_X0Y0_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 0.600 400.480 ;
    END
  END Tile_X0Y0_EE4END[4]
  PIN Tile_X0Y0_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 0.600 401.840 ;
    END
  END Tile_X0Y0_EE4END[5]
  PIN Tile_X0Y0_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 0.600 403.200 ;
    END
  END Tile_X0Y0_EE4END[6]
  PIN Tile_X0Y0_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 0.600 404.560 ;
    END
  END Tile_X0Y0_EE4END[7]
  PIN Tile_X0Y0_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 0.600 405.920 ;
    END
  END Tile_X0Y0_EE4END[8]
  PIN Tile_X0Y0_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 0.600 407.280 ;
    END
  END Tile_X0Y0_EE4END[9]
  PIN Tile_X0Y0_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 0.600 433.120 ;
    END
  END Tile_X0Y0_FrameData[0]
  PIN Tile_X0Y0_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 0.600 446.720 ;
    END
  END Tile_X0Y0_FrameData[10]
  PIN Tile_X0Y0_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 0.600 448.080 ;
    END
  END Tile_X0Y0_FrameData[11]
  PIN Tile_X0Y0_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 0.600 449.440 ;
    END
  END Tile_X0Y0_FrameData[12]
  PIN Tile_X0Y0_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 0.600 450.800 ;
    END
  END Tile_X0Y0_FrameData[13]
  PIN Tile_X0Y0_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 0.600 452.160 ;
    END
  END Tile_X0Y0_FrameData[14]
  PIN Tile_X0Y0_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 0.600 453.520 ;
    END
  END Tile_X0Y0_FrameData[15]
  PIN Tile_X0Y0_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 0.600 454.880 ;
    END
  END Tile_X0Y0_FrameData[16]
  PIN Tile_X0Y0_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 0.600 456.240 ;
    END
  END Tile_X0Y0_FrameData[17]
  PIN Tile_X0Y0_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 0.600 457.600 ;
    END
  END Tile_X0Y0_FrameData[18]
  PIN Tile_X0Y0_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 0.600 458.960 ;
    END
  END Tile_X0Y0_FrameData[19]
  PIN Tile_X0Y0_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 0.600 434.480 ;
    END
  END Tile_X0Y0_FrameData[1]
  PIN Tile_X0Y0_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 0.600 460.320 ;
    END
  END Tile_X0Y0_FrameData[20]
  PIN Tile_X0Y0_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 0.600 461.680 ;
    END
  END Tile_X0Y0_FrameData[21]
  PIN Tile_X0Y0_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 0.600 463.040 ;
    END
  END Tile_X0Y0_FrameData[22]
  PIN Tile_X0Y0_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 0.600 464.400 ;
    END
  END Tile_X0Y0_FrameData[23]
  PIN Tile_X0Y0_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 0.600 465.760 ;
    END
  END Tile_X0Y0_FrameData[24]
  PIN Tile_X0Y0_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 0.600 467.120 ;
    END
  END Tile_X0Y0_FrameData[25]
  PIN Tile_X0Y0_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 0.600 468.480 ;
    END
  END Tile_X0Y0_FrameData[26]
  PIN Tile_X0Y0_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 0.600 469.840 ;
    END
  END Tile_X0Y0_FrameData[27]
  PIN Tile_X0Y0_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 0.600 471.200 ;
    END
  END Tile_X0Y0_FrameData[28]
  PIN Tile_X0Y0_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 0.600 472.560 ;
    END
  END Tile_X0Y0_FrameData[29]
  PIN Tile_X0Y0_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 0.600 435.840 ;
    END
  END Tile_X0Y0_FrameData[2]
  PIN Tile_X0Y0_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 0.600 473.920 ;
    END
  END Tile_X0Y0_FrameData[30]
  PIN Tile_X0Y0_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 0.600 475.280 ;
    END
  END Tile_X0Y0_FrameData[31]
  PIN Tile_X0Y0_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 0.600 437.200 ;
    END
  END Tile_X0Y0_FrameData[3]
  PIN Tile_X0Y0_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 0.600 438.560 ;
    END
  END Tile_X0Y0_FrameData[4]
  PIN Tile_X0Y0_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 0.600 439.920 ;
    END
  END Tile_X0Y0_FrameData[5]
  PIN Tile_X0Y0_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 0.600 441.280 ;
    END
  END Tile_X0Y0_FrameData[6]
  PIN Tile_X0Y0_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 0.600 442.640 ;
    END
  END Tile_X0Y0_FrameData[7]
  PIN Tile_X0Y0_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 0.600 444.000 ;
    END
  END Tile_X0Y0_FrameData[8]
  PIN Tile_X0Y0_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 0.600 445.360 ;
    END
  END Tile_X0Y0_FrameData[9]
  PIN Tile_X0Y0_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 432.520 199.640 433.120 ;
    END
  END Tile_X0Y0_FrameData_O[0]
  PIN Tile_X0Y0_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 446.120 199.640 446.720 ;
    END
  END Tile_X0Y0_FrameData_O[10]
  PIN Tile_X0Y0_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 447.480 199.640 448.080 ;
    END
  END Tile_X0Y0_FrameData_O[11]
  PIN Tile_X0Y0_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 448.840 199.640 449.440 ;
    END
  END Tile_X0Y0_FrameData_O[12]
  PIN Tile_X0Y0_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 450.200 199.640 450.800 ;
    END
  END Tile_X0Y0_FrameData_O[13]
  PIN Tile_X0Y0_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 451.560 199.640 452.160 ;
    END
  END Tile_X0Y0_FrameData_O[14]
  PIN Tile_X0Y0_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 452.920 199.640 453.520 ;
    END
  END Tile_X0Y0_FrameData_O[15]
  PIN Tile_X0Y0_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 454.280 199.640 454.880 ;
    END
  END Tile_X0Y0_FrameData_O[16]
  PIN Tile_X0Y0_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 455.640 199.640 456.240 ;
    END
  END Tile_X0Y0_FrameData_O[17]
  PIN Tile_X0Y0_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 457.000 199.640 457.600 ;
    END
  END Tile_X0Y0_FrameData_O[18]
  PIN Tile_X0Y0_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 458.360 199.640 458.960 ;
    END
  END Tile_X0Y0_FrameData_O[19]
  PIN Tile_X0Y0_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 433.880 199.640 434.480 ;
    END
  END Tile_X0Y0_FrameData_O[1]
  PIN Tile_X0Y0_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 459.720 199.640 460.320 ;
    END
  END Tile_X0Y0_FrameData_O[20]
  PIN Tile_X0Y0_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 461.080 199.640 461.680 ;
    END
  END Tile_X0Y0_FrameData_O[21]
  PIN Tile_X0Y0_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 462.440 199.640 463.040 ;
    END
  END Tile_X0Y0_FrameData_O[22]
  PIN Tile_X0Y0_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 463.800 199.640 464.400 ;
    END
  END Tile_X0Y0_FrameData_O[23]
  PIN Tile_X0Y0_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 465.160 199.640 465.760 ;
    END
  END Tile_X0Y0_FrameData_O[24]
  PIN Tile_X0Y0_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 466.520 199.640 467.120 ;
    END
  END Tile_X0Y0_FrameData_O[25]
  PIN Tile_X0Y0_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 467.880 199.640 468.480 ;
    END
  END Tile_X0Y0_FrameData_O[26]
  PIN Tile_X0Y0_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 469.240 199.640 469.840 ;
    END
  END Tile_X0Y0_FrameData_O[27]
  PIN Tile_X0Y0_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 470.600 199.640 471.200 ;
    END
  END Tile_X0Y0_FrameData_O[28]
  PIN Tile_X0Y0_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 471.960 199.640 472.560 ;
    END
  END Tile_X0Y0_FrameData_O[29]
  PIN Tile_X0Y0_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 435.240 199.640 435.840 ;
    END
  END Tile_X0Y0_FrameData_O[2]
  PIN Tile_X0Y0_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 473.320 199.640 473.920 ;
    END
  END Tile_X0Y0_FrameData_O[30]
  PIN Tile_X0Y0_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 474.680 199.640 475.280 ;
    END
  END Tile_X0Y0_FrameData_O[31]
  PIN Tile_X0Y0_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 436.600 199.640 437.200 ;
    END
  END Tile_X0Y0_FrameData_O[3]
  PIN Tile_X0Y0_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 437.960 199.640 438.560 ;
    END
  END Tile_X0Y0_FrameData_O[4]
  PIN Tile_X0Y0_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 439.320 199.640 439.920 ;
    END
  END Tile_X0Y0_FrameData_O[5]
  PIN Tile_X0Y0_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 440.680 199.640 441.280 ;
    END
  END Tile_X0Y0_FrameData_O[6]
  PIN Tile_X0Y0_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 442.040 199.640 442.640 ;
    END
  END Tile_X0Y0_FrameData_O[7]
  PIN Tile_X0Y0_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 443.400 199.640 444.000 ;
    END
  END Tile_X0Y0_FrameData_O[8]
  PIN Tile_X0Y0_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 444.760 199.640 445.360 ;
    END
  END Tile_X0Y0_FrameData_O[9]
  PIN Tile_X0Y0_FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 158.790 519.240 159.070 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[0]
  PIN Tile_X0Y0_FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 172.590 519.240 172.870 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[10]
  PIN Tile_X0Y0_FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 519.240 174.250 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[11]
  PIN Tile_X0Y0_FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 175.350 519.240 175.630 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[12]
  PIN Tile_X0Y0_FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 176.730 519.240 177.010 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[13]
  PIN Tile_X0Y0_FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 178.110 519.240 178.390 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[14]
  PIN Tile_X0Y0_FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 179.490 519.240 179.770 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[15]
  PIN Tile_X0Y0_FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 180.870 519.240 181.150 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[16]
  PIN Tile_X0Y0_FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 182.250 519.240 182.530 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[17]
  PIN Tile_X0Y0_FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 519.240 183.910 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[18]
  PIN Tile_X0Y0_FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 185.010 519.240 185.290 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[19]
  PIN Tile_X0Y0_FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 160.170 519.240 160.450 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[1]
  PIN Tile_X0Y0_FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 161.550 519.240 161.830 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[2]
  PIN Tile_X0Y0_FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.930 519.240 163.210 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[3]
  PIN Tile_X0Y0_FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 519.240 164.590 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[4]
  PIN Tile_X0Y0_FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 165.690 519.240 165.970 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[5]
  PIN Tile_X0Y0_FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 167.070 519.240 167.350 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[6]
  PIN Tile_X0Y0_FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 168.450 519.240 168.730 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[7]
  PIN Tile_X0Y0_FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 169.830 519.240 170.110 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[8]
  PIN Tile_X0Y0_FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 171.210 519.240 171.490 519.520 ;
    END
  END Tile_X0Y0_FrameStrobe_O[9]
  PIN Tile_X0Y0_N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 13.890 519.240 14.170 519.520 ;
    END
  END Tile_X0Y0_N1BEG[0]
  PIN Tile_X0Y0_N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 15.270 519.240 15.550 519.520 ;
    END
  END Tile_X0Y0_N1BEG[1]
  PIN Tile_X0Y0_N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 16.650 519.240 16.930 519.520 ;
    END
  END Tile_X0Y0_N1BEG[2]
  PIN Tile_X0Y0_N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 18.030 519.240 18.310 519.520 ;
    END
  END Tile_X0Y0_N1BEG[3]
  PIN Tile_X0Y0_N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 519.240 19.690 519.520 ;
    END
  END Tile_X0Y0_N2BEG[0]
  PIN Tile_X0Y0_N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 20.790 519.240 21.070 519.520 ;
    END
  END Tile_X0Y0_N2BEG[1]
  PIN Tile_X0Y0_N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.170 519.240 22.450 519.520 ;
    END
  END Tile_X0Y0_N2BEG[2]
  PIN Tile_X0Y0_N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 23.550 519.240 23.830 519.520 ;
    END
  END Tile_X0Y0_N2BEG[3]
  PIN Tile_X0Y0_N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 24.930 519.240 25.210 519.520 ;
    END
  END Tile_X0Y0_N2BEG[4]
  PIN Tile_X0Y0_N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 26.310 519.240 26.590 519.520 ;
    END
  END Tile_X0Y0_N2BEG[5]
  PIN Tile_X0Y0_N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 27.690 519.240 27.970 519.520 ;
    END
  END Tile_X0Y0_N2BEG[6]
  PIN Tile_X0Y0_N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 519.240 29.350 519.520 ;
    END
  END Tile_X0Y0_N2BEG[7]
  PIN Tile_X0Y0_N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 30.450 519.240 30.730 519.520 ;
    END
  END Tile_X0Y0_N2BEGb[0]
  PIN Tile_X0Y0_N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 31.830 519.240 32.110 519.520 ;
    END
  END Tile_X0Y0_N2BEGb[1]
  PIN Tile_X0Y0_N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 33.210 519.240 33.490 519.520 ;
    END
  END Tile_X0Y0_N2BEGb[2]
  PIN Tile_X0Y0_N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 34.590 519.240 34.870 519.520 ;
    END
  END Tile_X0Y0_N2BEGb[3]
  PIN Tile_X0Y0_N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 35.970 519.240 36.250 519.520 ;
    END
  END Tile_X0Y0_N2BEGb[4]
  PIN Tile_X0Y0_N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 37.350 519.240 37.630 519.520 ;
    END
  END Tile_X0Y0_N2BEGb[5]
  PIN Tile_X0Y0_N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 519.240 39.010 519.520 ;
    END
  END Tile_X0Y0_N2BEGb[6]
  PIN Tile_X0Y0_N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 40.110 519.240 40.390 519.520 ;
    END
  END Tile_X0Y0_N2BEGb[7]
  PIN Tile_X0Y0_N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.490 519.240 41.770 519.520 ;
    END
  END Tile_X0Y0_N4BEG[0]
  PIN Tile_X0Y0_N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 55.290 519.240 55.570 519.520 ;
    END
  END Tile_X0Y0_N4BEG[10]
  PIN Tile_X0Y0_N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 56.670 519.240 56.950 519.520 ;
    END
  END Tile_X0Y0_N4BEG[11]
  PIN Tile_X0Y0_N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 519.240 58.330 519.520 ;
    END
  END Tile_X0Y0_N4BEG[12]
  PIN Tile_X0Y0_N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 59.430 519.240 59.710 519.520 ;
    END
  END Tile_X0Y0_N4BEG[13]
  PIN Tile_X0Y0_N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 60.810 519.240 61.090 519.520 ;
    END
  END Tile_X0Y0_N4BEG[14]
  PIN Tile_X0Y0_N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 62.190 519.240 62.470 519.520 ;
    END
  END Tile_X0Y0_N4BEG[15]
  PIN Tile_X0Y0_N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 42.870 519.240 43.150 519.520 ;
    END
  END Tile_X0Y0_N4BEG[1]
  PIN Tile_X0Y0_N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 44.250 519.240 44.530 519.520 ;
    END
  END Tile_X0Y0_N4BEG[2]
  PIN Tile_X0Y0_N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.630 519.240 45.910 519.520 ;
    END
  END Tile_X0Y0_N4BEG[3]
  PIN Tile_X0Y0_N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 47.010 519.240 47.290 519.520 ;
    END
  END Tile_X0Y0_N4BEG[4]
  PIN Tile_X0Y0_N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 519.240 48.670 519.520 ;
    END
  END Tile_X0Y0_N4BEG[5]
  PIN Tile_X0Y0_N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 49.770 519.240 50.050 519.520 ;
    END
  END Tile_X0Y0_N4BEG[6]
  PIN Tile_X0Y0_N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.150 519.240 51.430 519.520 ;
    END
  END Tile_X0Y0_N4BEG[7]
  PIN Tile_X0Y0_N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.530 519.240 52.810 519.520 ;
    END
  END Tile_X0Y0_N4BEG[8]
  PIN Tile_X0Y0_N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 53.910 519.240 54.190 519.520 ;
    END
  END Tile_X0Y0_N4BEG[9]
  PIN Tile_X0Y0_NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 63.570 519.240 63.850 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[0]
  PIN Tile_X0Y0_NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 519.240 77.650 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[10]
  PIN Tile_X0Y0_NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 78.750 519.240 79.030 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[11]
  PIN Tile_X0Y0_NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.130 519.240 80.410 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[12]
  PIN Tile_X0Y0_NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 81.510 519.240 81.790 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[13]
  PIN Tile_X0Y0_NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 82.890 519.240 83.170 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[14]
  PIN Tile_X0Y0_NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 84.270 519.240 84.550 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[15]
  PIN Tile_X0Y0_NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.950 519.240 65.230 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[1]
  PIN Tile_X0Y0_NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 66.330 519.240 66.610 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[2]
  PIN Tile_X0Y0_NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 519.240 67.990 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[3]
  PIN Tile_X0Y0_NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 69.090 519.240 69.370 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[4]
  PIN Tile_X0Y0_NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.470 519.240 70.750 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[5]
  PIN Tile_X0Y0_NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 71.850 519.240 72.130 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[6]
  PIN Tile_X0Y0_NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 73.230 519.240 73.510 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[7]
  PIN Tile_X0Y0_NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.610 519.240 74.890 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[8]
  PIN Tile_X0Y0_NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 75.990 519.240 76.270 519.520 ;
    END
  END Tile_X0Y0_NN4BEG[9]
  PIN Tile_X0Y0_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 85.650 519.240 85.930 519.520 ;
    END
  END Tile_X0Y0_S1END[0]
  PIN Tile_X0Y0_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 519.240 87.310 519.520 ;
    END
  END Tile_X0Y0_S1END[1]
  PIN Tile_X0Y0_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 88.410 519.240 88.690 519.520 ;
    END
  END Tile_X0Y0_S1END[2]
  PIN Tile_X0Y0_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 89.790 519.240 90.070 519.520 ;
    END
  END Tile_X0Y0_S1END[3]
  PIN Tile_X0Y0_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 102.210 519.240 102.490 519.520 ;
    END
  END Tile_X0Y0_S2END[0]
  PIN Tile_X0Y0_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 103.590 519.240 103.870 519.520 ;
    END
  END Tile_X0Y0_S2END[1]
  PIN Tile_X0Y0_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 104.970 519.240 105.250 519.520 ;
    END
  END Tile_X0Y0_S2END[2]
  PIN Tile_X0Y0_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 106.350 519.240 106.630 519.520 ;
    END
  END Tile_X0Y0_S2END[3]
  PIN Tile_X0Y0_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 107.730 519.240 108.010 519.520 ;
    END
  END Tile_X0Y0_S2END[4]
  PIN Tile_X0Y0_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 109.110 519.240 109.390 519.520 ;
    END
  END Tile_X0Y0_S2END[5]
  PIN Tile_X0Y0_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 110.490 519.240 110.770 519.520 ;
    END
  END Tile_X0Y0_S2END[6]
  PIN Tile_X0Y0_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 111.870 519.240 112.150 519.520 ;
    END
  END Tile_X0Y0_S2END[7]
  PIN Tile_X0Y0_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 91.170 519.240 91.450 519.520 ;
    END
  END Tile_X0Y0_S2MID[0]
  PIN Tile_X0Y0_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 519.240 92.830 519.520 ;
    END
  END Tile_X0Y0_S2MID[1]
  PIN Tile_X0Y0_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 93.930 519.240 94.210 519.520 ;
    END
  END Tile_X0Y0_S2MID[2]
  PIN Tile_X0Y0_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 95.310 519.240 95.590 519.520 ;
    END
  END Tile_X0Y0_S2MID[3]
  PIN Tile_X0Y0_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 519.240 96.970 519.520 ;
    END
  END Tile_X0Y0_S2MID[4]
  PIN Tile_X0Y0_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 98.070 519.240 98.350 519.520 ;
    END
  END Tile_X0Y0_S2MID[5]
  PIN Tile_X0Y0_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 99.450 519.240 99.730 519.520 ;
    END
  END Tile_X0Y0_S2MID[6]
  PIN Tile_X0Y0_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 100.830 519.240 101.110 519.520 ;
    END
  END Tile_X0Y0_S2MID[7]
  PIN Tile_X0Y0_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 113.250 519.240 113.530 519.520 ;
    END
  END Tile_X0Y0_S4END[0]
  PIN Tile_X0Y0_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 127.050 519.240 127.330 519.520 ;
    END
  END Tile_X0Y0_S4END[10]
  PIN Tile_X0Y0_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 128.430 519.240 128.710 519.520 ;
    END
  END Tile_X0Y0_S4END[11]
  PIN Tile_X0Y0_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 519.240 130.090 519.520 ;
    END
  END Tile_X0Y0_S4END[12]
  PIN Tile_X0Y0_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 131.190 519.240 131.470 519.520 ;
    END
  END Tile_X0Y0_S4END[13]
  PIN Tile_X0Y0_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 132.570 519.240 132.850 519.520 ;
    END
  END Tile_X0Y0_S4END[14]
  PIN Tile_X0Y0_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 133.950 519.240 134.230 519.520 ;
    END
  END Tile_X0Y0_S4END[15]
  PIN Tile_X0Y0_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 114.630 519.240 114.910 519.520 ;
    END
  END Tile_X0Y0_S4END[1]
  PIN Tile_X0Y0_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 519.240 116.290 519.520 ;
    END
  END Tile_X0Y0_S4END[2]
  PIN Tile_X0Y0_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 117.390 519.240 117.670 519.520 ;
    END
  END Tile_X0Y0_S4END[3]
  PIN Tile_X0Y0_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 118.770 519.240 119.050 519.520 ;
    END
  END Tile_X0Y0_S4END[4]
  PIN Tile_X0Y0_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 120.150 519.240 120.430 519.520 ;
    END
  END Tile_X0Y0_S4END[5]
  PIN Tile_X0Y0_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 121.530 519.240 121.810 519.520 ;
    END
  END Tile_X0Y0_S4END[6]
  PIN Tile_X0Y0_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 122.910 519.240 123.190 519.520 ;
    END
  END Tile_X0Y0_S4END[7]
  PIN Tile_X0Y0_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 124.290 519.240 124.570 519.520 ;
    END
  END Tile_X0Y0_S4END[8]
  PIN Tile_X0Y0_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 519.240 125.950 519.520 ;
    END
  END Tile_X0Y0_S4END[9]
  PIN Tile_X0Y0_SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 519.240 135.610 519.520 ;
    END
  END Tile_X0Y0_SS4END[0]
  PIN Tile_X0Y0_SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 149.130 519.240 149.410 519.520 ;
    END
  END Tile_X0Y0_SS4END[10]
  PIN Tile_X0Y0_SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 150.510 519.240 150.790 519.520 ;
    END
  END Tile_X0Y0_SS4END[11]
  PIN Tile_X0Y0_SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 151.890 519.240 152.170 519.520 ;
    END
  END Tile_X0Y0_SS4END[12]
  PIN Tile_X0Y0_SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 153.270 519.240 153.550 519.520 ;
    END
  END Tile_X0Y0_SS4END[13]
  PIN Tile_X0Y0_SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 519.240 154.930 519.520 ;
    END
  END Tile_X0Y0_SS4END[14]
  PIN Tile_X0Y0_SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 156.030 519.240 156.310 519.520 ;
    END
  END Tile_X0Y0_SS4END[15]
  PIN Tile_X0Y0_SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 136.710 519.240 136.990 519.520 ;
    END
  END Tile_X0Y0_SS4END[1]
  PIN Tile_X0Y0_SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 519.240 138.370 519.520 ;
    END
  END Tile_X0Y0_SS4END[2]
  PIN Tile_X0Y0_SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 139.470 519.240 139.750 519.520 ;
    END
  END Tile_X0Y0_SS4END[3]
  PIN Tile_X0Y0_SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 140.850 519.240 141.130 519.520 ;
    END
  END Tile_X0Y0_SS4END[4]
  PIN Tile_X0Y0_SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 142.230 519.240 142.510 519.520 ;
    END
  END Tile_X0Y0_SS4END[5]
  PIN Tile_X0Y0_SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 143.610 519.240 143.890 519.520 ;
    END
  END Tile_X0Y0_SS4END[6]
  PIN Tile_X0Y0_SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 519.240 145.270 519.520 ;
    END
  END Tile_X0Y0_SS4END[7]
  PIN Tile_X0Y0_SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 146.370 519.240 146.650 519.520 ;
    END
  END Tile_X0Y0_SS4END[8]
  PIN Tile_X0Y0_SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 147.750 519.240 148.030 519.520 ;
    END
  END Tile_X0Y0_SS4END[9]
  PIN Tile_X0Y0_UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 157.410 519.240 157.690 519.520 ;
    END
  END Tile_X0Y0_UserCLKo
  PIN Tile_X0Y0_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 0.600 302.560 ;
    END
  END Tile_X0Y0_W1BEG[0]
  PIN Tile_X0Y0_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 0.600 303.920 ;
    END
  END Tile_X0Y0_W1BEG[1]
  PIN Tile_X0Y0_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 0.600 305.280 ;
    END
  END Tile_X0Y0_W1BEG[2]
  PIN Tile_X0Y0_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 0.600 306.640 ;
    END
  END Tile_X0Y0_W1BEG[3]
  PIN Tile_X0Y0_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 301.960 199.640 302.560 ;
    END
  END Tile_X0Y0_W1END[0]
  PIN Tile_X0Y0_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 303.320 199.640 303.920 ;
    END
  END Tile_X0Y0_W1END[1]
  PIN Tile_X0Y0_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 304.680 199.640 305.280 ;
    END
  END Tile_X0Y0_W1END[2]
  PIN Tile_X0Y0_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 306.040 199.640 306.640 ;
    END
  END Tile_X0Y0_W1END[3]
  PIN Tile_X0Y0_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 0.600 308.000 ;
    END
  END Tile_X0Y0_W2BEG[0]
  PIN Tile_X0Y0_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 0.600 309.360 ;
    END
  END Tile_X0Y0_W2BEG[1]
  PIN Tile_X0Y0_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 0.600 310.720 ;
    END
  END Tile_X0Y0_W2BEG[2]
  PIN Tile_X0Y0_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 0.600 312.080 ;
    END
  END Tile_X0Y0_W2BEG[3]
  PIN Tile_X0Y0_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 0.600 313.440 ;
    END
  END Tile_X0Y0_W2BEG[4]
  PIN Tile_X0Y0_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 0.600 314.800 ;
    END
  END Tile_X0Y0_W2BEG[5]
  PIN Tile_X0Y0_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 0.600 316.160 ;
    END
  END Tile_X0Y0_W2BEG[6]
  PIN Tile_X0Y0_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 0.600 317.520 ;
    END
  END Tile_X0Y0_W2BEG[7]
  PIN Tile_X0Y0_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 0.600 318.880 ;
    END
  END Tile_X0Y0_W2BEGb[0]
  PIN Tile_X0Y0_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 0.600 320.240 ;
    END
  END Tile_X0Y0_W2BEGb[1]
  PIN Tile_X0Y0_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 0.600 321.600 ;
    END
  END Tile_X0Y0_W2BEGb[2]
  PIN Tile_X0Y0_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 0.600 322.960 ;
    END
  END Tile_X0Y0_W2BEGb[3]
  PIN Tile_X0Y0_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 0.600 324.320 ;
    END
  END Tile_X0Y0_W2BEGb[4]
  PIN Tile_X0Y0_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 0.600 325.680 ;
    END
  END Tile_X0Y0_W2BEGb[5]
  PIN Tile_X0Y0_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 0.600 327.040 ;
    END
  END Tile_X0Y0_W2BEGb[6]
  PIN Tile_X0Y0_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 0.600 328.400 ;
    END
  END Tile_X0Y0_W2BEGb[7]
  PIN Tile_X0Y0_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 318.280 199.640 318.880 ;
    END
  END Tile_X0Y0_W2END[0]
  PIN Tile_X0Y0_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 319.640 199.640 320.240 ;
    END
  END Tile_X0Y0_W2END[1]
  PIN Tile_X0Y0_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 321.000 199.640 321.600 ;
    END
  END Tile_X0Y0_W2END[2]
  PIN Tile_X0Y0_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 322.360 199.640 322.960 ;
    END
  END Tile_X0Y0_W2END[3]
  PIN Tile_X0Y0_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 323.720 199.640 324.320 ;
    END
  END Tile_X0Y0_W2END[4]
  PIN Tile_X0Y0_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 325.080 199.640 325.680 ;
    END
  END Tile_X0Y0_W2END[5]
  PIN Tile_X0Y0_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 326.440 199.640 327.040 ;
    END
  END Tile_X0Y0_W2END[6]
  PIN Tile_X0Y0_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 327.800 199.640 328.400 ;
    END
  END Tile_X0Y0_W2END[7]
  PIN Tile_X0Y0_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 307.400 199.640 308.000 ;
    END
  END Tile_X0Y0_W2MID[0]
  PIN Tile_X0Y0_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 308.760 199.640 309.360 ;
    END
  END Tile_X0Y0_W2MID[1]
  PIN Tile_X0Y0_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 310.120 199.640 310.720 ;
    END
  END Tile_X0Y0_W2MID[2]
  PIN Tile_X0Y0_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 311.480 199.640 312.080 ;
    END
  END Tile_X0Y0_W2MID[3]
  PIN Tile_X0Y0_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 312.840 199.640 313.440 ;
    END
  END Tile_X0Y0_W2MID[4]
  PIN Tile_X0Y0_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 314.200 199.640 314.800 ;
    END
  END Tile_X0Y0_W2MID[5]
  PIN Tile_X0Y0_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 315.560 199.640 316.160 ;
    END
  END Tile_X0Y0_W2MID[6]
  PIN Tile_X0Y0_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 316.920 199.640 317.520 ;
    END
  END Tile_X0Y0_W2MID[7]
  PIN Tile_X0Y0_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 0.600 351.520 ;
    END
  END Tile_X0Y0_W6BEG[0]
  PIN Tile_X0Y0_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 0.600 365.120 ;
    END
  END Tile_X0Y0_W6BEG[10]
  PIN Tile_X0Y0_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 0.600 366.480 ;
    END
  END Tile_X0Y0_W6BEG[11]
  PIN Tile_X0Y0_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 0.600 352.880 ;
    END
  END Tile_X0Y0_W6BEG[1]
  PIN Tile_X0Y0_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 0.600 354.240 ;
    END
  END Tile_X0Y0_W6BEG[2]
  PIN Tile_X0Y0_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 0.600 355.600 ;
    END
  END Tile_X0Y0_W6BEG[3]
  PIN Tile_X0Y0_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 0.600 356.960 ;
    END
  END Tile_X0Y0_W6BEG[4]
  PIN Tile_X0Y0_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 0.600 358.320 ;
    END
  END Tile_X0Y0_W6BEG[5]
  PIN Tile_X0Y0_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 0.600 359.680 ;
    END
  END Tile_X0Y0_W6BEG[6]
  PIN Tile_X0Y0_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 0.600 361.040 ;
    END
  END Tile_X0Y0_W6BEG[7]
  PIN Tile_X0Y0_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 0.600 362.400 ;
    END
  END Tile_X0Y0_W6BEG[8]
  PIN Tile_X0Y0_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 0.600 363.760 ;
    END
  END Tile_X0Y0_W6BEG[9]
  PIN Tile_X0Y0_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 350.920 199.640 351.520 ;
    END
  END Tile_X0Y0_W6END[0]
  PIN Tile_X0Y0_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 364.520 199.640 365.120 ;
    END
  END Tile_X0Y0_W6END[10]
  PIN Tile_X0Y0_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 365.880 199.640 366.480 ;
    END
  END Tile_X0Y0_W6END[11]
  PIN Tile_X0Y0_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 352.280 199.640 352.880 ;
    END
  END Tile_X0Y0_W6END[1]
  PIN Tile_X0Y0_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 353.640 199.640 354.240 ;
    END
  END Tile_X0Y0_W6END[2]
  PIN Tile_X0Y0_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 355.000 199.640 355.600 ;
    END
  END Tile_X0Y0_W6END[3]
  PIN Tile_X0Y0_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 356.360 199.640 356.960 ;
    END
  END Tile_X0Y0_W6END[4]
  PIN Tile_X0Y0_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 357.720 199.640 358.320 ;
    END
  END Tile_X0Y0_W6END[5]
  PIN Tile_X0Y0_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 359.080 199.640 359.680 ;
    END
  END Tile_X0Y0_W6END[6]
  PIN Tile_X0Y0_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 360.440 199.640 361.040 ;
    END
  END Tile_X0Y0_W6END[7]
  PIN Tile_X0Y0_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 361.800 199.640 362.400 ;
    END
  END Tile_X0Y0_W6END[8]
  PIN Tile_X0Y0_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 363.160 199.640 363.760 ;
    END
  END Tile_X0Y0_W6END[9]
  PIN Tile_X0Y0_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 0.600 329.760 ;
    END
  END Tile_X0Y0_WW4BEG[0]
  PIN Tile_X0Y0_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 0.600 343.360 ;
    END
  END Tile_X0Y0_WW4BEG[10]
  PIN Tile_X0Y0_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 0.600 344.720 ;
    END
  END Tile_X0Y0_WW4BEG[11]
  PIN Tile_X0Y0_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 0.600 346.080 ;
    END
  END Tile_X0Y0_WW4BEG[12]
  PIN Tile_X0Y0_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 0.600 347.440 ;
    END
  END Tile_X0Y0_WW4BEG[13]
  PIN Tile_X0Y0_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 0.600 348.800 ;
    END
  END Tile_X0Y0_WW4BEG[14]
  PIN Tile_X0Y0_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 0.600 350.160 ;
    END
  END Tile_X0Y0_WW4BEG[15]
  PIN Tile_X0Y0_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 0.600 331.120 ;
    END
  END Tile_X0Y0_WW4BEG[1]
  PIN Tile_X0Y0_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 0.600 332.480 ;
    END
  END Tile_X0Y0_WW4BEG[2]
  PIN Tile_X0Y0_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 0.600 333.840 ;
    END
  END Tile_X0Y0_WW4BEG[3]
  PIN Tile_X0Y0_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 0.600 335.200 ;
    END
  END Tile_X0Y0_WW4BEG[4]
  PIN Tile_X0Y0_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 0.600 336.560 ;
    END
  END Tile_X0Y0_WW4BEG[5]
  PIN Tile_X0Y0_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 0.600 337.920 ;
    END
  END Tile_X0Y0_WW4BEG[6]
  PIN Tile_X0Y0_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 0.600 339.280 ;
    END
  END Tile_X0Y0_WW4BEG[7]
  PIN Tile_X0Y0_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 0.600 340.640 ;
    END
  END Tile_X0Y0_WW4BEG[8]
  PIN Tile_X0Y0_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 0.600 342.000 ;
    END
  END Tile_X0Y0_WW4BEG[9]
  PIN Tile_X0Y0_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 329.160 199.640 329.760 ;
    END
  END Tile_X0Y0_WW4END[0]
  PIN Tile_X0Y0_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 342.760 199.640 343.360 ;
    END
  END Tile_X0Y0_WW4END[10]
  PIN Tile_X0Y0_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 344.120 199.640 344.720 ;
    END
  END Tile_X0Y0_WW4END[11]
  PIN Tile_X0Y0_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 345.480 199.640 346.080 ;
    END
  END Tile_X0Y0_WW4END[12]
  PIN Tile_X0Y0_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 346.840 199.640 347.440 ;
    END
  END Tile_X0Y0_WW4END[13]
  PIN Tile_X0Y0_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 348.200 199.640 348.800 ;
    END
  END Tile_X0Y0_WW4END[14]
  PIN Tile_X0Y0_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 349.560 199.640 350.160 ;
    END
  END Tile_X0Y0_WW4END[15]
  PIN Tile_X0Y0_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 330.520 199.640 331.120 ;
    END
  END Tile_X0Y0_WW4END[1]
  PIN Tile_X0Y0_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 331.880 199.640 332.480 ;
    END
  END Tile_X0Y0_WW4END[2]
  PIN Tile_X0Y0_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 333.240 199.640 333.840 ;
    END
  END Tile_X0Y0_WW4END[3]
  PIN Tile_X0Y0_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 334.600 199.640 335.200 ;
    END
  END Tile_X0Y0_WW4END[4]
  PIN Tile_X0Y0_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 335.960 199.640 336.560 ;
    END
  END Tile_X0Y0_WW4END[5]
  PIN Tile_X0Y0_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 337.320 199.640 337.920 ;
    END
  END Tile_X0Y0_WW4END[6]
  PIN Tile_X0Y0_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 338.680 199.640 339.280 ;
    END
  END Tile_X0Y0_WW4END[7]
  PIN Tile_X0Y0_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 340.040 199.640 340.640 ;
    END
  END Tile_X0Y0_WW4END[8]
  PIN Tile_X0Y0_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 341.400 199.640 342.000 ;
    END
  END Tile_X0Y0_WW4END[9]
  PIN Tile_X0Y1_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 107.480 199.640 108.080 ;
    END
  END Tile_X0Y1_E1BEG[0]
  PIN Tile_X0Y1_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 108.840 199.640 109.440 ;
    END
  END Tile_X0Y1_E1BEG[1]
  PIN Tile_X0Y1_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 110.200 199.640 110.800 ;
    END
  END Tile_X0Y1_E1BEG[2]
  PIN Tile_X0Y1_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 111.560 199.640 112.160 ;
    END
  END Tile_X0Y1_E1BEG[3]
  PIN Tile_X0Y1_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 0.600 108.080 ;
    END
  END Tile_X0Y1_E1END[0]
  PIN Tile_X0Y1_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 0.600 109.440 ;
    END
  END Tile_X0Y1_E1END[1]
  PIN Tile_X0Y1_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 0.600 110.800 ;
    END
  END Tile_X0Y1_E1END[2]
  PIN Tile_X0Y1_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 0.600 112.160 ;
    END
  END Tile_X0Y1_E1END[3]
  PIN Tile_X0Y1_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 112.920 199.640 113.520 ;
    END
  END Tile_X0Y1_E2BEG[0]
  PIN Tile_X0Y1_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 114.280 199.640 114.880 ;
    END
  END Tile_X0Y1_E2BEG[1]
  PIN Tile_X0Y1_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 115.640 199.640 116.240 ;
    END
  END Tile_X0Y1_E2BEG[2]
  PIN Tile_X0Y1_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 117.000 199.640 117.600 ;
    END
  END Tile_X0Y1_E2BEG[3]
  PIN Tile_X0Y1_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 118.360 199.640 118.960 ;
    END
  END Tile_X0Y1_E2BEG[4]
  PIN Tile_X0Y1_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 119.720 199.640 120.320 ;
    END
  END Tile_X0Y1_E2BEG[5]
  PIN Tile_X0Y1_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 121.080 199.640 121.680 ;
    END
  END Tile_X0Y1_E2BEG[6]
  PIN Tile_X0Y1_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 122.440 199.640 123.040 ;
    END
  END Tile_X0Y1_E2BEG[7]
  PIN Tile_X0Y1_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 123.800 199.640 124.400 ;
    END
  END Tile_X0Y1_E2BEGb[0]
  PIN Tile_X0Y1_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 125.160 199.640 125.760 ;
    END
  END Tile_X0Y1_E2BEGb[1]
  PIN Tile_X0Y1_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 126.520 199.640 127.120 ;
    END
  END Tile_X0Y1_E2BEGb[2]
  PIN Tile_X0Y1_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 127.880 199.640 128.480 ;
    END
  END Tile_X0Y1_E2BEGb[3]
  PIN Tile_X0Y1_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 129.240 199.640 129.840 ;
    END
  END Tile_X0Y1_E2BEGb[4]
  PIN Tile_X0Y1_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 130.600 199.640 131.200 ;
    END
  END Tile_X0Y1_E2BEGb[5]
  PIN Tile_X0Y1_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 131.960 199.640 132.560 ;
    END
  END Tile_X0Y1_E2BEGb[6]
  PIN Tile_X0Y1_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 133.320 199.640 133.920 ;
    END
  END Tile_X0Y1_E2BEGb[7]
  PIN Tile_X0Y1_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 0.600 124.400 ;
    END
  END Tile_X0Y1_E2END[0]
  PIN Tile_X0Y1_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 0.600 125.760 ;
    END
  END Tile_X0Y1_E2END[1]
  PIN Tile_X0Y1_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 0.600 127.120 ;
    END
  END Tile_X0Y1_E2END[2]
  PIN Tile_X0Y1_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 0.600 128.480 ;
    END
  END Tile_X0Y1_E2END[3]
  PIN Tile_X0Y1_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 0.600 129.840 ;
    END
  END Tile_X0Y1_E2END[4]
  PIN Tile_X0Y1_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 0.600 131.200 ;
    END
  END Tile_X0Y1_E2END[5]
  PIN Tile_X0Y1_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 0.600 132.560 ;
    END
  END Tile_X0Y1_E2END[6]
  PIN Tile_X0Y1_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 0.600 133.920 ;
    END
  END Tile_X0Y1_E2END[7]
  PIN Tile_X0Y1_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 0.600 113.520 ;
    END
  END Tile_X0Y1_E2MID[0]
  PIN Tile_X0Y1_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 0.600 114.880 ;
    END
  END Tile_X0Y1_E2MID[1]
  PIN Tile_X0Y1_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 0.600 116.240 ;
    END
  END Tile_X0Y1_E2MID[2]
  PIN Tile_X0Y1_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 0.600 117.600 ;
    END
  END Tile_X0Y1_E2MID[3]
  PIN Tile_X0Y1_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 0.600 118.960 ;
    END
  END Tile_X0Y1_E2MID[4]
  PIN Tile_X0Y1_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 0.600 120.320 ;
    END
  END Tile_X0Y1_E2MID[5]
  PIN Tile_X0Y1_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 0.600 121.680 ;
    END
  END Tile_X0Y1_E2MID[6]
  PIN Tile_X0Y1_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 0.600 123.040 ;
    END
  END Tile_X0Y1_E2MID[7]
  PIN Tile_X0Y1_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 156.440 199.640 157.040 ;
    END
  END Tile_X0Y1_E6BEG[0]
  PIN Tile_X0Y1_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 170.040 199.640 170.640 ;
    END
  END Tile_X0Y1_E6BEG[10]
  PIN Tile_X0Y1_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 171.400 199.640 172.000 ;
    END
  END Tile_X0Y1_E6BEG[11]
  PIN Tile_X0Y1_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 157.800 199.640 158.400 ;
    END
  END Tile_X0Y1_E6BEG[1]
  PIN Tile_X0Y1_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 159.160 199.640 159.760 ;
    END
  END Tile_X0Y1_E6BEG[2]
  PIN Tile_X0Y1_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 160.520 199.640 161.120 ;
    END
  END Tile_X0Y1_E6BEG[3]
  PIN Tile_X0Y1_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 161.880 199.640 162.480 ;
    END
  END Tile_X0Y1_E6BEG[4]
  PIN Tile_X0Y1_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 163.240 199.640 163.840 ;
    END
  END Tile_X0Y1_E6BEG[5]
  PIN Tile_X0Y1_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 164.600 199.640 165.200 ;
    END
  END Tile_X0Y1_E6BEG[6]
  PIN Tile_X0Y1_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 165.960 199.640 166.560 ;
    END
  END Tile_X0Y1_E6BEG[7]
  PIN Tile_X0Y1_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 167.320 199.640 167.920 ;
    END
  END Tile_X0Y1_E6BEG[8]
  PIN Tile_X0Y1_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 168.680 199.640 169.280 ;
    END
  END Tile_X0Y1_E6BEG[9]
  PIN Tile_X0Y1_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 0.600 157.040 ;
    END
  END Tile_X0Y1_E6END[0]
  PIN Tile_X0Y1_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 0.600 170.640 ;
    END
  END Tile_X0Y1_E6END[10]
  PIN Tile_X0Y1_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 0.600 172.000 ;
    END
  END Tile_X0Y1_E6END[11]
  PIN Tile_X0Y1_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 0.600 158.400 ;
    END
  END Tile_X0Y1_E6END[1]
  PIN Tile_X0Y1_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 0.600 159.760 ;
    END
  END Tile_X0Y1_E6END[2]
  PIN Tile_X0Y1_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 0.600 161.120 ;
    END
  END Tile_X0Y1_E6END[3]
  PIN Tile_X0Y1_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 0.600 162.480 ;
    END
  END Tile_X0Y1_E6END[4]
  PIN Tile_X0Y1_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 0.600 163.840 ;
    END
  END Tile_X0Y1_E6END[5]
  PIN Tile_X0Y1_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 0.600 165.200 ;
    END
  END Tile_X0Y1_E6END[6]
  PIN Tile_X0Y1_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 0.600 166.560 ;
    END
  END Tile_X0Y1_E6END[7]
  PIN Tile_X0Y1_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 0.600 167.920 ;
    END
  END Tile_X0Y1_E6END[8]
  PIN Tile_X0Y1_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 0.600 169.280 ;
    END
  END Tile_X0Y1_E6END[9]
  PIN Tile_X0Y1_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 134.680 199.640 135.280 ;
    END
  END Tile_X0Y1_EE4BEG[0]
  PIN Tile_X0Y1_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 148.280 199.640 148.880 ;
    END
  END Tile_X0Y1_EE4BEG[10]
  PIN Tile_X0Y1_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 149.640 199.640 150.240 ;
    END
  END Tile_X0Y1_EE4BEG[11]
  PIN Tile_X0Y1_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 151.000 199.640 151.600 ;
    END
  END Tile_X0Y1_EE4BEG[12]
  PIN Tile_X0Y1_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 152.360 199.640 152.960 ;
    END
  END Tile_X0Y1_EE4BEG[13]
  PIN Tile_X0Y1_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 153.720 199.640 154.320 ;
    END
  END Tile_X0Y1_EE4BEG[14]
  PIN Tile_X0Y1_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 155.080 199.640 155.680 ;
    END
  END Tile_X0Y1_EE4BEG[15]
  PIN Tile_X0Y1_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 136.040 199.640 136.640 ;
    END
  END Tile_X0Y1_EE4BEG[1]
  PIN Tile_X0Y1_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 137.400 199.640 138.000 ;
    END
  END Tile_X0Y1_EE4BEG[2]
  PIN Tile_X0Y1_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 138.760 199.640 139.360 ;
    END
  END Tile_X0Y1_EE4BEG[3]
  PIN Tile_X0Y1_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 140.120 199.640 140.720 ;
    END
  END Tile_X0Y1_EE4BEG[4]
  PIN Tile_X0Y1_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 141.480 199.640 142.080 ;
    END
  END Tile_X0Y1_EE4BEG[5]
  PIN Tile_X0Y1_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 142.840 199.640 143.440 ;
    END
  END Tile_X0Y1_EE4BEG[6]
  PIN Tile_X0Y1_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 144.200 199.640 144.800 ;
    END
  END Tile_X0Y1_EE4BEG[7]
  PIN Tile_X0Y1_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 145.560 199.640 146.160 ;
    END
  END Tile_X0Y1_EE4BEG[8]
  PIN Tile_X0Y1_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 146.920 199.640 147.520 ;
    END
  END Tile_X0Y1_EE4BEG[9]
  PIN Tile_X0Y1_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 0.600 135.280 ;
    END
  END Tile_X0Y1_EE4END[0]
  PIN Tile_X0Y1_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 0.600 148.880 ;
    END
  END Tile_X0Y1_EE4END[10]
  PIN Tile_X0Y1_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 0.600 150.240 ;
    END
  END Tile_X0Y1_EE4END[11]
  PIN Tile_X0Y1_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 0.600 151.600 ;
    END
  END Tile_X0Y1_EE4END[12]
  PIN Tile_X0Y1_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 0.600 152.960 ;
    END
  END Tile_X0Y1_EE4END[13]
  PIN Tile_X0Y1_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 0.600 154.320 ;
    END
  END Tile_X0Y1_EE4END[14]
  PIN Tile_X0Y1_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 0.600 155.680 ;
    END
  END Tile_X0Y1_EE4END[15]
  PIN Tile_X0Y1_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 0.600 136.640 ;
    END
  END Tile_X0Y1_EE4END[1]
  PIN Tile_X0Y1_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 0.600 138.000 ;
    END
  END Tile_X0Y1_EE4END[2]
  PIN Tile_X0Y1_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 0.600 139.360 ;
    END
  END Tile_X0Y1_EE4END[3]
  PIN Tile_X0Y1_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 0.600 140.720 ;
    END
  END Tile_X0Y1_EE4END[4]
  PIN Tile_X0Y1_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 0.600 142.080 ;
    END
  END Tile_X0Y1_EE4END[5]
  PIN Tile_X0Y1_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 0.600 143.440 ;
    END
  END Tile_X0Y1_EE4END[6]
  PIN Tile_X0Y1_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 0.600 144.800 ;
    END
  END Tile_X0Y1_EE4END[7]
  PIN Tile_X0Y1_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 0.600 146.160 ;
    END
  END Tile_X0Y1_EE4END[8]
  PIN Tile_X0Y1_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 0.600 147.520 ;
    END
  END Tile_X0Y1_EE4END[9]
  PIN Tile_X0Y1_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 0.600 173.360 ;
    END
  END Tile_X0Y1_FrameData[0]
  PIN Tile_X0Y1_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 0.600 186.960 ;
    END
  END Tile_X0Y1_FrameData[10]
  PIN Tile_X0Y1_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 0.600 188.320 ;
    END
  END Tile_X0Y1_FrameData[11]
  PIN Tile_X0Y1_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 0.600 189.680 ;
    END
  END Tile_X0Y1_FrameData[12]
  PIN Tile_X0Y1_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 0.600 191.040 ;
    END
  END Tile_X0Y1_FrameData[13]
  PIN Tile_X0Y1_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 0.600 192.400 ;
    END
  END Tile_X0Y1_FrameData[14]
  PIN Tile_X0Y1_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 0.600 193.760 ;
    END
  END Tile_X0Y1_FrameData[15]
  PIN Tile_X0Y1_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 0.600 195.120 ;
    END
  END Tile_X0Y1_FrameData[16]
  PIN Tile_X0Y1_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 0.600 196.480 ;
    END
  END Tile_X0Y1_FrameData[17]
  PIN Tile_X0Y1_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 0.600 197.840 ;
    END
  END Tile_X0Y1_FrameData[18]
  PIN Tile_X0Y1_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 0.600 199.200 ;
    END
  END Tile_X0Y1_FrameData[19]
  PIN Tile_X0Y1_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 0.600 174.720 ;
    END
  END Tile_X0Y1_FrameData[1]
  PIN Tile_X0Y1_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 0.600 200.560 ;
    END
  END Tile_X0Y1_FrameData[20]
  PIN Tile_X0Y1_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 0.600 201.920 ;
    END
  END Tile_X0Y1_FrameData[21]
  PIN Tile_X0Y1_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 0.600 203.280 ;
    END
  END Tile_X0Y1_FrameData[22]
  PIN Tile_X0Y1_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 0.600 204.640 ;
    END
  END Tile_X0Y1_FrameData[23]
  PIN Tile_X0Y1_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 0.600 206.000 ;
    END
  END Tile_X0Y1_FrameData[24]
  PIN Tile_X0Y1_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 0.600 207.360 ;
    END
  END Tile_X0Y1_FrameData[25]
  PIN Tile_X0Y1_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 0.600 208.720 ;
    END
  END Tile_X0Y1_FrameData[26]
  PIN Tile_X0Y1_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 0.600 210.080 ;
    END
  END Tile_X0Y1_FrameData[27]
  PIN Tile_X0Y1_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 0.600 211.440 ;
    END
  END Tile_X0Y1_FrameData[28]
  PIN Tile_X0Y1_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 0.600 212.800 ;
    END
  END Tile_X0Y1_FrameData[29]
  PIN Tile_X0Y1_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 0.600 176.080 ;
    END
  END Tile_X0Y1_FrameData[2]
  PIN Tile_X0Y1_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 0.600 214.160 ;
    END
  END Tile_X0Y1_FrameData[30]
  PIN Tile_X0Y1_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 0.600 215.520 ;
    END
  END Tile_X0Y1_FrameData[31]
  PIN Tile_X0Y1_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 0.600 177.440 ;
    END
  END Tile_X0Y1_FrameData[3]
  PIN Tile_X0Y1_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 0.600 178.800 ;
    END
  END Tile_X0Y1_FrameData[4]
  PIN Tile_X0Y1_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 0.600 180.160 ;
    END
  END Tile_X0Y1_FrameData[5]
  PIN Tile_X0Y1_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 0.600 181.520 ;
    END
  END Tile_X0Y1_FrameData[6]
  PIN Tile_X0Y1_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 0.600 182.880 ;
    END
  END Tile_X0Y1_FrameData[7]
  PIN Tile_X0Y1_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 0.600 184.240 ;
    END
  END Tile_X0Y1_FrameData[8]
  PIN Tile_X0Y1_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 0.600 185.600 ;
    END
  END Tile_X0Y1_FrameData[9]
  PIN Tile_X0Y1_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 172.760 199.640 173.360 ;
    END
  END Tile_X0Y1_FrameData_O[0]
  PIN Tile_X0Y1_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 186.360 199.640 186.960 ;
    END
  END Tile_X0Y1_FrameData_O[10]
  PIN Tile_X0Y1_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 187.720 199.640 188.320 ;
    END
  END Tile_X0Y1_FrameData_O[11]
  PIN Tile_X0Y1_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 189.080 199.640 189.680 ;
    END
  END Tile_X0Y1_FrameData_O[12]
  PIN Tile_X0Y1_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 190.440 199.640 191.040 ;
    END
  END Tile_X0Y1_FrameData_O[13]
  PIN Tile_X0Y1_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 191.800 199.640 192.400 ;
    END
  END Tile_X0Y1_FrameData_O[14]
  PIN Tile_X0Y1_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 193.160 199.640 193.760 ;
    END
  END Tile_X0Y1_FrameData_O[15]
  PIN Tile_X0Y1_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 194.520 199.640 195.120 ;
    END
  END Tile_X0Y1_FrameData_O[16]
  PIN Tile_X0Y1_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 195.880 199.640 196.480 ;
    END
  END Tile_X0Y1_FrameData_O[17]
  PIN Tile_X0Y1_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 197.240 199.640 197.840 ;
    END
  END Tile_X0Y1_FrameData_O[18]
  PIN Tile_X0Y1_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 198.600 199.640 199.200 ;
    END
  END Tile_X0Y1_FrameData_O[19]
  PIN Tile_X0Y1_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 174.120 199.640 174.720 ;
    END
  END Tile_X0Y1_FrameData_O[1]
  PIN Tile_X0Y1_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 199.960 199.640 200.560 ;
    END
  END Tile_X0Y1_FrameData_O[20]
  PIN Tile_X0Y1_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 201.320 199.640 201.920 ;
    END
  END Tile_X0Y1_FrameData_O[21]
  PIN Tile_X0Y1_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 202.680 199.640 203.280 ;
    END
  END Tile_X0Y1_FrameData_O[22]
  PIN Tile_X0Y1_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 204.040 199.640 204.640 ;
    END
  END Tile_X0Y1_FrameData_O[23]
  PIN Tile_X0Y1_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 205.400 199.640 206.000 ;
    END
  END Tile_X0Y1_FrameData_O[24]
  PIN Tile_X0Y1_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 206.760 199.640 207.360 ;
    END
  END Tile_X0Y1_FrameData_O[25]
  PIN Tile_X0Y1_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 208.120 199.640 208.720 ;
    END
  END Tile_X0Y1_FrameData_O[26]
  PIN Tile_X0Y1_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 209.480 199.640 210.080 ;
    END
  END Tile_X0Y1_FrameData_O[27]
  PIN Tile_X0Y1_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 210.840 199.640 211.440 ;
    END
  END Tile_X0Y1_FrameData_O[28]
  PIN Tile_X0Y1_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 212.200 199.640 212.800 ;
    END
  END Tile_X0Y1_FrameData_O[29]
  PIN Tile_X0Y1_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 175.480 199.640 176.080 ;
    END
  END Tile_X0Y1_FrameData_O[2]
  PIN Tile_X0Y1_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 213.560 199.640 214.160 ;
    END
  END Tile_X0Y1_FrameData_O[30]
  PIN Tile_X0Y1_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 214.920 199.640 215.520 ;
    END
  END Tile_X0Y1_FrameData_O[31]
  PIN Tile_X0Y1_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 176.840 199.640 177.440 ;
    END
  END Tile_X0Y1_FrameData_O[3]
  PIN Tile_X0Y1_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 178.200 199.640 178.800 ;
    END
  END Tile_X0Y1_FrameData_O[4]
  PIN Tile_X0Y1_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 179.560 199.640 180.160 ;
    END
  END Tile_X0Y1_FrameData_O[5]
  PIN Tile_X0Y1_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 180.920 199.640 181.520 ;
    END
  END Tile_X0Y1_FrameData_O[6]
  PIN Tile_X0Y1_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 182.280 199.640 182.880 ;
    END
  END Tile_X0Y1_FrameData_O[7]
  PIN Tile_X0Y1_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 183.640 199.640 184.240 ;
    END
  END Tile_X0Y1_FrameData_O[8]
  PIN Tile_X0Y1_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 185.000 199.640 185.600 ;
    END
  END Tile_X0Y1_FrameData_O[9]
  PIN Tile_X0Y1_FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.372000 ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[0]
  PIN Tile_X0Y1_FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[10]
  PIN Tile_X0Y1_FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[11]
  PIN Tile_X0Y1_FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[12]
  PIN Tile_X0Y1_FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[13]
  PIN Tile_X0Y1_FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[14]
  PIN Tile_X0Y1_FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[15]
  PIN Tile_X0Y1_FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[16]
  PIN Tile_X0Y1_FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[17]
  PIN Tile_X0Y1_FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[18]
  PIN Tile_X0Y1_FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[19]
  PIN Tile_X0Y1_FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[1]
  PIN Tile_X0Y1_FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[2]
  PIN Tile_X0Y1_FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[3]
  PIN Tile_X0Y1_FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[4]
  PIN Tile_X0Y1_FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[5]
  PIN Tile_X0Y1_FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639000 ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[6]
  PIN Tile_X0Y1_FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.552000 ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[7]
  PIN Tile_X0Y1_FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[8]
  PIN Tile_X0Y1_FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 0.280 ;
    END
  END Tile_X0Y1_FrameStrobe[9]
  PIN Tile_X0Y1_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 0.280 ;
    END
  END Tile_X0Y1_N1END[0]
  PIN Tile_X0Y1_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 0.280 ;
    END
  END Tile_X0Y1_N1END[1]
  PIN Tile_X0Y1_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 0.280 ;
    END
  END Tile_X0Y1_N1END[2]
  PIN Tile_X0Y1_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 0.280 ;
    END
  END Tile_X0Y1_N1END[3]
  PIN Tile_X0Y1_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 0.280 ;
    END
  END Tile_X0Y1_N2END[0]
  PIN Tile_X0Y1_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 0.280 ;
    END
  END Tile_X0Y1_N2END[1]
  PIN Tile_X0Y1_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 0.280 ;
    END
  END Tile_X0Y1_N2END[2]
  PIN Tile_X0Y1_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 0.280 ;
    END
  END Tile_X0Y1_N2END[3]
  PIN Tile_X0Y1_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 0.280 ;
    END
  END Tile_X0Y1_N2END[4]
  PIN Tile_X0Y1_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 0.280 ;
    END
  END Tile_X0Y1_N2END[5]
  PIN Tile_X0Y1_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 0.280 ;
    END
  END Tile_X0Y1_N2END[6]
  PIN Tile_X0Y1_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 0.280 ;
    END
  END Tile_X0Y1_N2END[7]
  PIN Tile_X0Y1_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 0.280 ;
    END
  END Tile_X0Y1_N2MID[0]
  PIN Tile_X0Y1_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 0.280 ;
    END
  END Tile_X0Y1_N2MID[1]
  PIN Tile_X0Y1_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 0.280 ;
    END
  END Tile_X0Y1_N2MID[2]
  PIN Tile_X0Y1_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 0.280 ;
    END
  END Tile_X0Y1_N2MID[3]
  PIN Tile_X0Y1_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 0.280 ;
    END
  END Tile_X0Y1_N2MID[4]
  PIN Tile_X0Y1_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 0.280 ;
    END
  END Tile_X0Y1_N2MID[5]
  PIN Tile_X0Y1_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 0.280 ;
    END
  END Tile_X0Y1_N2MID[6]
  PIN Tile_X0Y1_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 0.280 ;
    END
  END Tile_X0Y1_N2MID[7]
  PIN Tile_X0Y1_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 0.280 ;
    END
  END Tile_X0Y1_N4END[0]
  PIN Tile_X0Y1_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 0.280 ;
    END
  END Tile_X0Y1_N4END[10]
  PIN Tile_X0Y1_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 0.280 ;
    END
  END Tile_X0Y1_N4END[11]
  PIN Tile_X0Y1_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 0.280 ;
    END
  END Tile_X0Y1_N4END[12]
  PIN Tile_X0Y1_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 0.280 ;
    END
  END Tile_X0Y1_N4END[13]
  PIN Tile_X0Y1_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 0.280 ;
    END
  END Tile_X0Y1_N4END[14]
  PIN Tile_X0Y1_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 0.280 ;
    END
  END Tile_X0Y1_N4END[15]
  PIN Tile_X0Y1_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 0.280 ;
    END
  END Tile_X0Y1_N4END[1]
  PIN Tile_X0Y1_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 0.280 ;
    END
  END Tile_X0Y1_N4END[2]
  PIN Tile_X0Y1_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 0.280 ;
    END
  END Tile_X0Y1_N4END[3]
  PIN Tile_X0Y1_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 0.280 ;
    END
  END Tile_X0Y1_N4END[4]
  PIN Tile_X0Y1_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 0.280 ;
    END
  END Tile_X0Y1_N4END[5]
  PIN Tile_X0Y1_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 0.280 ;
    END
  END Tile_X0Y1_N4END[6]
  PIN Tile_X0Y1_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 0.280 ;
    END
  END Tile_X0Y1_N4END[7]
  PIN Tile_X0Y1_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 0.280 ;
    END
  END Tile_X0Y1_N4END[8]
  PIN Tile_X0Y1_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 0.280 ;
    END
  END Tile_X0Y1_N4END[9]
  PIN Tile_X0Y1_NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 0.280 ;
    END
  END Tile_X0Y1_NN4END[0]
  PIN Tile_X0Y1_NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 0.280 ;
    END
  END Tile_X0Y1_NN4END[10]
  PIN Tile_X0Y1_NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 0.280 ;
    END
  END Tile_X0Y1_NN4END[11]
  PIN Tile_X0Y1_NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 0.280 ;
    END
  END Tile_X0Y1_NN4END[12]
  PIN Tile_X0Y1_NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 0.280 ;
    END
  END Tile_X0Y1_NN4END[13]
  PIN Tile_X0Y1_NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 0.280 ;
    END
  END Tile_X0Y1_NN4END[14]
  PIN Tile_X0Y1_NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 0.280 ;
    END
  END Tile_X0Y1_NN4END[15]
  PIN Tile_X0Y1_NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 0.280 ;
    END
  END Tile_X0Y1_NN4END[1]
  PIN Tile_X0Y1_NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 0.280 ;
    END
  END Tile_X0Y1_NN4END[2]
  PIN Tile_X0Y1_NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 0.280 ;
    END
  END Tile_X0Y1_NN4END[3]
  PIN Tile_X0Y1_NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 0.280 ;
    END
  END Tile_X0Y1_NN4END[4]
  PIN Tile_X0Y1_NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 0.280 ;
    END
  END Tile_X0Y1_NN4END[5]
  PIN Tile_X0Y1_NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 0.280 ;
    END
  END Tile_X0Y1_NN4END[6]
  PIN Tile_X0Y1_NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 0.280 ;
    END
  END Tile_X0Y1_NN4END[7]
  PIN Tile_X0Y1_NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 0.280 ;
    END
  END Tile_X0Y1_NN4END[8]
  PIN Tile_X0Y1_NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 0.280 ;
    END
  END Tile_X0Y1_NN4END[9]
  PIN Tile_X0Y1_S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 0.280 ;
    END
  END Tile_X0Y1_S1BEG[0]
  PIN Tile_X0Y1_S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 0.280 ;
    END
  END Tile_X0Y1_S1BEG[1]
  PIN Tile_X0Y1_S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 0.280 ;
    END
  END Tile_X0Y1_S1BEG[2]
  PIN Tile_X0Y1_S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 0.280 ;
    END
  END Tile_X0Y1_S1BEG[3]
  PIN Tile_X0Y1_S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 0.280 ;
    END
  END Tile_X0Y1_S2BEG[0]
  PIN Tile_X0Y1_S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 0.280 ;
    END
  END Tile_X0Y1_S2BEG[1]
  PIN Tile_X0Y1_S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 0.280 ;
    END
  END Tile_X0Y1_S2BEG[2]
  PIN Tile_X0Y1_S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 0.280 ;
    END
  END Tile_X0Y1_S2BEG[3]
  PIN Tile_X0Y1_S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 0.280 ;
    END
  END Tile_X0Y1_S2BEG[4]
  PIN Tile_X0Y1_S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 0.280 ;
    END
  END Tile_X0Y1_S2BEG[5]
  PIN Tile_X0Y1_S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 0.280 ;
    END
  END Tile_X0Y1_S2BEG[6]
  PIN Tile_X0Y1_S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 0.280 ;
    END
  END Tile_X0Y1_S2BEG[7]
  PIN Tile_X0Y1_S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[0]
  PIN Tile_X0Y1_S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[1]
  PIN Tile_X0Y1_S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[2]
  PIN Tile_X0Y1_S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[3]
  PIN Tile_X0Y1_S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[4]
  PIN Tile_X0Y1_S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[5]
  PIN Tile_X0Y1_S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[6]
  PIN Tile_X0Y1_S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 0.280 ;
    END
  END Tile_X0Y1_S2BEGb[7]
  PIN Tile_X0Y1_S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 0.280 ;
    END
  END Tile_X0Y1_S4BEG[0]
  PIN Tile_X0Y1_S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 0.280 ;
    END
  END Tile_X0Y1_S4BEG[10]
  PIN Tile_X0Y1_S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 0.280 ;
    END
  END Tile_X0Y1_S4BEG[11]
  PIN Tile_X0Y1_S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 0.280 ;
    END
  END Tile_X0Y1_S4BEG[12]
  PIN Tile_X0Y1_S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 0.280 ;
    END
  END Tile_X0Y1_S4BEG[13]
  PIN Tile_X0Y1_S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 0.280 ;
    END
  END Tile_X0Y1_S4BEG[14]
  PIN Tile_X0Y1_S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 0.280 ;
    END
  END Tile_X0Y1_S4BEG[15]
  PIN Tile_X0Y1_S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 0.280 ;
    END
  END Tile_X0Y1_S4BEG[1]
  PIN Tile_X0Y1_S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 0.280 ;
    END
  END Tile_X0Y1_S4BEG[2]
  PIN Tile_X0Y1_S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 0.280 ;
    END
  END Tile_X0Y1_S4BEG[3]
  PIN Tile_X0Y1_S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 0.280 ;
    END
  END Tile_X0Y1_S4BEG[4]
  PIN Tile_X0Y1_S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 0.280 ;
    END
  END Tile_X0Y1_S4BEG[5]
  PIN Tile_X0Y1_S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 0.280 ;
    END
  END Tile_X0Y1_S4BEG[6]
  PIN Tile_X0Y1_S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 0.280 ;
    END
  END Tile_X0Y1_S4BEG[7]
  PIN Tile_X0Y1_S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 0.280 ;
    END
  END Tile_X0Y1_S4BEG[8]
  PIN Tile_X0Y1_S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 0.280 ;
    END
  END Tile_X0Y1_S4BEG[9]
  PIN Tile_X0Y1_SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[0]
  PIN Tile_X0Y1_SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[10]
  PIN Tile_X0Y1_SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[11]
  PIN Tile_X0Y1_SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[12]
  PIN Tile_X0Y1_SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[13]
  PIN Tile_X0Y1_SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[14]
  PIN Tile_X0Y1_SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[15]
  PIN Tile_X0Y1_SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[1]
  PIN Tile_X0Y1_SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[2]
  PIN Tile_X0Y1_SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[3]
  PIN Tile_X0Y1_SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[4]
  PIN Tile_X0Y1_SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[5]
  PIN Tile_X0Y1_SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[6]
  PIN Tile_X0Y1_SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[7]
  PIN Tile_X0Y1_SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[8]
  PIN Tile_X0Y1_SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 0.280 ;
    END
  END Tile_X0Y1_SS4BEG[9]
  PIN Tile_X0Y1_UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.704000 ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 0.280 ;
    END
  END Tile_X0Y1_UserCLK
  PIN Tile_X0Y1_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 0.600 42.800 ;
    END
  END Tile_X0Y1_W1BEG[0]
  PIN Tile_X0Y1_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 0.600 44.160 ;
    END
  END Tile_X0Y1_W1BEG[1]
  PIN Tile_X0Y1_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 0.600 45.520 ;
    END
  END Tile_X0Y1_W1BEG[2]
  PIN Tile_X0Y1_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 0.600 46.880 ;
    END
  END Tile_X0Y1_W1BEG[3]
  PIN Tile_X0Y1_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 42.200 199.640 42.800 ;
    END
  END Tile_X0Y1_W1END[0]
  PIN Tile_X0Y1_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 43.560 199.640 44.160 ;
    END
  END Tile_X0Y1_W1END[1]
  PIN Tile_X0Y1_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 44.920 199.640 45.520 ;
    END
  END Tile_X0Y1_W1END[2]
  PIN Tile_X0Y1_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 199.040 46.280 199.640 46.880 ;
    END
  END Tile_X0Y1_W1END[3]
  PIN Tile_X0Y1_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 0.600 48.240 ;
    END
  END Tile_X0Y1_W2BEG[0]
  PIN Tile_X0Y1_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 0.600 49.600 ;
    END
  END Tile_X0Y1_W2BEG[1]
  PIN Tile_X0Y1_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 0.600 50.960 ;
    END
  END Tile_X0Y1_W2BEG[2]
  PIN Tile_X0Y1_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 0.600 52.320 ;
    END
  END Tile_X0Y1_W2BEG[3]
  PIN Tile_X0Y1_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 0.600 53.680 ;
    END
  END Tile_X0Y1_W2BEG[4]
  PIN Tile_X0Y1_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 0.600 55.040 ;
    END
  END Tile_X0Y1_W2BEG[5]
  PIN Tile_X0Y1_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 0.600 56.400 ;
    END
  END Tile_X0Y1_W2BEG[6]
  PIN Tile_X0Y1_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 0.600 57.760 ;
    END
  END Tile_X0Y1_W2BEG[7]
  PIN Tile_X0Y1_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 0.600 59.120 ;
    END
  END Tile_X0Y1_W2BEGb[0]
  PIN Tile_X0Y1_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 0.600 60.480 ;
    END
  END Tile_X0Y1_W2BEGb[1]
  PIN Tile_X0Y1_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 0.600 61.840 ;
    END
  END Tile_X0Y1_W2BEGb[2]
  PIN Tile_X0Y1_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 0.600 63.200 ;
    END
  END Tile_X0Y1_W2BEGb[3]
  PIN Tile_X0Y1_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 0.600 64.560 ;
    END
  END Tile_X0Y1_W2BEGb[4]
  PIN Tile_X0Y1_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 0.600 65.920 ;
    END
  END Tile_X0Y1_W2BEGb[5]
  PIN Tile_X0Y1_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 0.600 67.280 ;
    END
  END Tile_X0Y1_W2BEGb[6]
  PIN Tile_X0Y1_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 0.600 68.640 ;
    END
  END Tile_X0Y1_W2BEGb[7]
  PIN Tile_X0Y1_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 58.520 199.640 59.120 ;
    END
  END Tile_X0Y1_W2END[0]
  PIN Tile_X0Y1_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 59.880 199.640 60.480 ;
    END
  END Tile_X0Y1_W2END[1]
  PIN Tile_X0Y1_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 61.240 199.640 61.840 ;
    END
  END Tile_X0Y1_W2END[2]
  PIN Tile_X0Y1_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 62.600 199.640 63.200 ;
    END
  END Tile_X0Y1_W2END[3]
  PIN Tile_X0Y1_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 63.960 199.640 64.560 ;
    END
  END Tile_X0Y1_W2END[4]
  PIN Tile_X0Y1_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 65.320 199.640 65.920 ;
    END
  END Tile_X0Y1_W2END[5]
  PIN Tile_X0Y1_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 66.680 199.640 67.280 ;
    END
  END Tile_X0Y1_W2END[6]
  PIN Tile_X0Y1_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 68.040 199.640 68.640 ;
    END
  END Tile_X0Y1_W2END[7]
  PIN Tile_X0Y1_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 47.640 199.640 48.240 ;
    END
  END Tile_X0Y1_W2MID[0]
  PIN Tile_X0Y1_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 49.000 199.640 49.600 ;
    END
  END Tile_X0Y1_W2MID[1]
  PIN Tile_X0Y1_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 50.360 199.640 50.960 ;
    END
  END Tile_X0Y1_W2MID[2]
  PIN Tile_X0Y1_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 51.720 199.640 52.320 ;
    END
  END Tile_X0Y1_W2MID[3]
  PIN Tile_X0Y1_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 53.080 199.640 53.680 ;
    END
  END Tile_X0Y1_W2MID[4]
  PIN Tile_X0Y1_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 54.440 199.640 55.040 ;
    END
  END Tile_X0Y1_W2MID[5]
  PIN Tile_X0Y1_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 55.800 199.640 56.400 ;
    END
  END Tile_X0Y1_W2MID[6]
  PIN Tile_X0Y1_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 57.160 199.640 57.760 ;
    END
  END Tile_X0Y1_W2MID[7]
  PIN Tile_X0Y1_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 0.600 91.760 ;
    END
  END Tile_X0Y1_W6BEG[0]
  PIN Tile_X0Y1_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 0.600 105.360 ;
    END
  END Tile_X0Y1_W6BEG[10]
  PIN Tile_X0Y1_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 0.600 106.720 ;
    END
  END Tile_X0Y1_W6BEG[11]
  PIN Tile_X0Y1_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 0.600 93.120 ;
    END
  END Tile_X0Y1_W6BEG[1]
  PIN Tile_X0Y1_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 0.600 94.480 ;
    END
  END Tile_X0Y1_W6BEG[2]
  PIN Tile_X0Y1_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 0.600 95.840 ;
    END
  END Tile_X0Y1_W6BEG[3]
  PIN Tile_X0Y1_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 0.600 97.200 ;
    END
  END Tile_X0Y1_W6BEG[4]
  PIN Tile_X0Y1_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 0.600 98.560 ;
    END
  END Tile_X0Y1_W6BEG[5]
  PIN Tile_X0Y1_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 0.600 99.920 ;
    END
  END Tile_X0Y1_W6BEG[6]
  PIN Tile_X0Y1_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 0.600 101.280 ;
    END
  END Tile_X0Y1_W6BEG[7]
  PIN Tile_X0Y1_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 0.600 102.640 ;
    END
  END Tile_X0Y1_W6BEG[8]
  PIN Tile_X0Y1_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 0.600 104.000 ;
    END
  END Tile_X0Y1_W6BEG[9]
  PIN Tile_X0Y1_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 91.160 199.640 91.760 ;
    END
  END Tile_X0Y1_W6END[0]
  PIN Tile_X0Y1_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 104.760 199.640 105.360 ;
    END
  END Tile_X0Y1_W6END[10]
  PIN Tile_X0Y1_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 106.120 199.640 106.720 ;
    END
  END Tile_X0Y1_W6END[11]
  PIN Tile_X0Y1_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 92.520 199.640 93.120 ;
    END
  END Tile_X0Y1_W6END[1]
  PIN Tile_X0Y1_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 93.880 199.640 94.480 ;
    END
  END Tile_X0Y1_W6END[2]
  PIN Tile_X0Y1_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 95.240 199.640 95.840 ;
    END
  END Tile_X0Y1_W6END[3]
  PIN Tile_X0Y1_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 96.600 199.640 97.200 ;
    END
  END Tile_X0Y1_W6END[4]
  PIN Tile_X0Y1_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 97.960 199.640 98.560 ;
    END
  END Tile_X0Y1_W6END[5]
  PIN Tile_X0Y1_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 99.320 199.640 99.920 ;
    END
  END Tile_X0Y1_W6END[6]
  PIN Tile_X0Y1_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 100.680 199.640 101.280 ;
    END
  END Tile_X0Y1_W6END[7]
  PIN Tile_X0Y1_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 102.040 199.640 102.640 ;
    END
  END Tile_X0Y1_W6END[8]
  PIN Tile_X0Y1_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 103.400 199.640 104.000 ;
    END
  END Tile_X0Y1_W6END[9]
  PIN Tile_X0Y1_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 0.600 70.000 ;
    END
  END Tile_X0Y1_WW4BEG[0]
  PIN Tile_X0Y1_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 0.600 83.600 ;
    END
  END Tile_X0Y1_WW4BEG[10]
  PIN Tile_X0Y1_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 0.600 84.960 ;
    END
  END Tile_X0Y1_WW4BEG[11]
  PIN Tile_X0Y1_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 0.600 86.320 ;
    END
  END Tile_X0Y1_WW4BEG[12]
  PIN Tile_X0Y1_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 0.600 87.680 ;
    END
  END Tile_X0Y1_WW4BEG[13]
  PIN Tile_X0Y1_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 0.600 89.040 ;
    END
  END Tile_X0Y1_WW4BEG[14]
  PIN Tile_X0Y1_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 0.600 90.400 ;
    END
  END Tile_X0Y1_WW4BEG[15]
  PIN Tile_X0Y1_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 0.600 71.360 ;
    END
  END Tile_X0Y1_WW4BEG[1]
  PIN Tile_X0Y1_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 0.600 72.720 ;
    END
  END Tile_X0Y1_WW4BEG[2]
  PIN Tile_X0Y1_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 0.600 74.080 ;
    END
  END Tile_X0Y1_WW4BEG[3]
  PIN Tile_X0Y1_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 0.600 75.440 ;
    END
  END Tile_X0Y1_WW4BEG[4]
  PIN Tile_X0Y1_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 0.600 76.800 ;
    END
  END Tile_X0Y1_WW4BEG[5]
  PIN Tile_X0Y1_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 0.600 78.160 ;
    END
  END Tile_X0Y1_WW4BEG[6]
  PIN Tile_X0Y1_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 0.600 79.520 ;
    END
  END Tile_X0Y1_WW4BEG[7]
  PIN Tile_X0Y1_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 0.600 80.880 ;
    END
  END Tile_X0Y1_WW4BEG[8]
  PIN Tile_X0Y1_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 0.600 82.240 ;
    END
  END Tile_X0Y1_WW4BEG[9]
  PIN Tile_X0Y1_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 69.400 199.640 70.000 ;
    END
  END Tile_X0Y1_WW4END[0]
  PIN Tile_X0Y1_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 83.000 199.640 83.600 ;
    END
  END Tile_X0Y1_WW4END[10]
  PIN Tile_X0Y1_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 84.360 199.640 84.960 ;
    END
  END Tile_X0Y1_WW4END[11]
  PIN Tile_X0Y1_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 85.720 199.640 86.320 ;
    END
  END Tile_X0Y1_WW4END[12]
  PIN Tile_X0Y1_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 87.080 199.640 87.680 ;
    END
  END Tile_X0Y1_WW4END[13]
  PIN Tile_X0Y1_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 88.440 199.640 89.040 ;
    END
  END Tile_X0Y1_WW4END[14]
  PIN Tile_X0Y1_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 89.800 199.640 90.400 ;
    END
  END Tile_X0Y1_WW4END[15]
  PIN Tile_X0Y1_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 70.760 199.640 71.360 ;
    END
  END Tile_X0Y1_WW4END[1]
  PIN Tile_X0Y1_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 72.120 199.640 72.720 ;
    END
  END Tile_X0Y1_WW4END[2]
  PIN Tile_X0Y1_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 73.480 199.640 74.080 ;
    END
  END Tile_X0Y1_WW4END[3]
  PIN Tile_X0Y1_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 74.840 199.640 75.440 ;
    END
  END Tile_X0Y1_WW4END[4]
  PIN Tile_X0Y1_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 76.200 199.640 76.800 ;
    END
  END Tile_X0Y1_WW4END[5]
  PIN Tile_X0Y1_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 77.560 199.640 78.160 ;
    END
  END Tile_X0Y1_WW4END[6]
  PIN Tile_X0Y1_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 78.920 199.640 79.520 ;
    END
  END Tile_X0Y1_WW4END[7]
  PIN Tile_X0Y1_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 80.280 199.640 80.880 ;
    END
  END Tile_X0Y1_WW4END[8]
  PIN Tile_X0Y1_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 199.040 81.640 199.640 82.240 ;
    END
  END Tile_X0Y1_WW4END[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.020 0.000 16.620 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.020 0.000 46.620 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.020 0.000 76.620 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.020 0.000 106.620 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.020 0.000 136.620 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 165.020 0.000 166.620 519.520 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 0.000 11.320 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.720 0.000 41.320 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.720 0.000 71.320 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.720 0.000 101.320 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 129.720 0.000 131.320 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.720 0.000 161.320 519.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.720 0.000 191.320 519.520 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 194.310 508.830 ;
      LAYER li1 ;
        RECT 5.520 10.795 194.120 508.725 ;
      LAYER met1 ;
        RECT 0.070 0.040 199.570 519.480 ;
      LAYER met2 ;
        RECT 0.100 518.960 13.610 519.510 ;
        RECT 14.450 518.960 14.990 519.510 ;
        RECT 15.830 518.960 16.370 519.510 ;
        RECT 17.210 518.960 17.750 519.510 ;
        RECT 18.590 518.960 19.130 519.510 ;
        RECT 19.970 518.960 20.510 519.510 ;
        RECT 21.350 518.960 21.890 519.510 ;
        RECT 22.730 518.960 23.270 519.510 ;
        RECT 24.110 518.960 24.650 519.510 ;
        RECT 25.490 518.960 26.030 519.510 ;
        RECT 26.870 518.960 27.410 519.510 ;
        RECT 28.250 518.960 28.790 519.510 ;
        RECT 29.630 518.960 30.170 519.510 ;
        RECT 31.010 518.960 31.550 519.510 ;
        RECT 32.390 518.960 32.930 519.510 ;
        RECT 33.770 518.960 34.310 519.510 ;
        RECT 35.150 518.960 35.690 519.510 ;
        RECT 36.530 518.960 37.070 519.510 ;
        RECT 37.910 518.960 38.450 519.510 ;
        RECT 39.290 518.960 39.830 519.510 ;
        RECT 40.670 518.960 41.210 519.510 ;
        RECT 42.050 518.960 42.590 519.510 ;
        RECT 43.430 518.960 43.970 519.510 ;
        RECT 44.810 518.960 45.350 519.510 ;
        RECT 46.190 518.960 46.730 519.510 ;
        RECT 47.570 518.960 48.110 519.510 ;
        RECT 48.950 518.960 49.490 519.510 ;
        RECT 50.330 518.960 50.870 519.510 ;
        RECT 51.710 518.960 52.250 519.510 ;
        RECT 53.090 518.960 53.630 519.510 ;
        RECT 54.470 518.960 55.010 519.510 ;
        RECT 55.850 518.960 56.390 519.510 ;
        RECT 57.230 518.960 57.770 519.510 ;
        RECT 58.610 518.960 59.150 519.510 ;
        RECT 59.990 518.960 60.530 519.510 ;
        RECT 61.370 518.960 61.910 519.510 ;
        RECT 62.750 518.960 63.290 519.510 ;
        RECT 64.130 518.960 64.670 519.510 ;
        RECT 65.510 518.960 66.050 519.510 ;
        RECT 66.890 518.960 67.430 519.510 ;
        RECT 68.270 518.960 68.810 519.510 ;
        RECT 69.650 518.960 70.190 519.510 ;
        RECT 71.030 518.960 71.570 519.510 ;
        RECT 72.410 518.960 72.950 519.510 ;
        RECT 73.790 518.960 74.330 519.510 ;
        RECT 75.170 518.960 75.710 519.510 ;
        RECT 76.550 518.960 77.090 519.510 ;
        RECT 77.930 518.960 78.470 519.510 ;
        RECT 79.310 518.960 79.850 519.510 ;
        RECT 80.690 518.960 81.230 519.510 ;
        RECT 82.070 518.960 82.610 519.510 ;
        RECT 83.450 518.960 83.990 519.510 ;
        RECT 84.830 518.960 85.370 519.510 ;
        RECT 86.210 518.960 86.750 519.510 ;
        RECT 87.590 518.960 88.130 519.510 ;
        RECT 88.970 518.960 89.510 519.510 ;
        RECT 90.350 518.960 90.890 519.510 ;
        RECT 91.730 518.960 92.270 519.510 ;
        RECT 93.110 518.960 93.650 519.510 ;
        RECT 94.490 518.960 95.030 519.510 ;
        RECT 95.870 518.960 96.410 519.510 ;
        RECT 97.250 518.960 97.790 519.510 ;
        RECT 98.630 518.960 99.170 519.510 ;
        RECT 100.010 518.960 100.550 519.510 ;
        RECT 101.390 518.960 101.930 519.510 ;
        RECT 102.770 518.960 103.310 519.510 ;
        RECT 104.150 518.960 104.690 519.510 ;
        RECT 105.530 518.960 106.070 519.510 ;
        RECT 106.910 518.960 107.450 519.510 ;
        RECT 108.290 518.960 108.830 519.510 ;
        RECT 109.670 518.960 110.210 519.510 ;
        RECT 111.050 518.960 111.590 519.510 ;
        RECT 112.430 518.960 112.970 519.510 ;
        RECT 113.810 518.960 114.350 519.510 ;
        RECT 115.190 518.960 115.730 519.510 ;
        RECT 116.570 518.960 117.110 519.510 ;
        RECT 117.950 518.960 118.490 519.510 ;
        RECT 119.330 518.960 119.870 519.510 ;
        RECT 120.710 518.960 121.250 519.510 ;
        RECT 122.090 518.960 122.630 519.510 ;
        RECT 123.470 518.960 124.010 519.510 ;
        RECT 124.850 518.960 125.390 519.510 ;
        RECT 126.230 518.960 126.770 519.510 ;
        RECT 127.610 518.960 128.150 519.510 ;
        RECT 128.990 518.960 129.530 519.510 ;
        RECT 130.370 518.960 130.910 519.510 ;
        RECT 131.750 518.960 132.290 519.510 ;
        RECT 133.130 518.960 133.670 519.510 ;
        RECT 134.510 518.960 135.050 519.510 ;
        RECT 135.890 518.960 136.430 519.510 ;
        RECT 137.270 518.960 137.810 519.510 ;
        RECT 138.650 518.960 139.190 519.510 ;
        RECT 140.030 518.960 140.570 519.510 ;
        RECT 141.410 518.960 141.950 519.510 ;
        RECT 142.790 518.960 143.330 519.510 ;
        RECT 144.170 518.960 144.710 519.510 ;
        RECT 145.550 518.960 146.090 519.510 ;
        RECT 146.930 518.960 147.470 519.510 ;
        RECT 148.310 518.960 148.850 519.510 ;
        RECT 149.690 518.960 150.230 519.510 ;
        RECT 151.070 518.960 151.610 519.510 ;
        RECT 152.450 518.960 152.990 519.510 ;
        RECT 153.830 518.960 154.370 519.510 ;
        RECT 155.210 518.960 155.750 519.510 ;
        RECT 156.590 518.960 157.130 519.510 ;
        RECT 157.970 518.960 158.510 519.510 ;
        RECT 159.350 518.960 159.890 519.510 ;
        RECT 160.730 518.960 161.270 519.510 ;
        RECT 162.110 518.960 162.650 519.510 ;
        RECT 163.490 518.960 164.030 519.510 ;
        RECT 164.870 518.960 165.410 519.510 ;
        RECT 166.250 518.960 166.790 519.510 ;
        RECT 167.630 518.960 168.170 519.510 ;
        RECT 169.010 518.960 169.550 519.510 ;
        RECT 170.390 518.960 170.930 519.510 ;
        RECT 171.770 518.960 172.310 519.510 ;
        RECT 173.150 518.960 173.690 519.510 ;
        RECT 174.530 518.960 175.070 519.510 ;
        RECT 175.910 518.960 176.450 519.510 ;
        RECT 177.290 518.960 177.830 519.510 ;
        RECT 178.670 518.960 179.210 519.510 ;
        RECT 180.050 518.960 180.590 519.510 ;
        RECT 181.430 518.960 181.970 519.510 ;
        RECT 182.810 518.960 183.350 519.510 ;
        RECT 184.190 518.960 184.730 519.510 ;
        RECT 185.570 518.960 199.540 519.510 ;
        RECT 0.100 0.560 199.540 518.960 ;
        RECT 0.100 0.010 13.610 0.560 ;
        RECT 14.450 0.010 14.990 0.560 ;
        RECT 15.830 0.010 16.370 0.560 ;
        RECT 17.210 0.010 17.750 0.560 ;
        RECT 18.590 0.010 19.130 0.560 ;
        RECT 19.970 0.010 20.510 0.560 ;
        RECT 21.350 0.010 21.890 0.560 ;
        RECT 22.730 0.010 23.270 0.560 ;
        RECT 24.110 0.010 24.650 0.560 ;
        RECT 25.490 0.010 26.030 0.560 ;
        RECT 26.870 0.010 27.410 0.560 ;
        RECT 28.250 0.010 28.790 0.560 ;
        RECT 29.630 0.010 30.170 0.560 ;
        RECT 31.010 0.010 31.550 0.560 ;
        RECT 32.390 0.010 32.930 0.560 ;
        RECT 33.770 0.010 34.310 0.560 ;
        RECT 35.150 0.010 35.690 0.560 ;
        RECT 36.530 0.010 37.070 0.560 ;
        RECT 37.910 0.010 38.450 0.560 ;
        RECT 39.290 0.010 39.830 0.560 ;
        RECT 40.670 0.010 41.210 0.560 ;
        RECT 42.050 0.010 42.590 0.560 ;
        RECT 43.430 0.010 43.970 0.560 ;
        RECT 44.810 0.010 45.350 0.560 ;
        RECT 46.190 0.010 46.730 0.560 ;
        RECT 47.570 0.010 48.110 0.560 ;
        RECT 48.950 0.010 49.490 0.560 ;
        RECT 50.330 0.010 50.870 0.560 ;
        RECT 51.710 0.010 52.250 0.560 ;
        RECT 53.090 0.010 53.630 0.560 ;
        RECT 54.470 0.010 55.010 0.560 ;
        RECT 55.850 0.010 56.390 0.560 ;
        RECT 57.230 0.010 57.770 0.560 ;
        RECT 58.610 0.010 59.150 0.560 ;
        RECT 59.990 0.010 60.530 0.560 ;
        RECT 61.370 0.010 61.910 0.560 ;
        RECT 62.750 0.010 63.290 0.560 ;
        RECT 64.130 0.010 64.670 0.560 ;
        RECT 65.510 0.010 66.050 0.560 ;
        RECT 66.890 0.010 67.430 0.560 ;
        RECT 68.270 0.010 68.810 0.560 ;
        RECT 69.650 0.010 70.190 0.560 ;
        RECT 71.030 0.010 71.570 0.560 ;
        RECT 72.410 0.010 72.950 0.560 ;
        RECT 73.790 0.010 74.330 0.560 ;
        RECT 75.170 0.010 75.710 0.560 ;
        RECT 76.550 0.010 77.090 0.560 ;
        RECT 77.930 0.010 78.470 0.560 ;
        RECT 79.310 0.010 79.850 0.560 ;
        RECT 80.690 0.010 81.230 0.560 ;
        RECT 82.070 0.010 82.610 0.560 ;
        RECT 83.450 0.010 83.990 0.560 ;
        RECT 84.830 0.010 85.370 0.560 ;
        RECT 86.210 0.010 86.750 0.560 ;
        RECT 87.590 0.010 88.130 0.560 ;
        RECT 88.970 0.010 89.510 0.560 ;
        RECT 90.350 0.010 90.890 0.560 ;
        RECT 91.730 0.010 92.270 0.560 ;
        RECT 93.110 0.010 93.650 0.560 ;
        RECT 94.490 0.010 95.030 0.560 ;
        RECT 95.870 0.010 96.410 0.560 ;
        RECT 97.250 0.010 97.790 0.560 ;
        RECT 98.630 0.010 99.170 0.560 ;
        RECT 100.010 0.010 100.550 0.560 ;
        RECT 101.390 0.010 101.930 0.560 ;
        RECT 102.770 0.010 103.310 0.560 ;
        RECT 104.150 0.010 104.690 0.560 ;
        RECT 105.530 0.010 106.070 0.560 ;
        RECT 106.910 0.010 107.450 0.560 ;
        RECT 108.290 0.010 108.830 0.560 ;
        RECT 109.670 0.010 110.210 0.560 ;
        RECT 111.050 0.010 111.590 0.560 ;
        RECT 112.430 0.010 112.970 0.560 ;
        RECT 113.810 0.010 114.350 0.560 ;
        RECT 115.190 0.010 115.730 0.560 ;
        RECT 116.570 0.010 117.110 0.560 ;
        RECT 117.950 0.010 118.490 0.560 ;
        RECT 119.330 0.010 119.870 0.560 ;
        RECT 120.710 0.010 121.250 0.560 ;
        RECT 122.090 0.010 122.630 0.560 ;
        RECT 123.470 0.010 124.010 0.560 ;
        RECT 124.850 0.010 125.390 0.560 ;
        RECT 126.230 0.010 126.770 0.560 ;
        RECT 127.610 0.010 128.150 0.560 ;
        RECT 128.990 0.010 129.530 0.560 ;
        RECT 130.370 0.010 130.910 0.560 ;
        RECT 131.750 0.010 132.290 0.560 ;
        RECT 133.130 0.010 133.670 0.560 ;
        RECT 134.510 0.010 135.050 0.560 ;
        RECT 135.890 0.010 136.430 0.560 ;
        RECT 137.270 0.010 137.810 0.560 ;
        RECT 138.650 0.010 139.190 0.560 ;
        RECT 140.030 0.010 140.570 0.560 ;
        RECT 141.410 0.010 141.950 0.560 ;
        RECT 142.790 0.010 143.330 0.560 ;
        RECT 144.170 0.010 144.710 0.560 ;
        RECT 145.550 0.010 146.090 0.560 ;
        RECT 146.930 0.010 147.470 0.560 ;
        RECT 148.310 0.010 148.850 0.560 ;
        RECT 149.690 0.010 150.230 0.560 ;
        RECT 151.070 0.010 151.610 0.560 ;
        RECT 152.450 0.010 152.990 0.560 ;
        RECT 153.830 0.010 154.370 0.560 ;
        RECT 155.210 0.010 155.750 0.560 ;
        RECT 156.590 0.010 157.130 0.560 ;
        RECT 157.970 0.010 158.510 0.560 ;
        RECT 159.350 0.010 159.890 0.560 ;
        RECT 160.730 0.010 161.270 0.560 ;
        RECT 162.110 0.010 162.650 0.560 ;
        RECT 163.490 0.010 164.030 0.560 ;
        RECT 164.870 0.010 165.410 0.560 ;
        RECT 166.250 0.010 166.790 0.560 ;
        RECT 167.630 0.010 168.170 0.560 ;
        RECT 169.010 0.010 169.550 0.560 ;
        RECT 170.390 0.010 170.930 0.560 ;
        RECT 171.770 0.010 172.310 0.560 ;
        RECT 173.150 0.010 173.690 0.560 ;
        RECT 174.530 0.010 175.070 0.560 ;
        RECT 175.910 0.010 176.450 0.560 ;
        RECT 177.290 0.010 177.830 0.560 ;
        RECT 178.670 0.010 179.210 0.560 ;
        RECT 180.050 0.010 180.590 0.560 ;
        RECT 181.430 0.010 181.970 0.560 ;
        RECT 182.810 0.010 183.350 0.560 ;
        RECT 184.190 0.010 184.730 0.560 ;
        RECT 185.570 0.010 199.540 0.560 ;
      LAYER met3 ;
        RECT 0.270 475.680 199.040 511.185 ;
        RECT 1.000 301.560 198.640 475.680 ;
        RECT 0.270 215.920 199.040 301.560 ;
        RECT 1.000 41.800 198.640 215.920 ;
        RECT 0.270 0.175 199.040 41.800 ;
      LAYER met4 ;
        RECT 0.295 0.855 9.320 511.185 ;
        RECT 11.720 0.855 14.620 511.185 ;
        RECT 17.020 0.855 39.320 511.185 ;
        RECT 41.720 0.855 44.620 511.185 ;
        RECT 47.020 0.855 69.320 511.185 ;
        RECT 71.720 0.855 74.620 511.185 ;
        RECT 77.020 0.855 99.320 511.185 ;
        RECT 101.720 0.855 104.620 511.185 ;
        RECT 107.020 0.855 129.320 511.185 ;
        RECT 131.720 0.855 134.620 511.185 ;
        RECT 137.020 0.855 159.320 511.185 ;
        RECT 161.720 0.855 164.620 511.185 ;
        RECT 167.020 0.855 189.320 511.185 ;
        RECT 191.720 0.855 199.330 511.185 ;
  END
END DSP
END LIBRARY

